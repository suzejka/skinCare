���      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.1.3�ub�n_estimators�KȌestimator_params�(�	criterion��	max_depth��min_samples_split��min_samples_leaf��min_weight_fraction_leaf��max_features��max_leaf_nodes��min_impurity_decrease��random_state��	ccp_alpha�t��	bootstrap���	oob_score���n_jobs�NhN�verbose�K �
warm_start��hN�max_samples�Nh�entropy�hKhK	hKhG        h�auto�hNhG        hG        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h6�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C�                                                                	       
                                                                      �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hh.hhhKhK	hKhG        h�sqrt�hNhJY��\hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��h?�f8�����R�(KhCNNNJ����J����K t�b�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGh3�scalar���h?�i8�����R�(KhCNNNJ����J����K t�bC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hK�
node_count�K�nodes�h5h8K ��h:��R�(KK��h?�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hyh\K ��hzh\K��h{h\K��h|h?�f8�����R�(KhCNNNJ����J����K t�bK��h}h�K ��h~h\K(��hh�K0��uK8KKt�b�B�                             �?i����@{	           ��@       	                   �;@�ʹ���@�           �@                            @
��#�d@F           �@                            �?��A�x@�           X�@������������������������       ��nѸ�Q@�           8�@������������������������       ����FO
@;             Y@                           �?��LxO@b           ��@������������������������       ���Ig�N@}            �g@������������������������       �YN�3L@�            �w@
                            @Ѯ����@�            `o@                           �?n�b@c             c@������������������������       ���Mc[)@             E@������������������������       ��ix�@E            �[@                           @^���B�@B            �X@������������������������       �92*%�@-            @P@������������������������       ��c�ۥ�	@             A@                          �3@��S��@�           �@                          �1@�^b��@O           h�@                           @�g�1@$           �~@������������������������       ��Ӝ���
@�            �x@������������������������       �`[)ιb	@<            �X@                            @��2sz�@+            ~@������������������������       �|����
@�            `w@������������������������       ��ӂ�!@B            �Z@                           @r��@A           �@                           @>��,L@Z           ��@������������������������       ��2��@�           P�@������������������������       �(��<$Y@�            �p@                          �:@��D��@�            @x@������������������������       �؁q~�@�             r@������������������������       �����|@-            �X@�t�b�values�h5h8K ��h:��R�(KKKK��h��B`       �s@     �`@     �R@     �w@      D@     �{@      @     �j@      ?@     @|@     �[@     �N@      C@     �Q@      l@     �S@     `v@     �u@     p{@     @W@     �`@     �P@     �G@     �c@      9@     @a@      @     �Y@      7@      a@     �I@     �A@      .@     �E@     �T@      @@     �b@     �c@     �c@      H@     @[@     �D@      B@     �_@      7@     @`@      @      U@      5@      ]@      E@      9@      @      ?@     @R@      8@      a@      a@     �a@     �E@     �O@      9@      6@     �V@      @     �P@              D@      .@      R@      .@      1@      @      3@      F@      2@     @R@      R@      W@      ;@     �J@      6@      6@     �S@      @     �N@              B@      .@     �H@      ,@      0@      @      3@     �C@      2@     �P@      O@     �S@      7@      $@      @              *@              @              @              7@      �?      �?                      @              @      $@      ,@      @      G@      0@      ,@      B@      3@      P@      @      F@      @      F@      ;@       @      @      (@      =@      @      P@      P@     �I@      0@      9@      @      @      &@      @      *@       @      (@      �?      *@      "@      �?              @      @       @      7@      4@      ;@      @      5@      $@       @      9@      (@     �I@      �?      @@      @      ?@      2@      @      @      "@      7@      @     �D@      F@      8@      (@      7@      9@      &@      @@       @       @              3@       @      5@      "@      $@       @      (@      $@       @      (@      5@      *@      @      @      ,@      @      4@              @              ,@      �?      1@      @       @      @      @      @       @      &@      &@      @      @      @      @              @              @               @              @      �?      @      @      �?                      @      @      �?              @      $@      @      0@              �?              (@      �?      &@      @      @      @      @      @       @      @      @       @      @      0@      &@      @      (@       @       @              @      �?      @      @       @      �?      @      @              �?      $@      $@      �?      &@      @      @      $@       @                       @      �?              @       @      �?      @      @              �?      @      @      �?      @      @      �?       @               @              @              @                              �?      �?                      @      @             �f@     @Q@      <@     @k@      .@     Ps@      �?      \@       @     �s@     �M@      :@      7@      ;@     �a@     �G@      j@      h@     �q@     �F@     �H@      8@      @      Y@       @     �c@             �L@              d@      .@      @      @      @     �O@      1@     @U@     �N@     �b@      (@      .@      (@       @      G@       @      W@              ;@             �V@      @      @       @      �?      >@      @     �G@      C@     �O@      (@      "@      @       @      :@       @     @R@              9@             �S@      @      �?       @      �?      4@      @      D@     �@@     �K@      (@      @       @              4@              3@               @              (@               @                      $@              @      @       @              A@      (@      @      K@             �P@              >@             �Q@       @       @      @      @     �@@      *@      C@      7@     �U@              8@      &@      @      D@              L@              1@              O@      @       @      @      @      7@       @      A@      2@     �Q@              $@      �?              ,@              $@              *@               @      @                              $@      &@      @      @      0@             �`@     �F@      7@     �]@      *@     �b@      �?     �K@       @     `c@      F@      5@      2@      6@     �S@      >@      _@     �`@     �`@     �@@     �W@      8@      "@     @U@      (@      ^@             �E@      @     @^@      =@      .@      *@      $@     �K@      8@     �Q@     �X@     �W@      9@     �O@      1@       @     �Q@      @     @X@              @@      @      X@      &@      @      &@      $@     �B@      *@     �H@      Q@     �O@      6@      @@      @      �?      .@      @      7@              &@      @      9@      2@       @       @              2@      &@      6@      ?@      ?@      @     �C@      5@      ,@     �@@      �?      ?@      �?      (@       @      A@      .@      @      @      (@      7@      @     �J@     �@@     �C@       @      8@      3@      @      =@      �?      ;@              $@       @      9@      @      �?       @      @      0@      �?      E@      ?@     �@@       @      .@       @      @      @              @      �?       @              "@      $@      @      @      @      @      @      &@       @      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ!�9<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@�`ߺT�@�	           ��@       	                    �?�B��l@t           �@                           @����@|           p�@                            @��$@           �z@������������������������       �L��a�	@�            �r@������������������������       ���"%+z@R             `@                          �1@���e�
@k            @d@������������������������       �{7׆�
@<            �V@������������������������       ���*�/@/            �Q@
                           @�t5�Р@�           ��@                           �?m��|r)@�             x@������������������������       �?c��4�
@<            @Y@������������������������       ��kĈ�@�            �q@                           @S-(�0@           `{@������������������������       ��u����
@�            �q@������������������������       �O��|��
@c            @c@                           �?�j��'l@0           ��@                           @�k8��z@           (�@                           �?3\����@�           `�@������������������������       ��jq0��@V            `a@������������������������       ��,�]�@P           �@                            �?���Q�{@r             g@������������������������       ���y+T�	@=            @Y@������������������������       �S���
@5             U@                          �7@xm�E�@           ��@                           �?�N]h @           Ȋ@������������������������       �=k�s��@�            Pv@������������������������       ��Y*#F@.           @@                           @U?��@           8�@������������������������       �,�뗲�@�           P�@������������������������       �%�6f��@[            @_@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@     �^@     @X@     �x@     �A@     }@      @     �j@     �A@     �|@     �[@      M@     �@@     �M@     `m@     �Q@     �v@     �q@     �{@      U@     �]@      ?@      8@      d@      @      j@             @S@      �?     @g@      <@      3@      @      @     �R@      0@     @a@     �W@     `i@      .@     �M@      @      @     �I@       @     �X@              D@      �?     @U@      &@      @              @     �B@       @     �G@     �B@     �V@      $@     �F@      @      @      A@      �?     @R@              ,@             @Q@      &@      @              �?      ?@      �?      A@      ;@     �P@      @      2@      @      �?      8@      �?     �K@              "@              M@              @              �?      3@              9@      6@      L@      @      ;@       @      @      $@              2@              @              &@      &@                              (@      �?      "@      @      $@       @      ,@              �?      1@      �?      9@              :@      �?      0@                              @      @      �?      *@      $@      8@      @      @              �?       @      �?      3@              &@               @                              @      @      �?      @      "@      .@      @      &@                      "@              @              .@      �?       @                                      @               @      �?      "@              N@      :@      1@     �[@      @     �[@             �B@             @Y@      1@      .@      @       @     �B@      ,@     �V@      M@     @\@      @      ;@      "@      ,@     �K@      @      G@              5@              7@      ,@      @               @      3@      @      H@      @@     �J@      @       @       @      @      *@              &@               @               @      �?      �?               @      @      �?      @      &@      <@      @      3@      @      &@      E@      @     �A@              3@              5@      *@      @                      *@      @     �D@      5@      9@       @     �@@      1@      @     �K@             @P@              0@             �S@      @      "@      @              2@       @     �E@      :@      N@              6@      @             �D@             �@@              ,@             �M@       @      @      @               @      @      <@      ,@     �C@              &@      $@      @      ,@              @@               @              3@      �?      @                      $@      �?      .@      (@      5@             @l@     �V@     @R@      m@      =@      p@      @     @a@      A@      q@     �T@     �C@      =@     �J@      d@      K@     �l@     @g@     `n@     @Q@     �R@      0@     �@@     �Q@      $@     �W@              O@      @     @Y@     �@@      $@      @      .@     �O@      @     @U@      Q@     �V@      ?@     �J@      *@      8@     �N@      $@     �S@             �M@      @     @R@      6@      "@      @      ,@      G@      @      O@      N@      M@      <@      4@      @      @      $@              1@              *@      �?      (@      @              �?       @      0@              @      $@      .@      @     �@@      $@      4@     �I@      $@     �N@              G@       @     �N@      .@      "@      @      (@      >@      @      M@      I@     �E@      8@      5@      @      "@      "@              0@              @              <@      &@      �?              �?      1@              7@       @      @@      @      .@      @      @      �?              ,@              �?              1@       @      �?                      @              $@      @      3@              @              @       @               @               @              &@      "@                      �?      $@              *@      @      *@      @      c@     �R@      D@     @d@      3@     @d@      @      S@      ?@     �e@     �H@      =@      8@      C@     �X@      H@      b@     �]@      c@      C@      T@      >@      (@      V@      @     @[@             �A@      1@      Y@      8@      1@      0@      "@      I@      ;@     @R@     �P@     �Q@      9@      E@      @       @      A@      @      K@              $@      @     �@@      ,@      @      @      @      8@      @      >@     �E@      @@      @      C@      8@      @      K@      @     �K@              9@      ,@     �P@      $@      ,@      &@      @      :@      5@     �E@      8@     �C@      6@      R@     �F@      <@     �R@      (@     �J@      @     �D@      ,@     @R@      9@      (@       @      =@      H@      5@     �Q@     �I@     �T@      *@     �M@      ?@      <@      Q@      "@      B@      @      ?@      (@     �P@      6@      &@      @      <@      E@      2@      L@      E@     �Q@      *@      *@      ,@              @      @      1@              $@       @      @      @      �?      @      �?      @      @      .@      "@      &@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��)hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@6�5[b@�	           ��@       	                    @/?VT�@S           ��@                            �?|y�̾2@�           0�@                          �1@��^�@�            �s@������������������������       ������@O            �[@������������������������       �,�_�Nb@�             i@                          �2@䌌Ŝ_@�            �r@������������������������       �L���@�            �i@������������������������       � �$�y�	@9            �X@
                           �?:�̟��
@�            �@                           @�M܋(�	@�            �r@������������������������       ��K���X@Y            �b@������������������������       �D�\>۲	@\            �b@                           @^���
@           @}@������������������������       ��+��5m
@�            �t@������������������������       ��	��@P            @a@                           �?8]�eA@G           ƣ@                          �8@i�@�S]@�           �@                           @�[O�u@,           �}@������������������������       �{Oo�O�@�            �p@������������������������       �6#}��@}            `i@                           @y��Ig�@�            �p@������������������������       ��\/��@�             l@������������������������       �z��װ@             D@                           �?V,`qh@p           �@                          �5@t�wdb@�           �@������������������������       ���2��@w             f@������������������������       �2��w�/@(            }@                            �?�)��@�            �@������������������������       �_�Y�"@�            pt@������������������������       ��ш��t@           ȉ@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        t@     �`@     �Y@     �v@     �A@      @      @     �j@      9@     �}@      Y@      N@      ?@     �O@     `l@     �J@     �v@     �r@     @}@      T@     �V@      4@      <@     @a@      @      l@              S@      @     `h@      9@      0@      @      @      S@      &@      a@      W@      k@      1@     �C@       @      7@     �N@      @      T@              8@      @     �P@      5@      @       @      @      F@      @      P@      K@     @W@      &@      ,@      @      (@     �C@      �?     �A@              @      @     �A@      @      @              �?      6@       @      =@      9@     �P@       @      "@      �?      @      ,@      �?      1@               @              &@               @              �?       @      �?      @      (@      6@      �?      @       @      @      9@              2@              @      @      8@      @      @                      ,@      �?      :@      *@     �F@      @      9@      @      &@      6@      @     �F@              2@              @@      0@               @       @      6@      @     �A@      =@      :@      @      ,@      @      @      .@      @      6@              .@              8@       @               @       @      0@      @      4@      9@      3@      @      &@              @      @              7@              @               @       @                              @              .@      @      @             �I@      (@      @     @S@       @      b@              J@              `@      @      &@       @      @      @@      @     @R@      C@     �^@      @      7@              @      9@       @     �M@              5@             �J@      �?                      @      &@       @      =@      .@      H@      @      ,@                      @       @      ?@              �?              ?@      �?                       @       @      �?      5@      @      9@      �?      "@              @      3@              <@              4@              6@                              �?      @      �?       @      "@      7@      @      <@      (@       @      J@             �U@              ?@             �R@      @      &@       @              5@       @      F@      7@     �R@      �?      .@      $@             �C@             �P@              :@             �M@      @      &@       @              .@       @      :@      (@      E@      �?      *@       @       @      *@              3@              @              0@                                      @              2@      &@     �@@             �l@     �\@     �R@     �l@      <@     q@      @      a@      6@     Pq@     �R@      F@      ;@     �L@     �b@      E@      l@     �i@     �o@     �O@     �J@      6@     �@@      P@      @     �T@             �E@              X@      <@      @      @      ,@     �E@       @     @Q@      P@     @R@      =@     �C@      *@      1@     �A@      @      P@             �@@             �K@      *@      �?              $@      7@       @      K@      F@      G@      5@      8@      $@      &@      .@      @      ?@              =@             �B@      @      �?              "@      "@       @      9@      5@      9@      &@      .@      @      @      4@             �@@              @              2@      @                      �?      ,@              =@      7@      5@      $@      ,@      "@      0@      =@              3@              $@             �D@      .@      @      @      @      4@      @      .@      4@      ;@       @      "@      @      *@      =@              2@              $@              @@      ,@      @      @      @      1@      @      (@      3@      .@       @      @       @      @                      �?                              "@      �?                              @              @      �?      (@              f@     @W@      E@     �d@      9@     �g@      @     @W@      6@     �f@     �G@      C@      4@     �E@      [@      A@     `c@     �a@     `f@      A@     @Q@      7@      ,@     �O@      $@     �R@       @      <@      "@     @S@      5@      @       @      @      >@      .@      P@     �E@     �R@      @      &@      @              1@              3@              *@              3@       @      @      @      �?      �?      @      5@      2@      ;@       @      M@      1@      ,@      G@      $@     �K@       @      .@      "@      M@      *@      �?      @       @      =@      &@     �E@      9@      H@      @      [@     �Q@      <@     @Y@      .@      ]@      @     @P@      *@      Z@      :@      ?@      (@      D@     �S@      3@     �V@      Y@      Z@      <@      6@      9@       @      <@      @      @@      @      0@      @      3@      @      (@      @      (@      =@       @      0@      6@      L@       @     �U@     �F@      4@     @R@      (@      U@             �H@      "@     @U@      4@      3@       @      <@     �H@      1@     �R@     �S@      H@      4@�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ _�?hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���{�r@�	           ��@       	                   �:@����@           ��@                           �?�+5 �J@=           `�@                           @�cs�@2           p~@������������������������       ���<͉%@�             p@������������������������       �+����@�            �l@                           @fn�@           ��@������������������������       �e�,���@�           ��@������������������������       ��_�[@�            �k@
                          �;@$��!��@�            �t@                           �?e�7'�@-             P@������������������������       ���x[
@             7@������������������������       �4^�rg
@            �D@                           �?��"�5�@�            �p@������������������������       �Ͱ����@+             N@������������������������       �5�y��@�            �i@                          �6@=j�B@�           ̡@                            �?�,���B@�           �@                           @:pכ�@           @z@������������������������       �?5��7�
@�            �p@������������������������       �H�7�
@Y            �b@                           �?VZ���O@�           |�@������������������������       ��O�c	/
@9           @~@������������������������       �����@�           ؅@                           �?EH=:�b@�           �@                            �?���w3@�             t@������������������������       �[����P@w            �e@������������������������       ��|iN�@W            @b@                           @�U��@�            0v@������������������������       �
��G@�             l@������������������������       �&!�v��@U            @`@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        s@     �b@     �U@     �s@      A@     0~@      *@     �m@      7@     �~@     �W@      M@      A@      P@     �l@      L@     �v@      t@     p}@     @S@     �a@     �Q@      L@     �`@      :@     �b@      "@     @[@      1@      d@     �H@     �A@      4@     �E@     �X@      4@     �b@     �`@     �d@      F@     �_@      E@     �C@     @Y@      6@     @a@      @     @S@      1@     �a@     �@@      6@      &@      @@     �T@      *@     ``@      X@      a@      C@     �J@       @      (@     �B@      @     �P@      @      7@      @     �O@      $@      @       @       @      ;@      @      I@     �A@      O@      ,@      1@      @      @      4@      �?      E@      @      .@             �D@      @      @       @       @       @      @      8@      5@      @@       @      B@      @      @      1@      @      8@               @      @      6@      @       @                      3@              :@      ,@      >@      @     @R@      A@      ;@      P@      .@      R@       @      K@      ,@     @S@      7@      0@      "@      >@      L@      $@     @T@     �N@     �R@      8@      K@      5@      7@      K@      @     �F@       @     �C@      $@     �I@      6@      *@      @      2@     �E@      @     �H@      J@     �L@      8@      3@      *@      @      $@      "@      ;@              .@      @      :@      �?      @      @      (@      *@      @      @@      "@      2@              .@      =@      1@      A@      @      (@      @      @@              5@      0@      *@      "@      &@      0@      @      3@      C@      =@      @      @              @      @      �?       @       @      $@              �?               @              �?      @      �?      @      *@      @      @      �?              @      @                       @       @                              �?                       @              �?      @      �?      @      @              �?      @      �?       @               @              �?              �?              �?       @      �?       @      $@      @              &@      =@      (@      <@      @      $@      �?      6@              4@      0@      &@      "@      $@      (@      @      0@      9@      7@      @      @      @      �?      @              @              @              @       @      @      @              �?      �?      @      �?      &@              @      7@      &@      8@      @      @      �?      2@              *@      ,@       @      @      $@      &@      @      (@      8@      (@      @     �d@     �S@      >@      g@       @     �t@      @     �_@      @     �t@     �F@      7@      ,@      5@     �`@      B@     �j@     @g@     s@     �@@      X@      G@      6@      a@      @     Pp@             �W@      @     �n@      7@      2@       @       @     @T@      0@     �d@     �_@      l@      4@      3@      .@      &@     �F@             �P@              ,@      �?     @S@      @      @      @      �?      (@      �?      E@     �A@     �M@      @      3@      @      @      <@              E@              $@      �?      P@      @      @      @              @      �?      9@      0@     �@@      @              (@      @      1@              9@              @              *@               @      �?      �?      @              1@      3@      :@             @S@      ?@      &@      W@      @     @h@              T@      @     @e@      0@      (@      @      @     @Q@      .@     �^@      W@     �d@      1@      >@       @              E@      �?     �Y@              :@              H@       @       @              @      >@              G@      A@      X@      @     �G@      7@      &@      I@       @     �V@              K@      @     �^@       @      $@      @      @     �C@      .@     @S@      M@     �Q@      &@     @Q@     �@@       @     �G@      @      R@      @     �@@             @U@      6@      @      @      *@     �I@      4@      I@     �M@      T@      *@      =@      @      @      ;@      @      A@      @      4@             �E@      *@      �?      @       @      :@      (@      1@      @@      A@      &@      0@      @      �?      *@      @      7@              *@              :@      "@                       @      *@      @      $@      *@      2@      @      *@               @      ,@      �?      &@      @      @              1@      @      �?      @              *@       @      @      3@      0@      @      D@      <@      @      4@      �?      C@              *@              E@      "@      @      @      &@      9@       @     �@@      ;@      G@       @      5@      3@       @      &@      �?      @@              @             �@@      @      @      @      @      .@       @      7@      1@      9@       @      3@      "@      @      "@              @              $@              "@      @                      @      $@      @      $@      $@      5@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ&h>hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �3@yxV��@�	           ��@       	                    @�{�oN�@~           ��@                           @;�A�@�           t�@                          �1@ �Z�2@�           h�@������������������������       ����6�@�            �q@������������������������       ������@�            0u@                            @�$�x1%@=            @������������������������       ��u�o�n
@	           �y@������������������������       �J�+#�7	@4             V@
                           @\��s��@�             r@������������������������       ��nv��@             7@                           @n�$M5�@�            �p@������������������������       ���f@j             e@������������������������       �����3@@            �X@                          �;@�q�I9@<           ��@                          �:@��J���@,           B�@                           �?~Ը@�           \�@������������������������       �`T�:�@           ��@������������������������       ��%��op@�           �@                           @���c�@]            @a@������������������������       ���#+�
@)            �P@������������������������       �2�p��B@4            �Q@                           @!�}FL�@           �z@                           �?�ۘ��@�            �r@������������������������       ���G�^�@�            �n@������������������������       ���g�
@"            �I@                           �?��e��@L             `@������������������������       ����&��@             I@������������������������       �O%'�@.            �S@�t�bh�h5h8K ��h:��R�(KKKK��h��B        �t@     �a@     @V@     pv@     �A@      ~@       @     @h@      <@     |@     @^@      J@      C@      S@     �i@     �K@     @w@     pu@     `|@     @S@      [@     �E@      <@     �`@      @     �i@              T@      @     �f@      ?@      *@      @      (@     �R@      2@      \@     @[@     @l@      0@     �S@      :@      4@     @Y@      @      d@             �Q@      @     �c@      6@      $@      @      (@     �M@      0@     �W@     @Q@     �g@      ,@     �@@      .@      ,@     �P@      @     �R@              9@      �?     @T@      4@      @              @      D@      *@     @P@      F@     �X@      (@      2@       @      $@      4@      @      H@              (@             �E@      "@       @               @      5@      @      9@      5@     �A@      @      .@      *@      @      G@       @      ;@              *@      �?      C@      &@      @              @      3@      @      D@      7@     �O@       @      G@      &@      @     �A@      �?     �U@              G@      @     �S@       @      @      @      @      3@      @      >@      9@     �V@       @      :@      $@      @      A@             �Q@              >@      @      Q@      �?      @      @              3@       @      <@      3@      U@      �?      4@      �?      �?      �?      �?      .@              0@              $@      �?                      @              �?       @      @      @      �?      =@      1@       @      A@             �F@              "@              6@      "@      @                      0@       @      1@      D@     �B@       @              @              �?                                              @       @      �?                      @              �?      "@                      =@      ,@       @     �@@             �F@              "@              3@      @       @                      *@       @      0@      ?@     �B@       @      3@       @      @      8@              @@              @              *@      @       @                      "@              @      1@      5@       @      $@      @      �?      "@              *@              @              @       @                              @       @      $@      ,@      0@              l@      Y@     �N@      l@      =@     @q@       @     �\@      8@     �p@     �V@     �C@      A@      P@     @`@     �B@     @p@     @m@     �l@     �N@      h@     �Q@     �G@      i@      4@     �o@       @     �U@      4@     �k@     �O@      A@      1@      I@     �[@      @@     @l@     �h@     `f@      K@     �f@     �Q@     �E@     �f@      4@     �n@      @     �S@      2@     �j@      M@      ;@      0@     �G@     @W@      ;@     �k@     �e@      e@     �J@      T@     �A@      4@      N@      .@     @U@      @      H@      .@      W@      :@      1@      @      ?@     �B@      2@     @Z@     �P@      P@      ;@     @Y@     �A@      7@     �^@      @      d@              >@      @     �^@      @@      $@      $@      0@      L@      "@     �\@      [@     @Z@      :@      (@              @      1@              @       @      "@       @      @      @      @      �?      @      2@      @      @      7@      $@      �?      @                      "@              �?              @       @       @      @       @               @      "@      �?      �?      4@      @      �?      @              @       @              @       @      @              @       @      @      �?      �?      "@      @      @      @      @              @@      >@      ,@      8@      "@      8@              ;@      @     �G@      ;@      @      1@      ,@      3@      @      A@     �B@     �H@      @      7@      9@      (@      0@      "@       @              2@      �?      A@      0@      @      0@      "@      *@      @      7@      <@      >@      @      *@      7@      (@      .@      @      @              2@      �?      5@      .@      @      ,@      "@      &@      @      6@      7@      8@      @      $@       @              �?       @       @                              *@      �?               @               @      �?      �?      @      @      @      "@      @       @       @              0@              "@      @      *@      &@      �?      �?      @      @      �?      &@      "@      3@              �?      @                              (@                      @      @      @                      �?      �?      �?      �?      @      @               @       @       @       @              @              "@              @      @      �?      �?      @      @              $@       @      *@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJDr�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@�{����@�	           ��@       	                     @�ri��@e           ��@                           @��$
�@|           0�@                            �?�ϹQ��@�           Є@������������������������       ��S��@K           H�@������������������������       ��.8)��@a             b@                          �2@~Z���@�            �t@������������������������       ��X�嗀@�            �n@������������������������       �y;�c��	@4            @U@
                           @����g@�            �u@                          �2@0���i@�            �q@������������������������       ���Q��Z@�             i@������������������������       �J`�y�
@=            �U@                           �?���N��@(             M@������������������������       ���gi�@             B@������������������������       �S:uc@             6@                           �?��ҙ�v@(           �@                            @<=T�ɽ@�           �@                           �?ά��B@�           `�@������������������������       �+�����@�            `p@������������������������       �����M@E           0�@                           @�f��&�@�            �p@������������������������       �뇶a�@o            �f@������������������������       ��5��K
@7            @V@                           @�U�=�@�           D�@                           �?�*��F�@:           ��@������������������������       ��%�2@           ��@������������������������       ���&���@5           P}@                            �?D��Yw�@f             e@������������������������       ��;���k@D            �[@������������������������       ��Sm0��	@"            �M@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �^@     @V@     Px@     �E@     �}@      &@     �o@      >@     0{@     �Z@     �I@      @@      M@      q@      O@     �v@     0s@     �y@     �W@     �R@      A@      5@      c@       @     �h@             �V@      �?      f@      >@      (@      @      @      U@      2@      a@     �W@     @g@      8@     �F@      :@      (@     �\@      �?     @b@              M@      �?     @a@      ,@      @      @       @     �P@      &@     �Z@      R@     `c@      2@      >@      ,@      @     �Q@      �?      Y@             �D@      �?     @\@      @      @      @      �?     �J@      @     �Q@     �C@      W@      *@      ;@      ,@      @     �L@             �Q@             �B@      �?      V@      @      @      @              F@      @      I@      @@     �P@      (@      @               @      *@      �?      >@              @              9@               @              �?      "@              5@      @      :@      �?      .@      (@      @     �F@              G@              1@              9@      $@      �?              �?      *@      @     �A@     �@@     �O@      @      *@      @      @      D@              >@              *@              9@      @      �?              �?      &@      @      3@      6@      H@       @       @      @      �?      @              0@              @                      @                               @      �?      0@      &@      .@      @      =@       @      "@     �B@      �?     �I@             �@@              C@      0@      @               @      2@      @      ?@      7@      ?@      @      :@      @      @      :@      �?     �D@              8@              ;@      0@      @                      1@      @      ?@      5@      ;@      @      0@      @       @      6@      �?      ;@              *@              4@      @      @                      *@      @      9@      .@      2@      @      $@              @      @              ,@              &@              @      &@                              @              @      @      "@              @       @       @      &@              $@              "@              &@                               @      �?                       @      @      �?       @       @      �?      &@              @              @               @                                      �?                              @      �?      �?              �?                      @              @              "@                               @                               @      �?              n@      V@      Q@     �m@     �D@     @q@      &@     �d@      =@     0p@     @S@     �C@      ;@      K@     �g@      F@     �k@     �j@     �k@     �Q@     @_@      8@      A@      V@      .@     �`@      "@     �Q@      $@     �_@      ?@      "@      $@      *@     @R@      $@     �Q@     �Y@     @W@      B@      X@      0@      *@      Q@      (@     @\@      @     �F@      @     �W@      ;@      @      "@      @      N@       @     �M@     �S@      O@      =@      >@      @      @      7@      @      0@      @      :@      �?      <@      @      @      �?      @      ;@      @      8@      6@      0@      @     �P@      (@      @     �F@      @     @X@      @      3@      @     �P@      4@      �?       @      @     �@@      @     �A@      L@      G@      6@      =@       @      5@      4@      @      3@       @      9@      @      @@      @      @      �?      @      *@       @      (@      8@      ?@      @      4@      @      5@      .@      @      (@       @      3@      @      &@       @      @      �?      @      @       @      "@      1@      3@       @      "@       @              @              @              @              5@       @                              $@              @      @      (@      @      ]@      P@      A@     �b@      :@      b@       @     �W@      3@     �`@      G@      >@      1@     �D@     �\@      A@      c@     �[@      `@      A@      Z@     �M@      8@     �`@      :@     �^@       @      W@      3@      _@      E@      >@      0@      @@     �V@      A@     �`@     @Y@     �Z@      >@      J@     �E@      3@      W@      6@      P@       @      N@      1@     �P@      =@      5@      *@      >@     �N@      8@     �U@     @P@     �N@      6@      J@      0@      @     �D@      @     �M@              @@       @     �L@      *@      "@      @       @      =@      $@     �F@      B@      G@       @      (@      @      $@      0@              5@               @              "@      @              �?      "@      9@              4@      "@      6@      @      (@       @      @      "@              1@               @              @      @                      @      ,@              $@      @      5@      @              @      @      @              @                              @                      �?      @      &@              $@      @      �?        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��d$hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�_~x�@�	           ��@       	                    �?,0�@�           F�@                          �3@�SQ� �@c           ��@                          �2@P�|�H
@            �y@������������������������       ��J�ٵ�	@�            @s@������������������������       ��N�{l	@@             Y@                          �;@c>�d�@c            �@������������������������       �Ξ��q�@.           `~@������������������������       �F}�n�@5            �V@
                           @�o��@�           ,�@                            �?_f�=�C@<           ȍ@������������������������       �v�m�%�@!            ~@������������������������       ����@           �}@                          �6@q�2V�)@D           ��@������������������������       �`3�6�@�           P�@������������������������       �3g�X�@�            �r@                           @p����@�           ��@                           �?��"�VZ@?           �@                          �4@/��{��@�            �r@������������������������       �A��B�@I            �[@������������������������       ��eC0O@y            �g@                           �?�o�5�@}            @j@������������������������       �XһA��@=            @X@������������������������       �X�`>W�
@@            @\@                           @%��DV@k           H�@                           @���1�@           �y@������������������������       ��<3 8I@V            �`@������������������������       �����@�            �q@                          �3@3�0�@X            @a@������������������������       �h�7�@             D@������������������������       �L�YI�	@=            �X@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �`@     @S@     0v@     �G@     @      $@     �k@      6@     �|@      W@     �S@     �@@     �P@     �o@      J@     �w@     �r@     z@     @V@     �l@     �W@      F@     0p@      6@     �x@      @     `b@      1@     �v@     �N@     �J@      :@      A@     �g@     �B@     �p@     �i@     �u@      M@     �S@      2@      .@      V@      @      c@             �O@       @     �a@      9@      ,@      @      @      N@      @     �R@     @Q@     `a@      7@      1@      @      @     �F@      �?     �T@              8@       @     @P@       @      "@               @      <@       @      :@      4@     �R@       @      (@      �?      @      ?@      �?     �O@              4@      �?      I@      �?      �?               @      5@       @      6@      3@      L@       @      @       @              ,@              3@              @      �?      .@      �?       @                      @              @      �?      3@              O@      .@      (@     �E@      @     �Q@             �C@              S@      7@      @      @      @      @@       @      H@     �H@      P@      5@      N@      $@       @      D@       @     @P@             �B@             �M@      *@       @      �?      @      =@       @      D@      D@     �J@      5@       @      @      @      @       @      @               @              1@      $@      @      @              @               @      "@      &@             �b@      S@      =@     `e@      1@     @n@      @      U@      .@     `k@      B@     �C@      4@      <@     @`@     �@@     �h@     �`@     �i@     �A@     �S@      D@      ;@      X@      ,@     �W@      @     �J@       @      V@      2@      1@      @      1@     �T@      4@     @Y@      Q@      W@      :@      <@      >@      (@     �E@      "@      F@      @     �@@      @      =@      @      $@      @      &@     �D@      @     �G@      D@     �M@      ,@      I@      $@      .@     �J@      @     �I@              4@      @     �M@      &@      @              @      E@      ,@      K@      <@     �@@      (@     �Q@      B@       @     �R@      @     `b@       @      ?@      @     ``@      2@      6@      *@      &@     �G@      *@     �W@     �P@     �\@      "@      =@      8@      �?     �K@             �\@              6@      @     �X@      &@      3@      "@              >@      @      P@      F@     @V@      @      E@      (@      �?      4@      @     �@@       @      "@      @     �@@      @      @      @      &@      1@      $@      ?@      7@      9@      @     @Z@      D@     �@@      X@      9@     �Y@      @      S@      @     @X@      ?@      9@      @      @@      P@      .@     @[@     �W@      R@      ?@      H@      2@      *@      D@      &@      J@       @     �D@       @     �C@      0@      .@              8@     �D@      @     �H@      F@      B@      *@      6@      (@      (@      8@      @      9@       @      ;@       @      ,@      $@      *@              6@      6@      @      =@      >@      .@      @      ,@      �?      @      �?      @      ,@              "@      �?      @      @      @              @       @       @      *@      @      $@               @      &@      @      7@      @      &@       @      2@      �?      &@      @      @              1@      ,@      @      0@      7@      @      @      :@      @      �?      0@      @      ;@              ,@              9@      @       @               @      3@              4@      ,@      5@      @      @      �?      �?      &@      @      0@              @              @      @       @                       @              @      @      0@      @      6@      @              @      �?      &@               @              2@      �?                       @      &@              ,@      "@      @      �?     �L@      6@      4@      L@      ,@      I@      �?     �A@      @      M@      .@      $@      @       @      7@      $@      N@      I@      B@      2@      B@      5@      2@     �C@      ,@     �D@      �?      <@      @      >@      .@       @      @      @      0@      @      E@      C@      ?@      .@      (@       @      @      "@       @      *@      �?      @       @      $@       @      @      @      @       @      �?      "@      "@      (@      @      8@      *@      &@      >@      @      <@              8@      �?      4@      @       @      @      @      ,@      @     �@@      =@      3@       @      5@      �?       @      1@              "@              @              <@               @              �?      @      @      2@      (@      @      @      @      �?      �?      $@              @              @              @              �?                      �?      @      �?      �?                      ,@              �?      @              @              @              6@              �?              �?      @              1@      &@      @      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ� LhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@W�؜�@�	           ��@       	                   �3@�*3��@a           ��@                            �?�]s��@l           ��@                           �?續@            ��@������������������������       �rB%F�
@�            `y@������������������������       �����@
           �y@                            @
l��@l           ��@������������������������       ���8xJ�
@�            �k@������������������������       �A�?�&}@�            v@
                           @�H'�@�             x@                           �?��丕@�            @r@������������������������       �����
@H            @]@������������������������       �8a4@n            �e@                            �?Y��d�@?             W@������������������������       �$�}���@             8@������������������������       ��� ��@-             Q@                          �:@��p@P           ��@                          �5@ +0e��@�           4�@                           �?5�p%�@�            �w@������������������������       ��sß@Y            @c@������������������������       ���{a�@�             l@                          �6@�ߺ�@           H�@������������������������       ��?V��@�            �q@������������������������       �3�HU
�@J           ��@                          �;@xOb���@j           `�@                           @���/@[            �a@������������������������       ��&F�9@E            �[@������������������������       ��bf]O?	@             >@                           �?ײ�Au�@           �{@������������������������       ��=�1�@<            @Y@������������������������       �W"d��s@�            �u@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     `c@     �X@     �u@     �B@     0}@      @     �j@      9@     @}@      X@     @P@      ?@     �R@      p@     �P@      v@     �s@     0|@      N@     �`@      E@      B@     �c@      ,@     �o@              U@      @     `m@      7@      7@      $@      2@      ^@      7@     �c@     �c@     �o@      :@     �Y@      =@      ;@      a@      @     �i@             �P@      @     �g@      7@      3@      @      .@     �U@      2@     �_@     �\@      j@      $@      J@      3@      (@     �W@      �?     @Y@              @@      @     @_@      (@      *@       @      @      H@      $@     �S@     �N@     �a@      @      =@      "@      @     �D@             �G@              2@              T@      @      @       @              4@      �?      D@      <@     �R@      @      7@      $@      @      K@      �?      K@              ,@      @     �F@      "@      "@              @      <@      "@      C@     �@@     �P@       @      I@      $@      .@     �D@      @     �Z@             �A@             �P@      &@      @       @      "@      C@       @      H@     �J@     �P@      @      .@      @      �?      0@       @     �K@              1@              :@              @      �?      @      0@              5@      0@      7@      �?     �A@      @      ,@      9@      @     �I@              2@              D@      &@       @      �?      @      6@       @      ;@     �B@     �E@      @      @@      *@      "@      5@      @      G@              1@      @      F@              @      @      @      A@      @     �@@      F@     �G@      0@      =@      @       @      4@      @      C@              .@       @      @@              @      @      �?      9@      @      7@     �A@      ?@      (@      (@      �?      @      @              4@              "@              1@                       @               @              @      *@      1@      @      1@      @      @      *@      @      2@              @       @      .@              @      @      �?      1@      @      4@      6@      ,@      "@      @      "@      �?      �?       @       @               @      �?      (@              �?      �?       @      "@      �?      $@      "@      0@      @      �?              �?                       @              �?              @              �?                      @              �?      �?      @       @       @      "@              �?       @      @              �?      �?      @                      �?       @      @      �?      "@       @      *@       @     @h@     @\@     �O@     �g@      7@     �j@      @      `@      3@      m@     @R@      E@      5@     �L@      a@     �E@     `h@     `c@     �h@      A@     �`@     @V@      D@     �b@      *@      g@      �?     �U@      ,@      g@      H@      8@      "@      D@     �V@      9@     �b@     �Z@     �_@      @@      >@      ?@      @     �G@             �K@              2@      @      F@      @      0@      @      @      1@      @     �C@      ;@      4@      @      0@      .@      @      4@              5@              &@      @      4@      �?      @              @       @      �?      8@       @              �?      ,@      0@              ;@              A@              @              8@      @      *@      @      @      .@      @      .@      3@      4@      @     @Z@      M@      B@     �Y@      *@      `@      �?      Q@      $@     �a@     �D@       @      @      A@     @R@      4@      \@      T@     �Z@      ;@      0@      "@      &@      1@      @     �J@              5@      @      E@      *@       @              @      6@      @      8@      "@      4@      @     @V@     �H@      9@     �U@       @      S@      �?     �G@      @     �X@      <@      @      @      ;@     �I@      1@      V@     �Q@     �U@      5@     �M@      8@      7@     �D@      $@      >@      @     �E@      @      H@      9@      2@      (@      1@      G@      2@      F@      H@     �Q@       @      *@              @      3@              (@      @      (@      �?       @       @      "@      �?       @      .@      @      &@      $@      5@              @              @      *@              $@      @      (@      �?      �?      �?      @                      (@      @      @      $@      4@              @                      @               @                              �?      �?      @      �?       @      @              @              �?              G@      8@      3@      6@      $@      2@       @      ?@      @      G@      7@      "@      &@      .@      ?@      ,@     �@@      C@     �H@       @      @      �?      @      @       @      $@               @              1@      �?      @      @      @      @      @      @      @      &@       @     �D@      7@      (@      0@       @       @       @      7@      @      =@      6@      @      @      (@      ;@      $@      :@      A@      C@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJyt hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@f�+��Z@�	           ��@       	                     @�h�4/q@           ��@                           �?z��O��@r           D�@                           @&��B�C@�           ��@������������������������       ��t�=�
@_           ��@������������������������       ���4&�
@H            �[@                          �1@=4���@�           Ȑ@������������������������       �:u��Y�@�            �r@������������������������       �$&,P�@           (�@
                          �3@�4��~@�           0�@                           @�Ƨ} ~@�            �y@������������������������       �J6�N�@@�            �v@������������������������       ���"o\�
@             H@                           �?:%Q�=@�            @m@������������������������       ��eh�d@Y            @`@������������������������       ��Oy�B@G             Z@                          �<@�W=^G@�           ȗ@                          �:@�c���@�           ��@                            @BR� �@S           ��@������������������������       �NO֖�@�           Ѓ@������������������������       ������D@�            �s@                           �?�-�^�@�            �m@������������������������       ��:����@2             T@������������������������       ��["U�@d            �c@                          �>@�l��.�@�            �t@                          �=@�����@_            �c@������������������������       ��t��.
@:            �V@������������������������       ��uRg&
@%             Q@                           �?΍��w@y             f@������������������������       ���L�F@W            �`@������������������������       ���B�z�	@"            �F@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �a@      W@     pw@      1@     p}@      @     �m@      ?@     p|@      ^@      L@     �@@     �I@     `n@     �J@     �t@     �s@     `}@     �T@     `g@      Q@     �J@      n@      @     `v@      �?     �a@      2@     �q@      N@     �C@      &@      0@     @^@      ;@     �i@     �f@     0t@      F@     �^@      H@      @@     �f@      @     �q@             �V@      1@     �k@      C@      >@      $@       @     �U@      0@     @b@     �^@     @p@     �@@      E@      0@      @     �P@       @     �`@             �B@       @     @V@      "@      @              @      B@             �M@     �F@     @Z@      *@      ?@      &@      @      O@       @     @^@             �@@      �?     �S@      @      @              @      :@              H@      @@     �T@      *@      &@      @              @              *@              @      �?      $@      @                      �?      $@              &@      *@      7@              T@      @@      :@     �\@       @     `b@             �J@      .@     ``@      =@      :@      $@      @     �I@      0@     �U@     @S@     `c@      4@      7@      @      @      9@      �?      D@              ;@             �D@      @      �?               @      &@      @      ;@      ;@      J@      @     �L@      ;@      5@     @V@      �?     �Z@              :@      .@     �V@      8@      9@      $@      �?      D@      (@      N@      I@     �Y@      .@     @P@      4@      5@     �M@      @     @S@      �?     �J@      �?     �P@      6@      "@      �?       @      A@      &@     �N@      N@     �O@      &@     �G@      "@      *@     �C@       @     �N@      �?     �C@             �B@      ,@       @      �?      @      8@      "@      @@     �@@      D@      @     �E@      @      *@      ?@       @      L@      �?     �@@             �@@      ,@      �?      �?       @      5@      "@      @@      :@     �B@      @      @      @               @              @              @              @              �?              �?      @                      @      @       @      2@      &@       @      4@      �?      0@              ,@      �?      =@       @      @              @      $@       @      =@      ;@      7@      @      ,@      @       @      "@      �?      @              @      �?      ,@      @      @              @      @       @      0@      3@      @      �?      @      @              &@              &@              "@              .@      �?      �?                      @              *@       @      0@      @     `b@     @R@     �C@     �`@      $@     @\@      @     �W@      *@      e@      N@      1@      6@     �A@     �^@      :@     �_@     �`@     `b@      C@      ]@      F@      6@     �Z@      "@      V@      @     �S@      *@     �a@     �C@      0@      "@      <@     @V@      8@     �\@      Z@      \@     �@@     �Y@      B@      3@      R@       @     �T@       @     �N@      "@     �^@      A@      @       @      7@      S@      0@     �T@     �S@     �U@      8@     �S@      ;@      (@      I@      @     �I@       @      B@      �?     �V@      3@      @       @      &@      I@      ,@      I@      F@      R@      .@      7@      "@      @      6@       @      @@              9@       @      @@      .@      @      @      (@      :@       @     �@@      A@      ,@      "@      ,@       @      @      A@      �?      @      �?      1@      @      2@      @      "@      �?      @      *@       @      ?@      :@      :@      "@      @              @      1@      �?              �?      @      @       @      �?      �?      �?       @      @       @      ,@       @      @       @      &@       @              1@              @              ,@              $@      @       @              @      $@      @      1@      2@      4@      @      ?@      =@      1@      =@      �?      9@              1@              =@      5@      �?      *@      @     �@@       @      (@      <@     �A@      @      4@      @      @      &@              @              @              .@      .@              @       @      :@      �?      @      .@      1@       @      "@      @      @      @              @              @              @      $@              @      �?      1@      �?       @      @      0@              &@       @              @                               @              &@      @               @      �?      "@              @      (@      �?       @      &@      6@      (@      2@      �?      5@              &@              ,@      @      �?      @      @      @      �?      @      *@      2@      @      @      4@      "@      0@      �?      *@              &@              "@      @      �?      @      @      @      �?      @      (@      "@       @      @       @      @       @               @                              @      �?                              @              @      �?      "@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�b��      hGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@8�c�[�@�	           ��@       	                    �?�"2!�4@`           ��@                            �?}d^�� @           ��@                           @'W�_�@�            `m@������������������������       ���H�ɿ
@u            �g@������������������������       �Z.t:@!            �F@                           @P�I�.�@�           H�@������������������������       ��(�Ae0@�            �j@������������������������       ���3�
@�            0y@
                           @-#���@G           Ȍ@                            �?0�L/��@�           ��@������������������������       �%� O�l@�            �w@������������������������       �֟s��6@�            �q@                            �?]��y�@�            0p@������������������������       �ݠ�  <@\            �b@������������������������       �?��^xH	@F             [@                           �?�ROq|@X           ��@                           @��f�	@�           P�@                           �?��{Y�#@�           x�@������������������������       ���1��/@�             l@������������������������       �#���#-@S           p�@                            �?uC�19�@�            Pr@������������������������       �.����@?             V@������������������������       ���b��@�            �i@                           @�UDhj|@�            �@                          �5@�t^5�@�           Ѓ@������������������������       �y��R8@A            @X@������������������������       �}��,@K           Ȁ@                          �9@�)��ղ@!           �|@������������������������       ��<�p�@�            �t@������������������������       ��P��|!@X            �`@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       0u@      a@     �S@      w@     �A@     �@      (@     �j@      9@     �{@      ]@      N@      F@      Q@     `m@     �P@     �t@     ps@     �z@     �U@     �]@      E@      8@     �f@      .@     Pq@      @     @U@      &@     `m@      B@      @@       @       @     �Y@      6@     �b@     �a@     �n@      A@     �M@      3@      @     �T@       @     �a@              H@             �Z@      ,@      &@       @       @     �F@      @      P@      V@     �`@      3@      1@      @      @      9@              <@              0@             �G@       @       @       @              (@              7@      3@      9@      $@      ,@      @              2@              5@              ,@             �F@       @       @      �?              $@              5@      (@      3@       @      @      �?      @      @              @               @               @                      �?               @               @      @      @       @      E@      .@      @      M@       @     �\@              @@             �M@      (@      "@               @     �@@      @     �D@     @Q@      [@      "@      5@      @      �?      .@      @     �@@               @              3@      "@                              *@      @      8@      ;@      ;@      @      5@       @       @     �E@      @     @T@              8@              D@      @      "@               @      4@              1@      E@     @T@      @     �M@      7@      2@     �X@      @     �`@      @     �B@      &@      `@      6@      5@      @      @     �L@      3@     �U@     �K@      \@      .@     �E@      .@      $@     �U@      @      X@      @      2@       @     @T@      0@      1@      �?      @     �F@      1@      Q@     �E@     @R@      $@      .@      @      @     �L@              O@              @      @      J@       @      *@              @      3@      ,@      C@      6@      H@      @      <@      $@      @      =@      @      A@      @      *@      @      =@       @      @      �?              :@      @      >@      5@      9@      @      0@       @       @      (@             �C@              3@      @      H@      @      @      @       @      (@       @      3@      (@     �C@      @      *@       @      �?      &@              .@              ,@      @      5@      @       @      @              @       @      @       @      <@      @      @              @      �?              8@              @              ;@       @       @               @      @              *@      @      &@       @     �k@     �W@      K@     `g@      4@      m@       @      `@      ,@     �j@      T@      <@      B@      N@     �`@      F@     �f@      e@      g@     �J@     �V@     �K@     �@@     �W@      ,@     �Q@      @     �U@      $@     @Z@      A@      .@      6@      B@     �N@      ;@     @U@     �U@     �V@      8@     �O@      A@      9@     @R@      $@      J@      @      R@      @      P@      @@      (@      2@      :@     �F@      3@     �N@      L@     �M@      2@      9@      $@      "@      6@              8@      @      5@       @      ,@      @      @      @      @      (@      @      0@      ,@      :@      @      C@      8@      0@     �I@      $@      <@       @     �I@      @      I@      :@       @      .@      7@     �@@      *@     �F@      E@     �@@      *@      ;@      5@       @      5@      @      2@              .@      @     �D@       @      @      @      $@      0@       @      8@      >@      @@      @      @       @              @       @      @              @       @      &@              �?       @      @      @      @      @      @      &@      @      8@      *@       @      0@       @      &@              &@      �?      >@       @       @       @      @      &@      @      4@      7@      5@      �?     ``@     �C@      5@     @W@      @     @d@      @      E@      @     �Z@      G@      *@      ,@      8@      R@      1@     �X@     �T@     @W@      =@     @Q@      9@      .@      J@      @     �Y@              A@       @     �P@      4@      @      $@      *@     �F@      .@     �G@     �D@      F@      8@      @      @      �?      @              7@              @              @      @      @      @      @      @      @       @      @      @      @     @P@      2@      ,@     �G@      @     �S@              >@       @     �O@      1@      @      @      "@     �D@      &@     �C@     �B@      C@      2@      O@      ,@      @     �D@      @      N@      @       @       @      D@      :@      @      @      &@      ;@       @     �I@     �D@     �H@      @     �B@      "@      @      B@       @      H@              @       @     �@@      0@      @              @      .@       @      D@     �@@     �A@      @      9@      @      @      @      �?      (@      @       @              @      $@      @      @      @      (@              &@       @      ,@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�o:}hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�H�"�@�	           ��@       	                   �5@�M�Zn�@           ԙ@                           �?�!��+�@�           ��@                            @�����@�             s@������������������������       ��U�(7 @f            �d@������������������������       ��5o/8@S            @a@                            @�4�`@           �|@������������������������       �-�b"L@�            0r@������������������������       �����=@c            �d@
                           @����)@M           �@                            @��:� C@�           h�@������������������������       ��6���@�            �u@������������������������       ��Ӯ]$@�             s@                          �;@Xu�Y��@�             n@������������������������       �� U�Ȋ@o            `c@������������������������       ����@>            @U@                            @�z�!��@�           ��@                          �4@���!Ӑ@~           ��@                           @JW��H�
@W           �@������������������������       ���qj� 
@�           ��@������������������������       �JD�׏�
@�            �s@                          �;@��f��@'           ��@������������������������       ��BD?O@�            �@������������������������       �c�B�@W            �a@                           �?~�v�L@           @z@                          �9@( B��@o            �f@������������������������       ��a���	@_            @c@������������������������       �<��]b@             <@                           @515�.@�            �m@������������������������       �LG*�@0            �S@������������������������       ��}0bK@d            �c@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       @s@     �_@     @Y@     pt@     �A@     p�@       @     �k@     �@@     �}@     �Y@     �P@      =@     �O@     �i@     �K@      v@     pt@     P|@     �W@     @]@     �Q@     @P@     �b@      9@     `d@      @     �[@      ;@     �c@     �H@      G@      .@      D@     @U@      B@      a@     `c@     �c@     �F@     @Q@      .@      5@     @U@      ,@     @U@             �C@      &@     @T@      3@      ;@      @      @      C@      &@      N@     @Q@     @S@      =@      ?@      @      @      :@      @      G@              (@             �@@      $@      @       @      �?      4@      �?     �@@      ;@     �B@      @      &@      @      �?      1@      �?      9@              @              7@       @      @              �?      &@      �?      1@      &@      ;@      @      4@              @      "@       @      5@              @              $@       @               @              "@              0@      0@      $@      @      C@      $@      .@     �M@      &@     �C@              ;@      &@      H@      "@      6@      �?      @      2@      $@      ;@      E@      D@      7@      ;@      @       @     �H@      �?      5@              &@      $@      <@      @      (@              �?      *@      @      3@      7@      =@      4@      &@      @      @      $@      $@      2@              0@      �?      4@      @      $@      �?      @      @      @       @      3@      &@      @      H@     �K@      F@      P@      &@     �S@      @     �Q@      0@      S@      >@      3@      (@     �@@     �G@      9@     @S@     �U@      T@      0@      C@     �C@     �A@     �H@       @      N@      @      L@      (@      H@      =@      0@      $@      9@      A@      ,@      L@     @P@     �D@      *@      9@      :@      3@      9@       @     �B@      @      6@      @      @@      ,@      @       @      @      4@      @      >@      <@      =@      "@      *@      *@      0@      8@      @      7@       @      A@      "@      0@      .@      (@       @      3@      ,@      @      :@     �B@      (@      @      $@      0@      "@      .@      @      2@              .@      @      <@      �?      @       @       @      *@      &@      5@      5@     �C@      @      $@       @      @      "@      @      ,@              @      @      2@              @      �?      @      $@       @      5@       @      5@      �?               @      @      @              @              "@              $@      �?              �?      @      @      @              *@      2@       @     �g@     �L@      B@     @f@      $@     �v@      @      \@      @      t@     �J@      5@      ,@      7@     �^@      3@     �j@     �e@     �r@     �H@     �b@     �F@      =@     `c@      @     0s@      @      U@      @     �p@      D@      ,@      &@      .@     @V@      (@     �e@     @a@     @p@     �A@      K@      .@      &@     @Y@       @     `f@             �F@             `c@      0@      $@      �?              F@      @     �W@     �Q@      f@      (@     �D@      @      @     �L@       @      ]@              B@             �_@      @       @      �?              ?@       @     �O@     �C@     �^@      @      *@      "@      @      F@             �O@              "@              <@      "@       @                      *@       @      ?@      ?@     �J@      @     �W@      >@      2@      K@      @      `@      @     �C@      @      \@      8@      @      $@      .@     �F@       @     @T@      Q@      U@      7@      S@      ;@      &@      I@      @      ]@              ?@      @     �Y@      2@      @      @      "@     �C@      @      Q@      M@      M@      7@      3@      @      @      @       @      (@      @       @              $@      @              @      @      @      �?      *@      $@      :@              E@      (@      @      7@      @      L@              <@      �?     �J@      *@      @      @       @     �@@      @      D@      A@      B@      ,@      ,@       @       @      @      @     �B@              &@              8@      &@      @              �?      0@      �?      (@      *@      0@      "@      ,@       @       @      @      �?     �B@              &@              6@      $@                      �?      "@              $@      *@      ,@      @                               @       @                                       @      �?      @                      @      �?       @               @      @      <@      $@      @      1@              3@              1@      �?      =@       @      @      @      @      1@      @      <@      5@      4@      @      @      @      @      @              &@              @      �?       @       @              @      @      "@              &@      @      @      �?      7@      @       @      &@               @              $@              ;@              @               @       @      @      1@      1@      1@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �3@��>U�@�	           ��@       	                    �?�)�ٴ�@           ܕ@                           �?E�r��v@            {@                            �?������@q            �e@������������������������       �P�1�d�
@            �C@������������������������       �	�͖@W            �`@                            �?/�ɶ��@�            Pp@������������������������       �'�M�@T            �_@������������������������       �י�]P�@T            �`@
                           @�'xI�@f           (�@                           �?z�)�c@�            �u@������������������������       ���N��@_            �a@������������������������       �m��P�f@|            `i@                           @�c�A/�
@�           h�@������������������������       �ߑ�}�
@�            `o@������������������������       �������
@�             w@                          @A@"l|��e@2           ��@                           @�X;S@           `�@                           �?������@�           p�@������������������������       ��\U��@�           �@������������������������       �+ʏ��@�           ��@                            �?���:jJ@T           ��@������������������������       �x�X�`@R            ``@������������������������       ���OK7�@           y@                           �?K�����	@             A@                             @����@z@             9@������������������������       ��swn`P@	             .@������������������������       ����N�@             $@������������������������       �u�&-�?             "@�t�bh�h5h8K ��h:��R�(KKKK��h��B        �t@     @\@     �X@     `u@     �C@      }@      @      m@      :@     p|@     @^@     �M@     �B@     @P@     @m@     @P@     w@     t@     0|@      T@     @Y@      8@      7@      b@      "@      k@       @      T@      @     �f@      >@      4@       @      @     �U@      .@     �^@     �\@     �h@      1@      >@      @      .@      L@      @     �M@       @      2@      @      B@      .@      $@              @      =@              >@     �F@      O@      @      .@      @      @      0@      @      @@              @              $@       @      �?                      *@              3@      ,@      :@       @              �?              @              @              @              @       @      �?                      @              @       @      @      �?      .@      @      @      *@      @      <@              @              @      @                              @              0@      (@      3@      �?      .@       @      (@      D@      @      ;@       @      &@      @      :@      @      "@              @      0@              &@      ?@      B@      @       @              @      ;@       @      $@              @      @      .@      @      @              @      @              @      &@      ,@       @      @       @      @      *@       @      1@       @      @              &@      @      @              �?      &@              @      4@      6@       @     �Q@      2@       @     @V@       @     �c@              O@             `b@      .@      $@       @      @     �L@      .@      W@     @Q@      a@      &@      7@      @       @      B@             �A@              5@             @P@      $@      @              �?      <@      (@      A@      :@      A@       @       @       @       @      $@              (@              ,@              =@      @      @                      (@      @      1@      .@      $@      @      5@       @              :@              7@              @              B@      @                      �?      0@      "@      1@      &@      8@      @      H@      ,@      @     �J@       @     �^@             �D@             �T@      @      @       @       @      =@      @      M@     �E@     �Y@      @      2@      @      �?      >@      �?      K@              &@              9@      @      @       @              (@      @      7@      (@      G@              >@       @      @      7@      �?      Q@              >@             �L@       @      �?               @      1@             �A@      ?@     �L@      @     �l@     @V@      S@     �h@      >@     @o@      @      c@      6@      q@     �V@     �C@     �A@      M@     �b@      I@     �n@     �i@     �o@     �O@     `l@     @U@     �Q@      h@      >@     @o@      @      c@      6@     �p@     @V@      B@      >@      M@     �b@      I@     �n@     �i@      o@     �O@     �c@     �Q@     �M@      b@      =@     `h@      @     �a@      3@     �j@      Q@      >@      :@      I@     �\@     �H@      g@      d@     �f@      K@     @U@      D@     �E@     �W@      4@      X@      @     �U@      .@     �^@     �D@      6@      0@      C@     �P@      8@     �^@     @W@     �Y@      9@      R@      ?@      0@      I@      "@     �X@             �J@      @     �V@      ;@       @      $@      (@     �G@      9@      O@     �P@     �S@      =@     �Q@      ,@      (@      H@      �?     �K@      �?      (@      @     �L@      5@      @      @       @      A@      �?      O@     �G@     �P@      "@      0@      @      "@       @              5@              @              "@      @      �?               @      @      �?      2@      @      0@              K@       @      @      D@      �?      A@      �?       @      @      H@      ,@      @      @      @      ;@              F@     �D@     �I@      "@      @      @      @      @                              �?               @       @      @      @                                              @              �?      @      @      @                              �?               @      �?      @      @                                                                      @       @      @                                                              @      @                                                              �?              @                                      �?               @      �?               @                                                              @                      �?                                                      �?                                                              @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�z1hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@��%S�@�	           ��@       	                   �1@9��8��@�           ޢ@                           �?7y̧@�           ��@                            @w��@1            �T@������������������������       ��Ls��@             �H@������������������������       ��aUݢ�	@             A@                            @����@�            �@������������������������       ���:��
@)           P~@������������������������       ������@Y            �_@
                           @#���l3@G           ��@                           �?ݝ��@K           ��@������������������������       ��v��˾@�           8�@������������������������       ��I(�4@�           H�@                           @�D�t[�@�            �x@������������������������       ������V@�            �j@������������������������       ��
��t�
@o            `f@                          �?@,�����@�           h�@                            @�{�s�@Z           D�@                           @- `�`�@J           ��@������������������������       ���u�@           �z@������������������������       ��-���@F           `�@                           @�u��L@           �y@������������������������       �sOS�;k@�            �u@������������������������       ��P%U��
@.            @P@                           @Z�LV@_             a@                           �?=��"�X@+             N@������������������������       �����@             >@������������������������       �<�%ŭ
@             >@                           �?U���1@4            @S@������������������������       �6�yFt�@)            �M@������������������������       ��xb嫯@             2@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@      a@     �X@     �u@     �H@     P|@      @     @m@      >@     �{@     @W@     �K@     �A@     �P@     `n@     @Q@     pw@     �r@     �}@     @S@     @g@      P@     �G@     �k@      7@     @v@       @      a@      .@     �q@      G@      A@      .@      <@     `a@      B@     �n@     @g@     s@      E@      F@      $@      $@     �J@      @     �\@       @      B@      �?     �Y@       @      @      �?      @      A@      @     �Q@      L@     �\@      ,@      @              @      @       @      "@              �?      �?      @      @      �?              @      @      �?              "@      6@              @              �?      �?       @      "@              �?      �?       @      �?                      �?       @                      @      1@              �?              @      @                                              @       @      �?              @      @      �?              @      @             �B@      $@      @      G@      @     �Z@       @     �A@             @X@      @      @      �?       @      =@      @     �Q@     �G@      W@      ,@      5@      @       @      C@       @     �S@              8@              S@      @      @      �?      �?      8@      @     �M@     �E@     �U@      "@      0@      @      @       @       @      ;@       @      &@              5@      �?      �?              �?      @              &@      @      @      @     �a@      K@     �B@     @e@      1@      n@              Y@      ,@      g@      C@      =@      ,@      5@     @Z@      >@     �e@     @`@     �g@      <@      \@     �@@      <@      c@      0@     �f@             @R@      @      c@      8@      4@      "@      .@     @T@      2@     @`@      W@      d@      ;@     �J@      6@      &@     @Q@      @     �X@             �A@       @     �T@      @      @       @      *@      A@      �?     �M@     �@@      R@      (@     �M@      &@      1@     �T@      *@     @T@              C@      @     @Q@      2@      ,@      @       @     �G@      1@     �Q@     �M@      V@      .@      >@      5@      "@      2@      �?     �N@              ;@       @      @@      ,@      "@      @      @      8@      (@     �F@      C@      ?@      �?      4@      ,@      "@      "@      �?      $@              .@      @      3@      (@       @      �?      @      1@      &@      5@      6@      .@              $@      @              "@             �I@              (@      @      *@       @      �?      @              @      �?      8@      0@      0@      �?      b@     @R@      J@      _@      :@     @X@      @     �X@      .@      c@     �G@      5@      4@     �C@      Z@     �@@     @`@     �\@     �d@     �A@     @`@     �K@     �D@     �\@      6@     �V@      @     �W@      .@     �b@     �E@      5@      *@     �@@      Y@      ;@     �]@     �X@     �c@      ?@     �W@      C@      6@      V@      ,@      R@       @      K@      @     �[@      <@      "@      $@      .@     �Q@      1@      U@     @R@     �^@      4@      G@      &@      (@      >@      �?      ?@      �?      9@              O@      0@       @      @              ?@      @     �C@      A@     �M@      @     �H@      ;@      $@      M@      *@     �D@      �?      =@      @     �H@      (@      �?      @      .@      D@      $@     �F@     �C@     �O@      .@     �A@      1@      3@      :@       @      3@      @      D@      &@     �C@      .@      (@      @      2@      =@      $@     �A@      :@      B@      &@      <@      0@      3@      6@      @      3@      @      C@      &@      6@      *@      (@       @      1@      4@       @      =@      7@      <@      $@      @      �?              @      �?                       @              1@       @              �?      �?      "@       @      @      @       @      �?      ,@      2@      &@      $@      @      @              @              @      @              @      @      @      @      &@      0@      "@      @       @      $@       @      @      @      @              @               @                      �?      @      @      @      @      @      �?              �?      @      @      @      @      @                              �?                              @                      �?       @                      �?      @      �?                       @              @              �?                      �?      �?      @      @      @      �?      �?              (@       @      @      @              �?              �?              �?      @              @      �?              @      @      *@       @      @      @       @      @      @              �?              �?              �?      @              @                      �?      @      $@      @       @      @                                                                              �?                      �?               @      �?      @       @       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJx��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @��<�@�	           ��@       	                   �3@�M#�'@�           6�@                           �?w(��@�           `�@                           @�e�W�@�            �p@������������������������       ���C��@�            �j@������������������������       ����v4@             M@                           �?��V�%@�           P�@������������������������       ��]��|7
@�            �w@������������������������       �.H�8;@�            �x@
                           �?���Ȳ@b           �@                            �?yZ��i8@�           ��@������������������������       ���ޚ�@�            @n@������������������������       ����Eb)@           0z@                           @����7@�           ��@������������������������       �6/���J@T           8�@������������������������       �����@g            �d@                           @�	���@�           ��@                           �? o_"C�@�           ȃ@                          �9@�ڿ�B@�            �w@������������������������       ���N�@�            `r@������������������������       � o>�j3@;             V@                           �?�n�c�.@�            `o@������������������������       �ݩ�m�@S            �`@������������������������       �W�5��@N            @]@                          �7@d�V,@           P{@                           �?TV	���@�            �p@������������������������       ������@K            �Y@������������������������       �a�o@d            �d@                          �8@����{@j            `e@������������������������       �ݩ��V@             9@������������������������       �,4=�>�@[            @b@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       0u@     �`@     �R@     �v@      E@     }@       @     @k@     �A@     �z@     @W@      J@      G@      K@     �n@      V@     �v@     �r@     �}@     �V@      l@     �X@     �D@     0r@      9@     �v@      @     �a@      8@     pt@      L@      @@      >@     �@@     �f@     �L@     Pp@      k@     0w@     �O@      J@      5@      $@     �^@       @     �d@             �I@      @     �`@      (@      ,@      @      @     �O@      $@     @\@      O@     �f@      3@      4@      @      @     �F@      �?      <@              *@      @      4@      �?       @      �?      @      (@      @      0@      3@     �L@       @      ,@      @      �?     �B@      �?      5@              @      @      3@      �?      @      �?      @      &@      �?      0@      *@     �D@       @      @               @       @              @              @              �?              �?                      �?      @              @      0@              @@      .@      @     �S@      �?      a@              C@             �\@      &@      @      @      �?     �I@      @     @X@     �E@      _@      &@      @      @       @      ?@      �?     @R@              :@             �J@      �?      @      �?      �?      :@             �I@      4@     @Q@       @      9@       @      @     �G@              P@              (@              O@      $@              @              9@      @      G@      7@     �K@      @     �e@     @S@      ?@      e@      7@      i@      @     �V@      5@      h@      F@      2@      8@      ;@     �]@     �G@     �b@     @c@     �g@      F@     �N@      7@      ,@      H@      @     @U@      �?     �B@              S@      5@      "@      $@      @     �D@      @      M@      M@      T@      4@      7@      @      "@      2@      @      :@      �?      9@              :@      @      �?      @      @      1@      @      &@      .@      ?@      @      C@      1@      @      >@             �M@              (@              I@      ,@       @      @      @      8@      @     �G@     �E@     �H@      *@      \@      K@      1@      ^@      1@      ]@      @     �J@      5@      ]@      7@      "@      ,@      5@     @S@      D@     �V@      X@     �[@      8@      X@      E@      1@     �\@      ,@     �X@      @     �D@      5@     �Y@      5@      "@      &@      3@     �L@      A@     �R@     @R@     �W@      8@      0@      (@              @      @      2@              (@              *@       @              @       @      4@      @      0@      7@      .@             �\@     �B@      A@     @R@      1@     �X@      @     @S@      &@     �X@     �B@      4@      0@      5@     �P@      ?@      Y@     �U@     @Y@      <@      L@      1@      5@     �F@      *@     @P@      @     �G@      @      G@      :@      (@      @      ,@     �@@      0@      O@      I@      R@      7@      :@      "@      4@      9@      "@      >@      @      ;@      @      6@      3@       @      @      (@      5@      ,@     �F@     �A@     �A@      $@      8@      @      "@      3@      "@      >@      �?      1@      @      5@      .@      @      @      "@      .@       @     �B@      ;@      8@      $@       @      @      &@      @                       @      $@       @      �?      @       @      �?      @      @      @       @       @      &@              >@       @      �?      4@      @     �A@              4@              8@      @      @               @      (@       @      1@      .@     �B@      *@      *@              �?      &@       @      0@              *@              (@      �?      @                      @      �?      @      $@      <@      "@      1@       @              "@       @      3@              @              (@      @                       @      @      �?      $@      @      "@      @      M@      4@      *@      <@      @      A@              >@      @     �J@      &@       @      $@      @     �@@      .@      C@      B@      =@      @     �@@      ,@      "@      3@       @      ;@              (@             �C@       @      @      @      �?      2@      *@      5@      9@      2@      �?      .@       @      @      @              .@              @              1@      @      �?                      @      �?      @       @      &@      �?      2@      (@      @      *@       @      (@              @              6@      @       @      @      �?      *@      (@      .@      1@      @              9@      @      @      "@       @      @              2@      @      ,@      @      @      @      @      .@       @      1@      &@      &@      @       @       @              �?                                      @      @                      �?       @                      @                      @      7@      @      @       @       @      @              2@      �?      @      @      @      @      @      .@       @      ,@      &@      &@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ&:�/hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @��4p��@�	           ��@       	                    @.�3��5@�           8�@                          �:@�K���@*           $�@                           @�<�Ґ@            �@������������������������       �fҭ�Lv@<           L�@������������������������       �����X@C            @[@                           �?�`��|@�            �p@������������������������       �C;��i�@9            @T@������������������������       �9_��'@r             g@
                          �2@>!fٚ�@�           L�@                          �1@�ƥ��	@�            0y@������������������������       �F�B;
@�            �n@������������������������       ���~kџ@a            �c@                           @��̨��@�            �@������������������������       ����@�            �i@������������������������       ��/�yNS@           {@                          �3@u���@�           ��@                           @�	�'��@�            pw@                           @7`��@�            @o@������������������������       ��$
�8�
@z             g@������������������������       ���,
�@%            @P@                           �?�j�V!|@P            @_@������������������������       ���o�G@#            �L@������������������������       ���v6�o@-             Q@                          �:@��R3@�           ��@                           �?��RB�@n           �@������������������������       �ۑ���@�            �l@������������������������       �!u(I(@�            �w@                          �;@��.^!@            �j@������������������������       �n,s�7@-            @S@������������������������       ���c�4@R             a@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       Ps@     �_@     �U@     �w@     �G@     �}@      $@     `k@      4@     0z@     �\@      O@     �H@      Q@     @k@     @Q@     0w@     �r@     p}@     @Y@     `i@      U@      K@     q@      5@     �v@      @     �_@      .@     �s@     �O@      D@     �A@      C@      c@     �D@     �p@     �i@     �u@     �N@      ^@     �M@      E@     �f@      1@     `f@      @      S@      @     �f@     �F@      ?@      8@      @@     �Y@     �A@     �e@      `@     �g@     �E@     @Z@      H@     �B@     @c@      1@     �c@      @     �J@      @      d@     �@@      <@      @      7@      U@      >@     �b@     �[@     �d@      B@     �W@     �B@      B@     �b@      &@     `b@      @      J@      @      c@      ;@      <@      @      7@      T@      8@     ``@     @Y@      c@      B@      $@      &@      �?      @      @      &@              �?              @      @                              @      @      2@      $@      *@              .@      &@      @      <@              5@      �?      7@      �?      6@      (@      @      1@      "@      3@      @      7@      2@      9@      @      &@              @       @              @      �?       @      �?      @      @              @      @      @      @       @      @      @      �?      @      &@      �?      :@              0@              .@              .@       @      @      (@      @      .@      �?      .@      *@      3@      @     �T@      9@      (@     �V@      @     �f@             �I@      $@     �`@      2@      "@      &@      @     �H@      @     �X@     @S@     �c@      2@      3@      @      @      9@      �?      U@              9@              Q@       @       @      @              .@             �@@      <@     �T@      @      "@      @      @      ,@      �?     �L@              (@             �A@      �?       @       @              (@              .@      5@     �G@      @      $@                      &@              ;@              *@             �@@      �?              �?              @              2@      @     �A@              P@      2@       @     �P@      @     �X@              :@      $@     �P@      0@      @       @      @      A@      @     �P@     �H@     �R@      *@      .@      @              7@              @@              "@       @      :@      @       @      �?      �?      &@      @      (@      5@      =@      @     �H@      .@       @     �E@      @     �P@              1@       @      D@      *@      @      @      @      7@              K@      <@      G@       @     �Z@     �E@     �@@      Z@      :@      \@      @      W@      @     �Y@     �I@      6@      ,@      >@     �P@      <@      Y@     �W@      _@      D@      ;@      @      @     �A@       @     �L@              9@             �D@      6@      @      �?       @      1@       @     �C@      6@      L@      @      0@              @      2@      �?      E@              4@              9@      1@              �?       @      (@      @      @@      *@     �D@      @      ,@               @      .@              ?@              2@              1@      0@              �?      �?      "@      �?      2@       @     �@@      �?       @              �?      @      �?      &@               @               @      �?                      �?      @      @      ,@      @       @       @      &@      @      @      1@      �?      .@              @              0@      @      @                      @      @      @      "@      .@       @      @      �?              *@      �?      @              �?              @      @      @                       @              @       @       @       @      @      @      @      @               @              @              *@      �?       @                      @      @      @      �?      *@             �S@     �C@      ;@     @Q@      8@     �K@      @     �P@      @      O@      =@      0@      *@      <@     �H@      4@     �N@     @R@      Q@     �A@      N@      <@      0@      C@      2@      J@             �I@      @     �H@      7@      $@      &@      9@     �@@      (@      J@     �J@     �D@     �@@     �@@      "@      $@      ,@      @      .@              4@       @      1@       @      @              @      (@      @      *@      5@      <@       @      ;@      3@      @      8@      &@     �B@              ?@       @      @@      .@      @      &@      6@      5@      @     �C@      @@      *@      9@      3@      &@      &@      ?@      @      @      @      0@      �?      *@      @      @       @      @      0@       @      "@      4@      ;@       @      @              @      "@      @      @      @      @      �?      @              @                      @      @      @      @      .@              (@      &@      @      6@      @                      $@              "@      @       @       @      @      *@      @      @      *@      (@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJʺ-ghG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@�� ��@�	           ��@       	                     @r��J��@r           �@                            �?�^-v2�@�           Џ@                           @~f��@           X�@������������������������       ���ʁ�@!           `}@������������������������       ��"*3)T
@�            Pu@                          �0@���8�I
@�            �i@������������������������       �/.\&�@             C@������������������������       �j�\cg
@o             e@
                          �1@ٴ���\@�            �x@                           �?��1@b            �c@������������������������       ���v��R	@%             L@������������������������       �-�!+d@=            �Y@                           @8՛��@�             m@������������������������       �s7D�r�
@T            �a@������������������������       �1�N5
@2            �V@                           @���[@           ��@                           @�R�b�?@G           ��@                           @iI��eu@f           ��@������������������������       ��霛�{@R           L�@������������������������       �x�4�@             E@                          �>@�����0@�            �v@������������������������       ����@�            �t@������������������������       �'>�N@             <@                           �?� r@�            �@                           @{H0�@�            �t@������������������������       ����y
@             E@������������������������       �[/����@�            0r@                           @�^��R@�            0y@������������������������       �1�S�@�            `o@������������������������       �9�ob@^             c@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       0u@     ``@     �Y@     �u@      H@     P@      @     �i@      ;@     �z@     �[@      I@     �D@      O@     �k@     �N@     �x@     �s@     �{@     �S@     �V@      B@      B@     @c@      $@     �l@      �?     �O@       @     �d@      9@      3@      "@      @      K@      .@      b@     �\@     �k@      2@      I@      6@      .@     �^@      @      e@              C@       @     ``@      ,@      2@       @      @     �E@       @     �W@      T@      g@      &@      B@      2@      *@     �Z@       @     @\@              >@       @     �Y@      *@      &@      @      @      B@       @      S@     �Q@     @c@      $@      3@      @      *@     �S@      �?      J@              "@       @      L@      &@       @      @      @      8@      @      H@      A@     �U@       @      1@      &@              <@      �?     �N@              5@             �G@       @      @       @              (@       @      <@     �B@     �P@       @      ,@      @       @      0@      �?      L@               @              <@      �?      @      @      �?      @              2@      "@      ?@      �?                       @       @              ,@                              @                              �?       @              @              @              ,@      @              ,@      �?      E@               @              6@      �?      @      @              @              (@      "@      :@      �?      D@      ,@      5@      ?@      @     �M@      �?      9@              A@      &@      �?      �?              &@      @     �I@      A@     �B@      @      *@      "@      @      3@      @      6@      �?      @              7@      @      �?                      @      �?      5@       @       @      @      @               @      @      @      0@              �?               @                                       @      �?      @      @              @       @      "@      @      0@       @      @      �?      @              .@      @      �?                      �?              0@      @       @       @      ;@      @      0@      (@       @     �B@              2@              &@      @              �?               @      @      >@      :@      =@              $@      @      0@      @       @      :@              @              @       @              �?              @      �?      <@      0@      .@              1@      �?              @              &@              &@               @      @                              @      @       @      $@      ,@              o@     �W@     �P@      h@      C@     q@      @     �a@      9@     Pp@     @U@      ?@      @@      M@      e@      G@     �o@     �h@     �k@     �N@      g@     �K@      J@      b@      7@      m@      @     @X@      3@     �d@     @P@      6@      7@      B@     �\@      @@     �d@      a@      c@      F@     �`@      D@      A@      `@      4@     �e@      @      V@      3@     �`@      M@      0@      0@      ?@     �V@      @@     �^@     @\@     �[@      D@     ``@      D@      A@     �_@      4@     @d@      @     �U@      *@      `@      M@      0@      0@      ?@     �V@      @@     �^@     �Z@      Z@      D@      @                      @              (@              �?      @      @                                                      �?      @      @             �I@      .@      2@      .@      @      M@      �?      "@              @@      @      @      @      @      7@              E@      8@      E@      @     �I@      *@      (@      .@      @      K@              "@              >@      @      @      @      @      7@              >@      8@     �D@      @               @      @                      @      �?                       @                                                      (@              �?              P@      D@      ,@     �H@      .@     �D@             �F@      @     @X@      4@      "@      "@      6@      K@      ,@      V@      O@     �Q@      1@      4@      4@      $@      2@      $@      ,@              ;@      �?     �I@      @      @      @      5@      :@      (@      A@      4@      >@      "@      �?       @              �?                               @                      �?                      @       @      @      @      @      @      @      3@      2@      $@      1@      $@      ,@              3@      �?     �I@       @      @      @      1@      8@      @      <@      .@      ;@      @      F@      4@      @      ?@      @      ;@              2@      @      G@      1@      @      @      �?      <@       @      K@      E@      D@       @      >@      (@      @      .@      @      4@              .@      @      A@      &@      @      @              1@      �?      ;@      *@      ?@      @      ,@       @              0@      �?      @              @              (@      @      @       @      �?      &@      �?      ;@      =@      "@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ7�@hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @%�"�y@�	           ��@       	                    �?r�F�Z�@�           �@                          �3@�\��X�@�           �@                           @��2��
@           P{@������������������������       ����e�@�            �j@������������������������       ������@�             l@                           �?;�9QA@�           8�@������������������������       ��e��1:@�            �m@������������������������       �*r0��@            �y@
                           �?�o0�@7           �@                          �5@��I��@�           ��@������������������������       �S�"4G�@�            �w@������������������������       ��*e�5�@�            �u@                          �6@,�����@z           �@������������������������       ���o�K@r           ȁ@������������������������       �� ��V�@           �z@                           @�[�>YL@�           L�@                           �?Gt.���@@           P�@                           �?�Ү{@�            �s@������������������������       ���rB�@0             R@������������������������       ����O�@�             n@                           �?ޑ�؀@�            @j@������������������������       ��~�3�t@i             e@������������������������       ����0c	@            �D@                           �?���Xd|@}           H�@                          �7@TXx�M�@�             x@������������������������       ���c��@�            �j@������������������������       �\ �@�@k            �e@                          �9@���õ'@�            �h@������������������������       ��F�Tv@}            �e@������������������������       ��+w1F&@             9@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       u@     �b@     �T@     �u@      @@     �@      @     �m@      >@     �{@     �Z@     �L@     �@@      L@      m@     �J@      v@     �u@     �y@     �T@     �l@     �Z@     �F@     Pp@      0@     �x@      @      d@      1@     Pu@     @P@     �B@      :@      @@     �e@     �@@     �o@     �k@     Pt@      P@      S@      :@      0@     �V@       @     �h@      �?     �M@      @     @c@      >@      *@      "@      "@      M@              Z@     @V@     �_@      6@      4@      @      @     �@@      �?     �X@              8@      @     �S@      @      $@              �?      8@              A@      ?@      O@      @       @      @      @      4@              A@              @       @     �D@      @      $@              �?      0@              4@      *@      :@       @      (@                      *@      �?      P@              2@       @     �B@                                       @              ,@      2@      B@      �?      L@      5@      (@     �L@      �?     �X@      �?     �A@              S@      9@      @      "@       @      A@             �Q@      M@      P@      3@      1@      &@      @      9@      �?      A@      �?      1@              =@      &@       @      "@      @      &@              :@      .@      &@       @     �C@      $@      @      @@              P@              2@             �G@      ,@      �?              @      7@              F@     �E@     �J@      &@     @c@      T@      =@     `e@      ,@      i@      @     �Y@      *@     `g@     �A@      8@      1@      7@     �\@     �@@     �b@     ``@     �h@      E@     �Q@      =@      @     �R@      $@     �Z@      @     �D@      @     @R@      $@      @      &@       @     �J@      .@     �P@     �F@     �U@      .@      ,@      4@      @     �C@      @      P@              ;@             �A@      @      @      @      �?      :@      @     �C@     �@@      K@      @     �L@      "@      @     �A@      @      E@      @      ,@      @      C@      @              @      �?      ;@      $@      ;@      (@      @@      "@     �T@     �I@      6@     @X@      @     �W@             �N@      @     �\@      9@      4@      @      5@     �N@      2@     @U@     �U@     @\@      ;@      H@      .@      ,@     �K@      �?     �O@             �B@      @     @R@      ,@      ,@      @      @      ?@       @      H@     �K@     �N@      .@     �A@      B@       @      E@      @      ?@              8@             �D@      &@      @       @      .@      >@      $@     �B@      ?@      J@      (@     �Z@     �F@      C@     @V@      0@     �\@       @     @S@      *@     �Z@      E@      4@      @      8@     �N@      4@     @X@     �_@      U@      2@     �I@      :@      &@     �B@       @      M@      �?     �H@      @     �F@      8@      $@              ,@      <@      $@      E@     �O@      D@       @      =@      $@      "@      4@       @      =@      �?      @@      @      :@      0@      @              &@      (@       @     �@@     �F@      2@      �?      $@      @       @       @              @      �?      @       @      @      @      @               @       @       @      @       @      @              3@      @      @      (@       @      6@              ;@      �?      6@      $@      @              "@      $@      @      >@     �B@      ,@      �?      6@      0@       @      1@              =@              1@              3@       @      @              @      0@       @      "@      2@      6@      @      3@      @       @      *@              :@              *@              &@      @      @              @      0@       @      @      .@      3@      @      @      "@              @              @              @               @      �?                                               @      @      @      �?      L@      3@      ;@      J@      ,@      L@      �?      <@      $@     �N@      2@      $@      @      $@     �@@      $@     �K@      P@      F@      $@     �B@      &@      4@      ;@      ,@      ?@      �?      3@      "@      A@      1@      "@      @       @      7@       @     �B@     �F@      <@       @      3@      @      "@      .@      ,@      6@              @      �?      6@      (@      @      �?               @              6@      <@      4@      @      2@      @      &@      (@              "@      �?      (@       @      (@      @      @      @       @      .@       @      .@      1@       @      @      3@       @      @      9@              9@              "@      �?      ;@      �?      �?      �?       @      $@       @      2@      3@      0@       @      2@       @      @      9@              3@              @      �?      :@      �?      �?                       @       @      *@      3@      *@       @      �?              �?                      @              @              �?                      �?       @       @              @              @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�n/hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�3�Ft�@�	           ��@       	                   �4@E��-��@�           �@                           �?��Nd�@^           �@                          �2@��#,_@h           P�@������������������������       �
ЍR�F@�            �r@������������������������       �C�}	�@�            �q@                           �?���	�@�           Ē@������������������������       �m=��SS@/           @~@������������������������       �atѝ3�@�           h�@
                            �?���Ɇ�@�           ��@                           �?���0@�            v@������������������������       �'7�f@Z            �a@������������������������       �ĵ���@�            `j@                           @�jfeQn@�            pq@������������������������       �"�ʏ��@w            �h@������������������������       �1����@4            @T@                           @����@�           X�@                            @��D�@�           �@                           �?$�
}C@�           ��@������������������������       �k|��{@�            ps@������������������������       ������@0           �@                           �?�u�Ic@           `x@������������������������       �[O%2�@(             N@������������������������       ��ni��B@�            �t@                           @C��
+@�            �q@                            �?u�O9�
@D            @[@������������������������       ��i�H�_@             8@������������������������       �nM�l
@2            @U@                           �?���r1$@q            �e@������������������������       �>+���-@1            �R@������������������������       ��l�@�@@            �X@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     @c@      V@     v@      B@     `{@      "@     �m@      <@     }@     @Z@     �M@      ;@     �R@     �l@     �P@     �u@     pt@     `|@      W@     �h@     �U@      G@     �k@      0@      s@      @     `a@      &@     s@     �F@      F@      ,@      @@      _@      <@     �m@     `j@     `s@      E@     �`@      F@      C@     �c@      $@     �k@       @      Y@      "@      m@      A@      A@      (@      1@     @W@      8@     `d@     �d@     0p@     �A@     �K@      (@      8@     �J@       @     �J@       @      =@       @     �I@      0@      4@      @      "@     �C@      @      F@      M@     @T@      .@      :@      @      &@     �A@      @      @@       @      .@      �?      5@       @      $@      �?      @      6@      @      .@      B@      F@      @      =@      @      *@      2@       @      5@              ,@      @      >@       @      $@       @      @      1@      �?      =@      6@     �B@      (@     �S@      @@      ,@      Z@       @     @e@             �Q@      �?     �f@      2@      ,@      "@       @      K@      2@     �]@     @[@     @f@      4@     �@@       @      �?      @@      �?     �S@              A@             @S@      $@      �?              @      1@      @      H@      I@     @R@      &@      G@      8@      *@      R@      �?      W@             �B@      �?      Z@       @      *@      "@      �?     �B@      .@     �Q@     �M@     @Z@      "@      O@      E@       @     �P@      @     �T@      �?     �C@       @     @R@      &@      $@       @      .@      ?@      @     �R@      F@     �I@      @     �C@      >@      @      G@       @     �E@      �?      5@      �?      :@      @      @       @      @      .@      @      F@      3@     �D@       @      3@      *@              "@              5@      �?      @              @      @              �?      @      @              :@      $@      1@       @      4@      1@      @     �B@       @      6@              ,@      �?      5@              @      �?      @      $@      @      2@      "@      8@              7@      (@      @      4@      @      D@              2@      �?     �G@       @      @               @      0@      �?      ?@      9@      $@      @      2@      &@      @       @      @      7@              .@              E@      @       @              @      @      �?      9@      7@      �?      �?      @      �?      �?      (@              1@              @      �?      @      �?      @               @      "@              @       @      "@      @     �`@      Q@      E@     @`@      4@     �`@      @     @X@      1@      d@      N@      .@      *@      E@      Z@      C@      [@      ]@      b@      I@     @V@      L@      C@     �Z@      3@      Z@      @     �V@      0@     �_@      K@      ,@      (@      @@     @U@     �A@     @U@     @W@     �Z@      G@     �M@      G@      .@      R@      $@      T@      �?     �K@       @     �Y@     �A@      "@      "@      ,@     �N@      :@     �K@      O@     @S@      @@      ;@      @       @      7@      @      :@      �?      6@       @      E@      $@              �?      @      ?@      &@      9@      =@      8@      0@      @@     �E@      @     �H@      @      K@             �@@              N@      9@      "@       @      &@      >@      .@      >@     �@@     �J@      0@      >@      $@      7@      A@      "@      8@      @      B@      ,@      8@      3@      @      @      2@      8@      "@      >@      ?@      =@      ,@      @      �?      @      @       @      @      @      @      �?       @      @                              @              $@      �?      @      @      7@      "@      2@      =@      @      4@              @@      *@      6@      0@      @      @      2@      3@      "@      4@      >@      :@      &@     �E@      (@      @      8@      �?      <@      �?      @      �?      A@      @      �?      �?      $@      3@      @      7@      7@      C@      @      5@       @              @      �?      ,@                      �?      $@       @      �?               @      $@              @      @      6@      @      @                       @              @                              @      �?                       @       @              �?                              ,@       @              @      �?       @                      �?      @      �?      �?                       @              @      @      6@      @      6@      $@      @      2@              ,@      �?      @              8@      @              �?       @      "@      @      1@      0@      0@               @       @       @      @               @      �?      @              (@      �?                              @      @      @      $@      @              ,@       @       @      (@              @              �?              (@      @              �?       @      @              $@      @      &@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ���YhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@���Ӆ�@�	           ��@       	                    �?܎�vk@�           Ƣ@                            �?�S{Hm�@�           ��@                          �4@5~r�D@�            �m@������������������������       ���b��@e            �c@������������������������       �&!Э�@0            @T@                           �?e���@b           8�@������������������������       ��^��@�            �i@������������������������       �;���F@�            �s@
                           @�<��@�           ��@                          �5@��6@           ��@������������������������       �;f�$@�           ��@������������������������       ����2�=
@N             ^@                          �2@��#�2b@�            �x@������������������������       ���$I@h             f@������������������������       �B�Lt@~            `k@                           �?)�`9ݵ@�           ��@                           @��p�@�           �@                           �?%���O@           @z@������������������������       ��#�F@�            @n@������������������������       ����=%�@o            @f@                           �?�m��"@y            �g@������������������������       ���:�"W	@.            @T@������������������������       �E�`�k�@K            �[@                           @��ٮ��@<           �@                           �?'�O@�           ��@������������������������       ��>5�_@�             l@������������������������       ��P]�@X           ��@                           @|$�{�1@b            @b@������������������������       � i���
@             C@������������������������       ��O�*-<@E             [@�t�b��     h�h5h8K ��h:��R�(KKKK��h��B`       �t@     `a@     @\@      u@      ?@     0�@      @     �n@      :@     �|@      Y@      N@      :@     �Q@      m@      N@      v@     @q@     �{@     �S@     �g@      M@      K@      k@      3@     pw@      �?     `b@      $@     @s@      L@      C@      @      ;@      `@      =@     �k@     �c@     �s@      F@     �O@      4@      =@     �R@      (@     �V@      �?      L@      @     �U@      3@      *@      �?      5@     �C@      $@      O@      M@     �S@      0@      0@       @      $@     �A@              5@              6@      @      =@      �?      @              @      0@      @      (@      3@      @@      @      "@              $@      5@              2@              *@              4@      �?      �?              �?      .@       @      @      ,@      6@      @      @       @              ,@              @              "@      @      "@               @              @      �?      @      @      @      $@      �?     �G@      2@      3@      D@      (@     �Q@      �?      A@      @     �L@      2@      $@      �?      .@      7@      @      I@     �C@     �G@      "@      4@       @      @      ,@      @      A@              &@              1@      "@      @              @      @      @      8@      1@      ;@              ;@      0@      ,@      :@      @      B@      �?      7@      @      D@      "@      @      �?      (@      0@      �?      :@      6@      4@      "@     �_@      C@      9@     �a@      @     �q@             �V@      @     �k@     �B@      9@      @      @     �V@      3@      d@      Y@     `m@      <@     @U@      5@      1@     @^@      @     @m@             �P@              e@      6@      9@      @      @      O@      2@     �_@     �Q@     �e@      9@      R@      5@      .@     @]@      @     @i@             �O@             �b@      3@      8@      @      @     �H@      2@      ]@     @P@     �d@      5@      *@               @      @      @      @@              @              2@      @      �?                      *@              &@      @      @      @      E@      1@       @      5@              I@              8@      @     �J@      .@              �?      @      <@      �?      A@      >@     �O@      @      "@      $@      @      @              2@              1@              C@       @              �?      @      "@      �?      (@      ,@      @@      @     �@@      @      @      1@              @@              @      @      .@      *@                              3@              6@      0@      ?@              b@     @T@     �M@     �]@      (@     �a@      @      Y@      0@     �b@      F@      6@      4@      F@      Z@      ?@     ``@     �]@     @`@      A@     �R@      9@      5@     �G@       @      O@      @      D@      (@     @S@      *@      @      @      "@      E@      @     �K@      F@      H@      ,@      E@      6@      3@      6@      @      E@      �?      A@       @     �K@      $@      @      @      "@     �@@       @     �A@      <@      <@      ,@      2@      "@      2@      .@      @      0@      �?      4@      @      @@       @      @      @      @      3@              7@      4@      2@      @      8@      *@      �?      @       @      :@              ,@      @      7@       @      �?      �?      @      ,@       @      (@       @      $@      "@     �@@      @       @      9@       @      4@       @      @      @      6@      @       @                      "@       @      4@      0@      4@              &@               @      @              @              @              0@                                      @      �?      $@      @      ,@              6@      @              2@       @      ,@       @      �?      @      @      @       @                      @      �?      $@      &@      @             �Q@      L@      C@      R@      @     @T@      @      N@      @     �R@      ?@      0@      ,@     �A@      O@      ;@      S@     �R@     �T@      4@      J@      H@      >@     �P@      @     �Q@      @     �M@      @      N@      <@      0@      (@      <@      H@      :@     �L@     @P@      O@      .@      "@      @      @      3@              5@              5@      �?      6@      *@      @      @      @      5@      &@      1@       @      6@      $@     �E@     �D@      7@     �G@      @     �H@      @      C@      @      C@      .@      &@      @      9@      ;@      .@      D@     �L@      D@      @      2@       @       @      @              &@              �?              ,@      @               @      @      ,@      �?      3@      "@      4@      @      @      @      �?      �?              @                              @       @                              @              @      @      "@       @      ,@      @      @      @               @              �?              &@      �?               @      @      &@      �?      .@      @      &@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ1P�ShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?
�{-��@�	           ��@       	                   �<@LE���@$           4�@                          �4@��[�s�@�           �@                           @�nԩ��@w           ��@������������������������       ��$Ї��@)           P}@������������������������       �����@N            �`@                           @^o���@0           8�@������������������������       �WǕ�Az@�           @�@������������������������       �u|�KO@:            �W@
                           @��3@}            @i@                          �>@�K�*]@l            �e@������������������������       �Kd��@-            @P@������������������������       ���	�'�@?             [@                            @�'�@P�@             =@������������������������       ���1�@
             1@������������������������       �Z��h W@             (@                          �2@���R|i@~           x�@                           @uV��M@�           H�@                            @o�@Q             a@������������������������       ��ܷj'�	@9            �W@������������������������       �z�0�
@             E@                           @���2|@�           �@������������������������       ��x��
@!           �}@������������������������       �/��t�@c             e@                           @������@�           ̖@                          �;@�R�K�@�           Ȅ@������������������������       �G���M@�           ��@������������������������       �Y9X�� @1            �P@                           @�X��a�@�           Ј@������������������������       ��|�@           �y@������������������������       ��t�s��@�            �w@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       t@     @a@     @W@     �u@      D@     0@       @      m@      E@     �y@     @W@     @P@     �E@     @S@     `o@     �H@     �v@     �s@     @}@     �O@     �a@     @Q@     �O@     �b@      <@     `c@       @     �^@      ?@      `@      F@      A@      9@     �I@      Z@      3@      a@     `b@     �g@      >@     �]@     �G@     �G@      a@      ;@     �b@      @     �]@      =@     �\@     �@@      ?@      0@     �F@     @V@      .@     �_@     @_@     �e@      >@      J@      *@      4@     �N@      "@     �Q@      �?      B@      @     �H@      5@      *@      @      "@     �C@      @     �B@      J@     �V@      2@      @@      @      &@      J@      "@     �K@      �?      6@      @      E@      ,@      &@      @      "@      >@      @      A@      D@     @R@      *@      4@      @      "@      "@              .@              ,@              @      @       @                      "@              @      (@      1@      @     �P@      A@      ;@     �R@      2@     �S@      @     �T@      8@     @P@      (@      2@      $@      B@      I@      (@     @V@     @R@      U@      (@      K@      ;@      8@     �R@      ,@     �R@      @     @S@      5@      L@      (@      ,@       @      ?@      E@      @      T@      Q@      S@      $@      (@      @      @              @      @              @      @      "@              @       @      @       @      @      "@      @       @       @      8@      6@      0@      ,@      �?      @       @      @       @      .@      &@      @      "@      @      .@      @      $@      6@      .@              8@      4@      0@      "@      �?      @       @      @       @      .@       @      @      @      @      &@      @      @      3@      $@              "@      @      @      @              @       @                      "@      @       @      @      �?      $@               @      @      @              .@      1@      (@      @      �?       @              @       @      @      @      �?      @      @      �?      @      @      .@      @                       @              @               @                                      @               @              @              @      @      @                                       @               @                                                       @              @              @      �?      @                       @              @                                                      @                                                       @       @             `f@     @Q@      >@     @h@      (@     �u@             @[@      &@     �q@     �H@      ?@      2@      :@     `b@      >@      l@     @e@     pq@     �@@     �F@      0@      @     �R@      �?      `@              H@             @]@      $@      &@      @      $@      @@      (@      T@      L@     �\@      &@      $@      �?      �?      6@              4@              @              ,@      @                      @      @      @      "@      5@       @      @      @              �?      4@              *@              @              *@      @                      @                      @      0@      @      @      @      �?               @              @              �?              �?      @                              @      @      @      @      �?      �?     �A@      .@      @      J@      �?      [@             �E@             �Y@      @      &@      @      @      <@      @     �Q@     �A@     �Z@      @      ?@      @       @     �D@      �?     �U@              9@             @R@      @      $@       @       @      3@      @      K@      <@     �T@      @      @      $@      @      &@              6@              2@              >@              �?       @      @      "@       @      1@      @      9@       @     �`@     �J@      7@      ^@      &@      k@             �N@      &@     `d@     �C@      4@      ,@      0@     �\@      2@      b@     �\@     �d@      6@     �L@      @@      "@      J@      "@      X@              ?@             �S@      .@      (@      @      @     �J@      $@     @P@     �L@     �P@      "@     �H@      ?@       @      I@      @     �V@              >@             �Q@      (@      (@       @      @     �I@      @      N@      K@      M@      @       @      �?      �?       @      @      @              �?              "@      @              @      �?       @      @      @      @       @       @     @S@      5@      ,@      Q@       @      ^@              >@      &@      U@      8@       @      @      $@      O@       @      T@     �L@     �X@      *@      E@       @      @      C@             �S@              4@       @      E@      @      @      @      @     �A@      @      B@      =@      I@      @     �A@      3@      $@      >@       @     �D@              $@      @      E@      4@      @      @      @      ;@      @      F@      <@      H@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJa�5chG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@Ë�M�@�	           ��@       	                    @d)�VB�@�           ��@                           �?��$�h�@�           ��@                           �?�=˶�k@           �z@������������������������       ��9ym@u            �g@������������������������       ��RCn@�             n@                          �4@E��.@�           ��@������������������������       ��ž�.<@X           ��@������������������������       ��h�al@�            �m@
                           @'b-�@�           ��@                            �?�?0�:�@�            �p@������������������������       �f\s�I
@j             d@������������������������       ��.��
@B            @[@                           @A.�kP�@=           ��@������������������������       �J�d��@�           Ѕ@������������������������       �`�s��
@�            �l@                           �?2��k�@�           ��@                           @��I�'@�           ��@                            @�=r'@Y           ��@������������������������       ��vL]x�@�            �s@������������������������       �{iOW�
@�            `l@                           �?x�g���@�            p@������������������������       ����#��
@)            �Q@������������������������       ���PVT@r            @g@                          �9@(_�0@�           ��@                           @P���@�            @w@������������������������       ��d���@�            @i@������������������������       ��TY��1@s            @e@                           @[Jv++@�            �u@������������������������       �)���@�            �j@������������������������       �B�ɴ�@V             a@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       Pt@     �^@     �T@     @v@     �H@     `}@       @      n@      ?@      {@     @_@      Q@      =@     �O@     �m@      L@     �y@     �r@     p{@     �Q@     @f@     �O@      G@     �l@      9@     Pv@      �?      a@      .@     �q@      M@     �I@      &@      9@      ^@      6@     �o@     �f@     pr@     �C@     �[@     �@@      <@      ^@      6@      a@      �?     @Q@      $@     @]@     �F@      6@      @      4@      P@      0@     @^@     @Z@      _@      ;@     �E@      *@      @     �H@       @      I@              9@      @     �J@       @      @      �?       @      5@      �?      A@      @@     �N@       @      4@      �?              "@              7@              2@              <@      @      @      �?      �?      &@              ,@      4@      >@      @      7@      (@      @      D@       @      ;@              @      @      9@      @       @              @      $@      �?      4@      (@      ?@      @      Q@      4@      8@     �Q@      ,@     �U@      �?      F@      @      P@     �B@      .@      @      (@     �E@      .@     �U@     @R@     �O@      3@     �G@      &@      7@      J@      (@      F@              :@      @     �C@      ?@      *@      �?       @      >@      $@     �M@     �G@      L@      2@      5@      "@      �?      3@       @      E@      �?      2@      @      9@      @       @      @      @      *@      @      <@      :@      @      �?     �P@      >@      2@     @[@      @     �k@              Q@      @      e@      *@      =@      @      @      L@      @     ``@     �S@     `e@      (@      @       @      @      @@              D@              @              G@       @      "@      �?              (@      @     �A@      6@     �A@      @       @       @       @      5@              5@              @              =@                      �?              @      @      ;@      $@      5@      @      @               @      &@              3@              @              1@       @      "@                      @               @      (@      ,@       @      N@      6@      ,@     @S@      @     �f@             �N@      @     �^@      &@      4@      @      @      F@      �?      X@      L@      a@      @      G@      0@      *@      O@      @      ^@             �K@      �?     �Y@      $@      *@      @       @      ;@      �?     @Q@      C@     �[@      @      ,@      @      �?      .@             �N@              @      @      5@      �?      @              @      1@              ;@      2@      9@      @     `b@     �M@      B@     �_@      8@     @\@      @     �Y@      0@     �b@     �P@      1@      2@      C@     @]@      A@     �c@     �\@      b@      @@      J@     �C@      9@      R@      .@     �D@      @      R@      (@     �O@      C@      *@      *@      <@      O@      4@     �U@     �K@     �Q@      2@      C@      ;@      2@      J@      @      9@      @     �E@      &@      B@     �B@      $@       @      3@      H@      ,@     �N@     �C@     �A@      &@      ;@      3@      @      9@      @      0@      �?      ;@              >@      5@       @      @      @     �B@      @      A@      0@      9@      @      &@       @      *@      ;@              "@      @      0@      &@      @      0@       @      @      (@      &@      $@      ;@      7@      $@      @      ,@      (@      @      4@      $@      0@              =@      �?      ;@      �?      @      @      "@      ,@      @      9@      0@     �A@      @              @      @      @      @      $@              @              @                              �?      @              $@      @      0@      �?      ,@       @      @      ,@      @      @              7@      �?      7@      �?      @      @       @      $@      @      .@      *@      3@      @     �W@      4@      &@     �K@      "@      R@       @      ?@      @     @U@      =@      @      @      $@     �K@      ,@      R@      N@     �R@      ,@     �L@      *@      @      @@             �C@              "@             �J@      .@                      @     �A@       @     �B@     �C@      9@      @     �B@      $@      @      ,@              2@              @              9@      &@                      �?      4@      �?      8@      3@       @      @      4@      @      @      2@              5@               @              <@      @                      @      .@      �?      *@      4@      1@              C@      @      @      7@      "@     �@@       @      6@      @      @@      ,@      @      @      @      4@      (@     �A@      5@     �H@      $@      ,@      @       @      1@      @      8@              6@      @      4@       @      �?       @      @      @      &@      1@      ,@      <@       @      8@      @       @      @      @      "@       @                      (@      @      @      @       @      *@      �?      2@      @      5@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�WhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�W\K�@�	           ��@       	                    �?_f��pD@           �@                          �6@���D�@T           ��@                          �3@i��5�C@:            @������������������������       �{D�F@�            �p@������������������������       �GB��1@�             l@                          �?@_	ZV�@           |@������������������������       �9��@�            �y@������������������������       ����&�
@             D@
                           @����<R@�           �@                           @�uG��@~           ��@������������������������       �{	��Y\@�           ��@������������������������       ���1�Km@�             t@                            �?K�B��@/           �}@������������������������       ��p8B��@�            0v@������������������������       ���]��?@M            �^@                          �3@F3oU�@�           L�@                           @}ό��@�            �y@                           �?h&�}@�            @k@������������������������       ���e�D@]            @d@������������������������       � g�N�	@%             L@                          �1@Y���y@n            @h@������������������������       �ᚿ��@3            �V@������������������������       ���$��@;            �Y@                           �?Ƅp��@�           ��@                           @!�`�@�            �n@������������������������       ��Nj,@m            �d@������������������������       �WS�	@2             T@                           @78s�@            |@������������������������       �W��D�@�             s@������������������������       ��%�}��@Y             b@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        u@     �a@     �U@     �v@     �E@     }@      (@     `l@      9@     �{@      [@     �F@     �C@     �S@     @o@      P@     �u@     �s@      {@     @U@     �m@     �Y@     �H@     �p@      1@     @v@       @     �a@      .@     @u@     �O@      B@      <@      G@      f@      F@     pp@     @k@     �t@      P@     �R@      E@      ;@      W@       @      U@      @     �N@       @     @X@      3@      ,@      1@      9@      J@      2@     @V@     @U@      W@     �A@     �G@      ,@      "@      N@       @      O@              :@      @     �K@      @       @      @      &@      7@      @     �B@      D@     �K@      7@      :@      @      @      D@      �?     �@@              0@      @      7@      @      @      @       @      1@              (@      7@      D@      &@      5@      "@      @      4@      �?      =@              $@      @      @@      �?       @       @      "@      @      @      9@      1@      .@      (@      ;@      <@      2@      @@      @      6@      @     �A@      �?      E@      ,@      @      (@      ,@      =@      &@      J@     �F@     �B@      (@      :@      3@      ,@      >@      @      .@      @      ?@      �?      E@      ,@      @      &@      ,@      =@       @     �H@     �E@      B@      $@      �?      "@      @       @              @              @                              �?      �?                      @      @       @      �?       @     �d@     �N@      6@     �e@      "@      q@       @     �T@      @     `n@      F@      6@      &@      5@      _@      :@     �e@     �`@      n@      =@     �Z@      B@      2@     @`@      @     �l@       @     �P@      @     �g@      :@      4@      $@      ,@     �T@      ,@     �^@      V@     �h@      5@     @R@      5@      $@     �[@       @     `h@              J@       @     �b@      0@      ,@      "@      (@     �P@      *@     @X@      P@     @a@      1@      A@      .@       @      3@      @      B@       @      ,@       @      C@      $@      @      �?       @      0@      �?      :@      8@     �M@      @     �L@      9@      @      F@      @     �D@              0@      @      K@      2@       @      �?      @      E@      (@     �I@     �F@      F@       @      F@      ,@      @     �A@      �?      :@              (@       @      B@      1@              �?      @      6@      &@     �E@     �D@     �@@      @      *@      &@              "@      @      .@              @      �?      2@      �?       @              �?      4@      �?       @      @      &@      �?      Y@      C@     �B@     �W@      :@     @[@      @      U@      $@     @Z@     �F@      "@      &@      @@     �R@      4@      V@     @Y@     �X@      5@      E@      @      &@      E@      @     �M@      �?      9@              F@      9@      �?               @      1@      @      ;@     �E@     �C@      $@      =@      �?      @      7@              B@              *@              6@      *@                      @       @       @      "@      :@      5@      @      :@      �?      @      .@              8@              "@              .@      &@                      @      @       @      @      2@      0@      @      @              �?       @              (@              @              @       @                      �?      �?              @       @      @              *@      @      @      3@      @      7@      �?      (@              6@      (@      �?              �?      "@      @      2@      1@      2@      @      "@      @      �?      &@      �?      $@      �?      @              .@      $@      �?                      @      �?      @       @      @      @      @              @       @      @      *@               @              @       @                      �?      @      @      &@      .@      .@      �?      M@      ?@      :@      J@      5@      I@      @     �M@      $@     �N@      4@       @      &@      8@     �L@      ,@     �N@      M@      N@      &@      ;@      @      $@      4@      "@      *@       @      7@       @      <@      @      @       @      @      <@      @      $@      6@      8@      �?      7@      @      "@      0@       @       @       @      4@       @      @      @      @       @      @      *@      @      @      0@      .@      �?      @      �?      �?      @      �?      @              @              5@       @      �?                      .@              @      @      "@              ?@      :@      0@      @@      (@     �B@      �?      B@       @     �@@      ,@       @      "@      4@      =@      &@     �I@      B@      B@      $@      1@      3@      .@      =@      $@      =@      �?      5@      @      .@      *@               @      2@      *@      $@      A@      :@      4@       @      ,@      @      �?      @       @       @              .@       @      2@      �?       @      @       @      0@      �?      1@      $@      0@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ���6hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @,��9�@�	           ��@       	                    �?g�lo�D@�           ��@                            �?^7�N�@j           X�@                           �?�P@�            `s@������������������������       ��³���
@g            @b@������������������������       �@UO��@j            �d@                            �?_&c��@�           ��@������������������������       �G�ݟ�@           �y@������������������������       ����7�[@�            �k@
                          �5@�����@�           ��@                           �?���'U@\           8�@������������������������       �h-ߤ�@�            �w@������������������������       �I�]�@^           H�@                           �?�G �@7           �@������������������������       ��%��Q@�            @u@������������������������       �� al@b           x�@                           �?���:�r@�           Б@                          �:@�����@�           �@                          �7@��X�@P           ��@������������������������       �	"�t�%@�            �w@������������������������       �d��7� @a            `d@                           @ݧ��gU@]            @d@������������������������       �=k�̺@3             T@������������������������       �je���@*            �T@                           �?/Z���@           0{@                          �8@q_�oT@�            @i@������������������������       �A�`P;@k            �c@������������������������       �j��;;	@            �E@                          �1@��2`N(@�             m@������������������������       �0ˮFC@             E@������������������������       �-#�v�I@o            �g@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       @s@      b@      V@     �v@      F@     �}@      @      l@     �D@     `|@     �X@     �M@     �J@     �M@     �k@     @Q@     �u@     `s@     �}@     �R@      i@     @X@      G@      q@      :@     �u@      @     �b@      7@     pu@      L@      C@     �B@      C@     �e@      J@     @p@     �h@     @v@      J@     �K@      6@      (@      X@       @     �a@             �N@      @     �_@      .@      @      @      &@      Q@       @      U@      L@     �a@      1@      0@       @      @      H@      @      D@              <@       @     �D@      @              �?       @      8@      @      0@      8@     �D@      @      &@       @       @      2@      @      8@              .@              <@      �?              �?              @      �?      @      @      6@      @      @              @      >@      �?      0@              *@       @      *@      @                       @      2@       @      *@      3@      3@      �?     �C@      4@      @      H@      @     �Y@             �@@      @     �U@      "@      @      @      "@      F@      @      Q@      @@     @Y@      *@     �@@      .@      �?      @@      @     �K@              :@      @      J@      @      @      @      @      >@      @      F@      6@     �P@      @      @      @      @      0@             �G@              @              A@      @       @              @      ,@       @      8@      $@      A@      @     @b@     �R@      A@     @f@      2@      j@      @     �V@      2@      k@     �D@     �@@      @@      ;@      Z@      F@      f@     �a@     �j@     �A@      K@      @@      (@     �W@      �?     �a@              B@       @      ]@      $@      5@      ,@      @     �E@      4@     �X@     @U@     @^@      7@      5@      .@      @      H@      �?     �Q@              3@              ?@      @      @      @              *@      @     �D@      E@     �H@       @     �@@      1@      "@     �G@             �Q@              1@       @     @U@      @      ,@       @      @      >@      0@      M@     �E@      R@      .@      W@     �E@      6@     �T@      1@      Q@      @      K@      $@      Y@      ?@      (@      2@      7@     �N@      8@     @S@      L@     @W@      (@      D@      (@      "@      =@      &@      C@       @      .@      @      F@      ,@      �?       @      @      ;@      @     �@@      *@      6@      @      J@      ?@      *@      K@      @      >@      �?     �C@      @      L@      1@      &@      $@      3@      A@      2@      F@     �E@     �Q@      @     �Z@     �G@      E@      V@      2@     @_@      �?     �R@      2@     �[@      E@      5@      0@      5@      I@      1@     �V@     @\@      ]@      6@     �Q@      ;@      @@     �G@      0@     �O@      �?     �G@      1@     �J@     �@@      1@      (@      3@      :@      @      J@      T@     �R@      *@     �K@      *@      8@      @@      (@     �N@      �?     �D@      1@      G@      <@      .@      @      (@      4@      @      G@      I@     �G@      (@     �D@      (@      ,@      >@      $@      C@      �?      <@      @     �B@      9@      &@      @      @      .@       @      =@     �@@      C@      @      ,@      �?      $@       @       @      7@              *@      (@      "@      @      @      @       @      @      @      1@      1@      "@       @      .@      ,@       @      .@      @       @              @              @      @       @      @      @      @      �?      @      >@      ;@      �?       @      @       @      "@      �?                       @                      �?      �?      @      @      @      �?      @      0@      &@              @      $@              @      @       @              @              @      @      �?      @      �?       @              �?      ,@      0@      �?     �B@      4@      $@     �D@       @      O@              ;@      �?      M@      "@      @      @       @      8@      &@     �C@     �@@      E@      "@      1@      @      @      3@              ?@              $@      �?      =@      �?      @                      &@      @      1@      3@      <@      @      (@       @      @      1@              ?@              "@      �?      4@      �?      �?                      @      �?      &@      3@      4@       @      @      �?               @                              �?              "@              @                      @       @      @               @       @      4@      1@      @      6@       @      ?@              1@              =@       @              @       @      *@       @      6@      ,@      ,@      @      @      �?      �?      �?               @              "@              ,@                              �?                       @      �?                      0@      0@      @      5@       @      =@               @              .@       @              @      �?      *@       @      ,@      *@      ,@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhM�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@��4��r@�	           ��@       	                    @O�\�@�           8�@                           @��:&F@f           @�@                            @��"���@�           ��@������������������������       ��F;>�@           P{@������������������������       ��ٿ
W@�            �k@                           �?ωJ��	@�            ps@������������������������       �sk$0�@l            �e@������������������������       �vϲmv	@Y            `a@
                           @xE>"�@%           `|@                          �2@����@�            v@������������������������       ���#�>�@�            �o@������������������������       �p���
@=             Y@                           @�nm��	@<            @Y@������������������������       �j�g*  @             6@������������������������       �`Ѐ㎎	@0            �S@                            @$���;-@=           v�@                           @�[���@{           @�@                            �?��|B@�           �@������������������������       ���=n�U@           @y@������������������������       ����#��@�           (�@                           @�=���o@�           ��@������������������������       ��SB�P@e           h�@������������������������       ���{iޡ@o            @e@                          �?@Z��hn@�           X�@                          �;@J�@�           ��@������������������������       �`�|��	@y           ��@������������������������       �"_��
@)             L@                           �?_߄[S�@             �J@������������������������       ������
@             >@������������������������       �+<�F]	@             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �r@     @a@     �W@     �v@      :@     �~@       @      i@      =@     p|@     �Y@     �P@      A@     �I@      n@     �N@      y@     @r@     P}@     @W@     �V@      :@      8@     `b@      @     �j@      �?     �R@      �?     �g@      ?@      7@      @      $@     @U@      *@      a@     �Z@     �j@      7@     �M@      *@      (@      V@      @     `b@      �?      J@      �?     �b@      (@      ,@      @      @     @P@      @      V@     �Q@      c@      1@      I@      $@      &@     �H@      @      Z@      �?      <@             @U@      (@      *@      @      @      K@      @      P@      K@     @V@      *@      7@       @      @      B@      @      Q@              4@              P@      @      *@      @      @      C@             �C@      @@      O@      &@      ;@       @      @      *@      @      B@      �?       @              5@      @                      �?      0@      @      9@      6@      ;@       @      "@      @      �?     �C@             �E@              8@      �?     @P@              �?      @       @      &@      �?      8@      1@     �O@      @      �?                      9@              =@              4@      �?      :@                               @       @      �?      &@      @      E@      �?       @      @      �?      ,@              ,@              @             �C@              �?      @              @              *@      (@      5@      @      @@      *@      (@     �M@             �P@              6@              C@      3@      "@              @      4@       @     �H@     �A@      O@      @      :@      @      (@      K@             �B@              4@              8@      0@       @              @      &@       @     �C@      ;@      L@      @      9@      @       @      F@              7@              0@              6@      "@      @              @      @      @      1@      1@     �D@       @      �?      �?      @      $@              ,@              @               @      @      �?                      @      �?      6@      $@      .@      @      @      @              @              >@               @              ,@      @      �?                      "@              $@       @      @                                                      *@               @              �?      �?                               @               @              �?              @      @              @              1@                              *@       @      �?                      @               @       @      @             �i@      \@     �Q@     �k@      3@     @q@      @     �_@      <@     �p@     �Q@     �E@      ;@     �D@     �c@      H@     pp@     @g@     �o@     �Q@     `c@      S@      E@     �c@       @     �k@      @      R@      7@     �j@      F@      >@      0@      5@     �Z@      A@     �h@     �`@     `i@     �G@     �X@     �H@      8@     �U@      @      c@      @      K@      @     �`@      <@      1@      *@      &@      G@      ,@      \@      R@     @]@      C@     �E@      3@       @     �B@       @     �M@      @      8@       @      D@       @      @       @      @      5@      @     �@@      7@     �H@      (@      L@      >@      0@      I@      �?     @W@       @      >@       @     �W@      4@      *@      @      @      9@      &@     �S@     �H@      Q@      :@      L@      ;@      2@      R@      @     �Q@              2@      3@     @S@      0@      *@      @      $@     �N@      4@      U@     �O@     �U@      "@      C@      *@      0@      Q@      @     �I@              *@      3@      L@      ,@      $@      �?      $@     �D@      &@     �P@     �I@     �P@      "@      2@      ,@       @      @      �?      3@              @              5@       @      @       @              4@      "@      2@      (@      4@              I@      B@      <@     �N@      &@      K@      �?     �K@      @     �K@      ;@      *@      &@      4@     �H@      ,@     �P@     �I@      J@      7@      H@      ?@      6@      K@      $@      K@      �?      J@      @      I@      7@      *@      $@      .@     �H@      ,@      N@     �G@     �I@      5@      D@      :@      6@     �H@      "@      K@      �?      F@      @      I@      7@      *@      $@      *@     �C@      (@     �L@     �F@      F@      2@       @      @              @      �?                       @                                               @      $@       @      @       @      @      @       @      @      @      @      �?                      @              @      @              �?      @                      @      @      �?       @              @      @       @                              @              @      @              �?      @                      @      �?      �?               @       @      @      @      �?                                       @                               @                      �?      @               @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJFn�MhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@��q��@�	           ��@       	                     �?c��Y@�           ��@                           @�D���1@�           (�@                           �?r�
~@�            �u@������������������������       ���0��K@V            �`@������������������������       ��/2�,h@�            �j@                           @�%���
@�            �r@������������������������       ��7�x��
@}            @h@������������������������       �(ͭ�W	@A            �Z@
                           �?����%@V           X�@                           �?=��1�8@�           �@������������������������       ����rX�@�            �k@������������������������       ��E�z�
@2           0~@                           @ �n�Zy@�           P�@������������������������       �6O��ؘ@�           ��@������������������������       ��
�Z �@�            �w@                           �?w��a�@�           ��@                          �;@�P�.@e           �@                           �?��#��@           �x@������������������������       ��u��U@\             a@������������������������       �(���ډ@�             p@                           �?(����Z@b            @b@������������������������       ��y�U,L@9            �U@������������������������       �䣙�@)             N@                            @!��@e           ��@                            �?6��d�|@�           0�@������������������������       ��[�+��@�            �o@������������������������       ���X�B�@�            px@                           �?D�! �8@�            �t@������������������������       �����@A            �Y@������������������������       ��c�M�@�            �l@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     @b@     @S@     �w@      C@     @}@      @     �j@     �A@     |@     �Z@     �L@      C@      P@     �o@     �L@     �v@     �r@     �}@     @R@      d@     �L@      B@     `m@      4@     �v@             �`@      3@     �s@     �M@      @@      0@      1@     �b@      :@     �m@     `e@     `s@     �D@      B@      .@      .@      Y@      �?     @U@              ;@      *@     �T@       @      $@      @      @     �@@      "@     �L@     �@@     �W@      ,@      6@      @      @      E@      �?      E@              1@      *@     �C@      @      @      @      @      1@      @      ;@      8@     �I@      *@      *@      @              (@              4@              @              2@      �?       @      @              @              ,@      @      7@      @      "@      �?      @      >@      �?      6@              &@      *@      5@      @      @      �?      @      *@      @      *@      3@      <@      @      ,@      &@      $@      M@             �E@              $@             �E@      @      @       @              0@      @      >@      "@     �E@      �?      &@      @       @     �A@              =@              "@              >@      @      @       @              .@      @      3@      @      :@              @       @       @      7@              ,@              �?              *@              �?                      �?              &@      @      1@      �?     @_@      E@      5@     �`@      3@     @q@             @Z@      @     @m@     �I@      6@      "@      &@     @]@      1@     `f@     @a@      k@      ;@      G@      2@      "@     �N@      @     @_@              D@       @     �U@      &@      @       @       @     �B@             @R@      L@     @Z@      .@      1@      @       @      6@       @      :@              .@       @      8@      @      @       @      @      ,@              @@      .@      6@      @      =@      &@      �?     �C@       @     �X@              9@             �O@      @      @              @      7@             �D@     �D@     �T@      (@     �S@      8@      (@     �R@      .@     �b@             @P@      @     `b@      D@      .@      @      @      T@      1@     �Z@     �T@     �[@      (@      I@      *@      @     �K@      ,@     �Q@              E@      �?     �W@      :@      $@      @       @     �K@      *@     �P@      G@      U@      $@      =@      &@       @      3@      �?      T@              7@      @     �J@      ,@      @       @      �?      9@      @      D@      B@      ;@       @     �c@     @V@     �D@     �a@      2@     �Z@      @     �T@      0@     �`@      H@      9@      6@     �G@     @Z@      ?@     �_@     @_@     �d@      @@     �O@      2@      5@      J@      @     �H@      @      >@      &@     �L@      5@      �?      @      @     �@@      "@      F@      F@     �I@      .@     �J@      .@      *@     �E@      @      E@              7@      @      E@      @      �?      �?       @      9@      @     �@@      B@      D@      @      &@       @      &@      @      @      @              *@      @      .@                              �?      &@      �?      2@      0@      5@      �?      E@      *@       @     �B@      �?      C@              $@       @      ;@      @      �?      �?      �?      ,@      @      .@      4@      3@      @      $@      @       @      "@       @      @      @      @      @      .@      .@              @      @       @      @      &@       @      &@      "@      @       @       @       @      �?      �?      �?      @      @      "@      "@              @      @      @      @      @       @      @              @      �?              �?      �?      @      @              �?      @      @              �?      �?       @      �?      @      @      @      "@     �W@     �Q@      4@     �V@      (@      M@      @      J@      @      S@      ;@      8@      0@     �D@      R@      6@     �T@     @T@     �\@      1@      P@      I@      @     �I@      @     �G@              @@             �N@      4@      ,@      @      7@     �G@      1@     �M@      G@     �V@       @      :@      ;@       @      1@      @      .@              7@              &@      (@              @      &@      7@      @      8@      (@     �B@       @      C@      7@      @      A@      �?      @@              "@              I@       @      ,@      @      (@      8@      &@     �A@      A@      K@      @      >@      5@      .@     �C@      @      &@      @      4@      @      .@      @      $@      $@      2@      9@      @      7@     �A@      7@      "@       @       @              (@      �?      @              "@      @      @       @       @              &@      "@      �?      @      2@      @      @      <@      *@      .@      ;@      @      @      @      &@      �?      $@      @       @      $@      @      0@      @      2@      1@      3@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�X]hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �4@ ���o@�	           ��@       	                    �?��ֈ��@z           ��@                          �2@{�QA�@'           0�@                           @���c��@Y           P�@������������������������       ��ׇ�$�@I           ��@������������������������       �����g�@             :@                           �?/
�S,@�            �s@������������������������       ���OSQ	@^            �a@������������������������       ��'B�y@p            �e@
                           @O�Z&b@S           8�@                          �3@�-�|~@5            @������������������������       �m����@�            �v@������������������������       �&bt���@Q            �`@                           @��9"Q@           p}@������������������������       �?য��@�             w@������������������������       �J՝�6'@9            @Y@                            @��gN�[@N           8�@                           @��S���@�           ��@                          �:@�r:�[�@Q           x�@������������������������       �BX?b�@c            �@������������������������       �q³0%r@�            �w@                          �9@yv.1�U@\             a@������������������������       ��4T ��@6            �S@������������������������       ��-�Bvy
@&            �L@                          �?@#�p�@�           ��@                           @d��j��@|            �@������������������������       �2��f�@-           �|@������������������������       ��&b�!@O            @]@������������������������       � �u�s�@%             I@�t�bh�h5h8K ��h:��R�(KKKK��h��B        �r@     @[@     �V@     @x@      D@     ~@       @     @o@      ;@     �|@     @W@      M@      ;@      O@     �p@     @Q@     �u@     �s@     �{@      V@     @]@      ?@      @@      h@      3@      r@             �\@       @     �k@     �@@      5@      �?      (@     �^@      2@      d@     `b@      p@     �E@     �O@      3@      "@     �T@      @     @c@              O@             �Z@      ,@       @      �?      @     �G@      @     �K@      Q@      b@      5@      9@      *@      @      L@      @     �V@              H@             �Q@      @      @              @     �@@       @     �B@     �J@      V@      ,@      2@      *@      @      K@      @      V@              F@             �Q@      @      @              @     �@@      �?      B@      G@     �U@      ,@      @                       @               @              @                      �?                                      �?      �?      @      �?              C@      @      @      ;@              P@              ,@              B@      @      @      �?              ,@       @      2@      .@     �L@      @      1@      �?      @      "@              C@              @              5@       @      @                      $@              @       @      4@              5@      @      �?      2@              :@              "@              .@      @       @      �?              @       @      *@      @     �B@      @      K@      (@      7@     �[@      ,@     �`@             �J@       @     �\@      3@      *@              @      S@      ,@     @Z@     �S@     �[@      6@      ;@      @      1@     �N@      ,@     �K@              ;@      @     �I@      .@      (@              @     �G@       @      E@     �G@     �F@      &@      2@      @      *@     �H@      @     �G@              8@      @     �B@      *@       @              @      ?@      @      :@      B@      A@       @      "@      �?      @      (@       @       @              @       @      ,@       @      @               @      0@       @      0@      &@      &@      "@      ;@      @      @     �H@             �S@              :@      @     �O@      @      �?                      =@      @     �O@      @@     �P@      &@      6@      @      @     �E@             �L@              9@       @      I@      @      �?                      :@      @     �G@      6@     �F@      $@      @      �?              @              6@              �?      �?      *@                                      @      �?      0@      $@      5@      �?      g@     �S@      M@     `h@      5@      h@       @     �`@      3@     �m@      N@     �B@      :@      I@     �a@     �I@     `g@      e@     �g@     �F@      `@      J@     �@@     @b@      &@     �b@      �?     �Q@       @     �e@     �B@      6@      4@     �A@     �X@     �B@     @`@     @\@     �a@     �B@     �\@     �C@     �@@      b@      @      a@      �?     �N@       @     `d@      @@      6@      2@      A@     �U@      =@     �\@     �X@     ``@     �B@     �T@      =@      8@     @Z@      @     �]@      �?     �C@      @     �^@      3@      &@      @      7@      P@      &@     @T@      P@     �W@      8@      @@      $@      "@     �C@              2@              6@      �?      D@      *@      &@      ,@      &@      7@      2@      A@      A@      B@      *@      ,@      *@               @      @      &@              $@              (@      @               @      �?      &@       @      .@      .@      (@               @       @               @      @      @              @              @      @              �?              "@      @      &@       @      �?              @      @                               @              @              @                      �?      �?       @      @      @      @      &@             �K@      :@      9@     �H@      $@     �F@      �?      P@      &@     �N@      7@      .@      @      .@     �F@      ,@     �L@     �K@     �F@       @      J@      2@      6@      G@      @      F@      �?     �O@      &@      K@      3@      .@      @      ,@      F@      ,@     �J@     �G@     �F@       @     �C@      .@      6@     �C@      @      @@      �?     �M@      &@     �A@      ,@      *@       @      *@      @@      *@      D@     �C@      A@      @      *@      @              @      @      (@              @              3@      @       @      �?      �?      (@      �?      *@       @      &@       @      @       @      @      @      @      �?              �?              @      @              @      �?      �?              @       @                �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�Ȑ��@�	           ��@       	                     @^�`Ɏ@            ��@                           �?��9z�@a           L�@                          �7@�h���@�           ��@������������������������       �\�޽	@�            0w@������������������������       ���*�@�            �m@                          �5@j�n�@�           Б@������������������������       ����D@�           ��@������������������������       ����Z#�@           `y@
                           �?����{�@�           `�@                           @ML��@           �y@������������������������       �q� C�@�            0t@������������������������       �:6�d�@:            �V@                          �;@8M�7��@�            �p@������������������������       ���	M�@�            �o@������������������������       �D/d{&@
             2@                          �3@�|��@�           (�@                            �?�����@           �{@                           @��0��g@O            @\@������������������������       ���˷d
@-             P@������������������������       �v6�`h@"            �H@                           �?���w�@�            �t@������������������������       �h�e`�
@_            `a@������������������������       �����_@p            �g@                           �?���^k@�           <�@                           �?@��i@J            �@������������������������       ��|�7�s@c             d@������������������������       � ;�~��@�             x@                           @�&QG%�@C           �~@������������������������       �[� |�x@�            �w@������������������������       ��G�V��@N            @]@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       `u@      a@     �V@     �t@     �C@     �}@      &@      k@      >@     `z@      ^@     �N@     �D@      O@     @o@      M@     �v@     �s@     �|@     @W@     �i@      P@     �O@      h@      =@     �t@      $@     �b@      4@     �q@     �S@      7@      7@      C@      b@      @@     @k@     �d@     @r@     �N@     �c@      I@     �B@      b@      1@      p@      @     @X@      &@      m@     �G@      2@      .@      3@     �X@      4@      d@     �X@     �k@     �B@     �I@      >@      1@      M@      *@      L@      @     �C@      $@      O@      9@       @       @      &@      B@      ,@     �I@     �A@      N@      0@     �B@       @      *@     �G@      $@     �E@      �?      0@       @      A@      @      @      �?      $@      1@      $@      ?@      4@     �E@      $@      ,@      6@      @      &@      @      *@      @      7@       @      <@      2@      @      @      �?      3@      @      4@      .@      1@      @     �Z@      4@      4@     �U@      @     @i@              M@      �?     @e@      6@      $@      @       @     �O@      @     @[@      P@     @d@      5@     �L@      &@      @     �J@             �`@              D@             �Y@      $@      @      @      @      A@      @     @S@     �F@      `@      (@     �H@      "@      ,@      A@      @     �P@              2@      �?     �P@      (@      @              @      =@      �?      @@      3@     �@@      "@      I@      ,@      :@     �G@      (@     �R@      @      K@      "@     �K@      @@      @       @      3@      G@      (@      M@     @P@     �Q@      8@      ?@       @      7@      <@       @     �@@      @      ?@      @      =@      7@      @       @      1@      9@      $@     �E@      D@      A@      "@      8@      @      1@      8@      @      8@       @      ?@      @      6@      0@      �?      @      ,@      0@      $@      A@     �B@      7@      @      @       @      @      @      @      "@      �?                      @      @       @      @      @      "@              "@      @      &@      @      3@      @      @      3@      @      E@              7@       @      :@      "@       @               @      5@       @      .@      9@      B@      .@      3@      @      @      3@      �?      E@              7@       @      9@      "@       @               @      0@              .@      9@      A@      $@                                      @                                      �?                                      @       @                       @      @     �`@      R@      <@     �a@      $@      b@      �?     @P@      $@     �`@     �D@      C@      2@      8@     @Z@      :@     �a@     �b@     �d@      @@      A@      ,@      @     �N@             �K@              3@             �E@      &@      @              @     �A@      @      D@     �I@      I@      @      @      @       @      4@              .@              @               @       @                      �?       @              (@      $@      1@      @      @              �?      &@              @              @              �?       @                      �?       @              @      $@      &@      @      @      @      �?      "@               @                              @                                                      @              @      �?      ;@      @      @     �D@              D@              *@             �A@      "@      @               @     �@@      @      <@     �D@     �@@      @      $@       @              8@              7@               @              (@       @      �?                       @       @       @      0@      5@       @      1@      @      @      1@              1@              @              7@      @      @               @      9@      @      4@      9@      (@      �?     @Y@      M@      5@     �T@      $@     @V@      �?      G@      $@      W@      >@      @@      2@      5@     �Q@      3@     �Y@     @X@     �\@      9@      K@      D@      (@     �@@       @      ;@             �A@       @      G@      $@      (@      *@      *@     �D@       @      K@     �K@     �O@      (@      9@      @      &@      @       @      @              &@       @      "@      @              @      @      (@      @      *@      .@      6@      �?      =@      A@      �?      :@      @      5@              8@      @     �B@      @      (@      "@       @      =@      @     �D@      D@     �D@      &@     �G@      2@      "@     �H@       @      O@      �?      &@       @      G@      4@      4@      @       @      =@      &@      H@      E@      J@      *@      B@      *@      @      G@       @     �D@      �?       @       @      B@      .@      .@      �?       @      0@      @      E@      :@     �E@      *@      &@      @       @      @              5@              @              $@      @      @      @              *@      @      @      0@      "@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ}3jhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��j��@�	           ��@       	                   �5@�`yO.�@'           ��@                          �2@]Ug�4@q           @�@                            @&fi�)�@a           �@������������������������       �th�ɾ
@           �z@������������������������       ��a��Ɔ@]            �a@                          �3@.����@           �z@������������������������       �WH]�e,	@V            �a@������������������������       ��@�F�@�            �q@
                          �;@�6k)2@�           0�@                           �?60we�@U            �@������������������������       �0��>@            �i@������������������������       �s9{�DV@�            0u@                           @��k��+@a            �d@������������������������       �y5�H �@H            �^@������������������������       ���ӹ/�@            �E@                          �7@��,��@z           6�@                           @�>���@�           �@                            @����@           X�@������������������������       �wj��@]           ��@������������������������       ����6@�            �p@                           @N �:�@�           ��@������������������������       ��x�g@f            �b@������������������������       �;�����@           P|@                           @N����@�           ��@                           �?NQF��@�           ��@������������������������       �����@M            �\@������������������������       �#�-�@G           P�@                           @Z�c`�k@Z             c@������������������������       �Ni�-h�@?            @Z@������������������������       � ���.	@            �G@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       ps@     `a@     �U@     @v@     �E@     �@      @     �m@      6@     @}@     @X@      I@      F@     @Q@      k@     �P@     �v@     �r@      |@     �S@     �`@      M@     �@@     ``@      6@     pq@      @     �]@       @     �l@     �D@      2@      ,@      1@     �V@      :@     �`@     @Z@     @j@     �B@      O@      @@      (@     �U@      @      g@             �P@             �`@      2@      (@       @      @     �F@      "@     @W@     �P@     �b@      0@      9@      ,@      "@      M@      @      Z@              I@              V@       @      @      @      �?      >@      @     �K@      A@     �R@      @      1@      $@      @      D@       @     @S@             �E@             �S@      @      @      @      �?      2@      �?      B@      :@      N@       @       @      @      @      2@       @      ;@              @              "@      @              �?              (@      @      3@       @      ,@      @     �B@      2@      @      <@              T@              0@              F@      $@      @      @       @      .@      @      C@     �@@     @S@      &@      (@       @      �?       @              C@              @              2@               @                      @       @      (@      @      :@      �?      9@      $@       @      4@              E@              *@              :@      $@      @      @       @      &@      @      :@      ;@     �I@      $@     �Q@      :@      5@     �F@      2@     �W@      @     �J@       @     �X@      7@      @      @      ,@     �F@      1@      E@      C@     �M@      5@      M@      2@      &@     �C@      ,@     @U@      @      E@      @     �T@      ,@      @              @     �B@      @      <@      @@     �E@      ,@      3@      @      @      @      $@      2@      @      2@      @      <@      @       @              @      &@      @      (@      2@      :@      @     �C@      (@      @      @@      @     �P@              8@      @     �K@      &@      @                      :@       @      0@      ,@      1@      @      *@       @      $@      @      @      $@              &@       @      0@      "@              @      "@       @      &@      ,@      @      0@      @      @      @      $@       @       @      $@              @       @      *@      "@              @      @       @      @      (@      @      (@      @       @      �?              @       @                      @              @                      @       @              @       @      �?      @      @     @f@     @T@     �J@      l@      5@     �m@      @     @]@      ,@     �m@      L@      @@      >@      J@     �_@     �D@     @l@     `h@     �m@      E@      ]@     �H@      <@     �d@       @     �g@              P@      *@     �d@      @@      5@      @      5@     �R@      7@     `b@     �^@     �b@      6@      M@      =@      4@     @]@       @      V@              D@       @     �V@      9@      .@      @      5@     �E@      .@     �Q@      Q@     @S@      0@      F@      0@      (@      X@       @      K@              6@      @     @P@      .@      &@      �?      ,@     �@@       @     �C@      F@     �H@      "@      ,@      *@       @      5@      @      A@              2@       @      9@      $@      @       @      @      $@      @      ?@      8@      <@      @      M@      4@       @     �G@             �Y@              8@      @      S@      @      @      �?              @@       @     @S@     �K@     �Q@      @      "@      @       @      *@              ;@              �?              7@      @       @                      @       @      7@      &@      .@       @     �H@      *@      @      A@              S@              7@      @     �J@      @      @      �?              ;@              K@      F@      L@      @      O@      @@      9@     �N@      *@     �F@      @     �J@      �?     �Q@      8@      &@      :@      ?@     �I@      2@     �S@      R@     �V@      4@      E@      ;@      6@      K@      *@      ;@      @     �I@      �?      M@      5@      $@      8@      7@      G@      1@      M@     �L@     @P@      1@      @      @      "@       @       @      @      �?      "@              &@      @      �?       @      �?      (@               @       @      8@      @     �A@      6@      *@      G@      &@      6@       @      E@      �?     �G@      1@      "@      6@      6@      A@      1@      I@     �K@     �D@      ,@      4@      @      @      @              2@               @              *@      @      �?       @       @      @      �?      5@      .@      9@      @      (@      @      @       @              0@                              @      @      �?       @      @      @      �?      *@      @      5@       @       @                      @               @               @              @                              �?       @               @       @      @      �?�t�bub��     hhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�?�QhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?h�P�@�	           ��@       	                   �:@�UC���@�           <�@                            @�Ou��@           |�@                          �3@_�Wi$@@           P�@������������������������       ���\�
@           �y@������������������������       ��΃�#�@4           �~@                           @0�u���@�            Pu@������������������������       ���g�@�            0r@������������������������       ��gd�Q�	@             I@
                           �?�R���n@n             f@                           @�q��o*@b             c@������������������������       ��ʑ�d$@Q             _@������������������������       ��*q���@             <@������������������������       ���M5�@             8@                           @��ǆ�@           t�@                           @��n+��@�           �@                          �3@�OKdD@�           |�@������������������������       �ѥ�x~e@;           0�@������������������������       �:V�t�@�           d�@                           @�rI�4@�            �q@������������������������       ��*�#T�@�            `m@������������������������       �����-	@            �H@                           @.4��w�@q           ��@                           @1�`B�
@�            �p@������������������������       �Ԅ�/�@.            �R@������������������������       �w���
@t            �g@                           @�pː@�            `s@������������������������       �vN�T��@f            �c@������������������������       ���H�"v@i             c@�t�bh�h5h8K ��h:��R�(KKKK��h��B        @t@     �d@      Q@     �u@     �B@     �@      @     `k@      C@     0~@      [@     @Q@     �G@     �N@     �n@     �Q@      v@     `s@     �x@     @P@     �\@      C@      8@      ^@      @      o@       @     �V@       @      f@     �A@      =@      "@      3@     @W@      $@     @]@     �\@     �a@      ;@     �[@      ;@      7@     @Y@      �?     �m@      �?     �T@       @      d@      <@      0@      @      3@     @T@      @     @[@     @U@     �_@      8@     @S@      3@      ,@     �T@             `f@      �?      H@      �?      _@      (@      &@      @      (@     �N@       @     �S@     �K@      [@      1@      6@      @      @      H@              V@              2@      �?     �M@               @       @      @      @@      �?      C@      >@      J@      @     �K@      .@      &@      A@             �V@      �?      >@             @P@      (@      @       @      "@      =@      �?     �D@      9@      L@      (@     �@@       @      "@      3@      �?      M@              A@      @      B@      0@      @              @      4@       @      >@      >@      3@      @     �@@      @      "@      &@      �?     �H@              <@      @      =@      0@      @              @      .@       @      ;@      ;@      2@      @               @               @              "@              @              @                              @      @              @      @      �?      @      @      &@      �?      3@      @      (@      �?      "@              1@      @      *@      @              (@      @       @      >@      ,@      @      @      @      �?      0@      �?      (@      �?      "@              1@      @      "@      @              (@      @       @      9@      *@      @      @      @      �?      *@      �?       @      �?       @              "@      @      "@      @              (@      @      @      8@       @      @                              @              @              �?               @       @                                              @      �?      @               @      @              @       @                                               @      @                                              @      �?              j@     �_@      F@      l@     �@@      p@      @      `@      >@      s@     @R@      D@      C@      E@      c@     �N@     `m@     `h@     �o@      C@      c@     �X@      D@     �f@      >@     �f@       @      [@      ;@     �k@     �L@     �@@      =@     �C@      [@     �N@      g@      b@     `f@     �@@     �^@     �Q@      C@     �d@      4@     @c@       @     @X@      ;@     @i@      I@      ;@      2@     �@@     �U@     �D@     �c@      _@     `d@      ?@      6@      *@      *@     �P@      @      J@      �?      @@      �?      N@      0@      @       @      @      5@      1@     �Q@     �A@      S@      @     @Y@     �L@      9@     @Y@      1@     �Y@      �?     @P@      :@     �a@      A@      4@      0@      =@     @P@      8@      V@     @V@     �U@      8@      >@      =@       @      .@      $@      <@              &@              5@      @      @      &@      @      6@      4@      ;@      5@      0@       @      ;@      7@       @      (@       @      <@               @              2@      @      @      $@      @      3@      1@      ,@      5@      *@       @      @      @              @       @                      @              @                      �?              @      @      *@              @              L@      <@      @      E@      @      S@      �?      4@      @     �T@      0@      @      "@      @     �F@              I@      I@     �R@      @      ?@      �?              9@             �F@              *@      �?      B@       @      @       @              <@              4@      3@      B@       @      @                      �?              1@              @      �?      @                                      @              @      @      9@              9@      �?              8@              <@              "@              ?@       @      @       @              5@              ,@      0@      &@       @      9@      ;@      @      1@      @      ?@      �?      @       @     �G@      ,@      @      @      @      1@              >@      ?@      C@      @      $@      3@      �?      "@              1@              @              8@      @              @              &@              $@      (@      8@      �?      .@       @      @       @      @      ,@      �?               @      7@       @      @      �?      @      @              4@      3@      ,@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJl�`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?^�t��@�	           ��@       	                   �@@��e<N�@           ��@                           �?�r��@�           �@                          �6@ w�eb�@I           �@������������������������       ���i�@�            �s@������������������������       ��Th�9i@}            �h@                          �:@m�Z��@�           �@������������������������       �:���@#           @�@������������������������       �f�;݆�@�            `k@
                            @^�TOv@             F@������������������������       ���sA
@             9@������������������������       ��<�"R@             3@                           �? :�^�|@�           ��@                          �5@�s+�w�@*           ��@                           �?�p���
@j           �@������������������������       ��* ��
@M           `�@������������������������       ��/P�_@            �K@                           @:�}}4@�            �r@������������������������       �b��U�e@\            �b@������������������������       �xȣ��1@d             c@                          �6@�`!A�-@q           ��@                           @o����@L           ��@������������������������       ���o��@�             i@������������������������       ��G��f@�           ��@                          �>@�r��$@%           �|@������������������������       ������@           z@������������������������       ����-UC@            �C@�t�bh�h5h8K ��h:��R�(KKKK��h��B�       �r@      ]@     �V@     �v@     �F@     P~@       @      k@      :@     �{@      \@     �P@     �C@      S@     p@      K@     @x@     pr@     @|@     @T@     @\@     �K@      L@      d@     �A@     @b@      @      ]@      1@     �b@     �K@     �C@      4@     �F@      Z@      >@      d@     @`@      f@      @@      \@      F@     �J@     �c@     �A@     @b@      @     �[@      1@     �b@      J@     �B@      0@      F@     �Y@      =@     �c@      `@      f@      @@     �C@      $@      8@      K@      �?     �N@      @      8@      @     �F@      *@      @      @      *@     �@@      (@     �G@      C@      Q@      ,@      ?@      @      "@     �B@             �A@      �?      &@       @      9@      &@      �?      �?      $@      (@      &@      ;@      =@     �F@      &@       @      @      .@      1@      �?      :@       @      *@       @      4@       @      @      @      @      5@      �?      4@      "@      7@      @     @R@      A@      =@     �Y@      A@     @U@      @     �U@      *@      Z@     �C@      @@      &@      ?@     @Q@      1@     �[@     �V@      [@      2@      O@      7@      6@      S@      >@      T@      @     �Q@      &@     @X@      =@      9@       @      ;@     �J@      "@     �V@     �P@     @R@      0@      &@      &@      @      ;@      @      @              1@       @      @      $@      @      @      @      0@       @      4@      7@     �A@       @      �?      &@      @      @                              @              �?      @       @      @      �?       @      �?      @       @                              @      �?      @                              @              �?               @      �?               @      �?      @       @                      �?      @       @                                       @                      @              @      �?                                                     @g@     �N@      A@     @i@      $@     0u@      �?     @Y@      "@     Pr@     �L@      <@      3@      ?@      c@      8@     `l@     �d@     @q@     �H@     �Q@      "@      "@      S@       @      d@             �E@             �\@      5@      @      @      @     �O@      @      V@     �Q@     @\@      9@      F@      @             �J@              ]@              8@             �R@      *@       @       @      @      ?@              K@      H@      W@      0@      F@      @              I@             �X@              8@             �P@      *@       @              @      >@             �H@     �G@     �R@      0@                              @              1@                               @                       @              �?              @      �?      2@              :@      @      "@      7@       @     �F@              3@              D@       @      @      �?              @@      @      A@      6@      5@      "@      1@       @      @      (@       @      9@              "@              0@      @      @      �?              4@       @       @      "@      @      "@      "@       @      @      &@              4@              $@              8@      @      �?                      (@       @      :@      *@      .@              ]@      J@      9@     �_@       @     @f@      �?      M@      "@     `f@      B@      6@      0@      :@     �V@      4@     `a@     �W@     `d@      8@     �L@      9@      7@     �T@      @     �a@              E@       @     @a@      .@      2@       @      �?     �M@      .@     @[@      N@     �]@      &@      (@      @      "@      3@             �@@              @              :@      "@      @      @      �?      2@      @      8@      0@      &@             �F@      4@      ,@      P@      @     �Z@              B@       @      \@      @      *@      @             �D@      (@     @U@      F@     �Z@      &@     �M@      ;@       @     �E@      @      C@      �?      0@      @     �D@      5@      @       @      9@      ?@      @      >@     �A@     �F@      *@     �L@      :@             �E@      @      A@              0@      @     �A@      5@      @       @      3@      ?@      @      9@      A@     �A@      (@       @      �?       @                      @      �?                      @                              @                      @      �?      $@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�~�7hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?<��*p�@�	           ��@       	                    �?~)�v @           ��@                            @o nЙ@^            �@                           @� �)!@�            �s@������������������������       ���)��@f             c@������������������������       ��{!k�@i            @d@                          �7@⍶+�@�            �l@������������������������       ��:%�rD@c            `d@������������������������       �����4@,            �P@
                            @P�a��@�           $�@                          �3@��H5@�           ��@������������������������       �L�f�f�@^            `a@������������������������       ���\?@-           �~@                          �:@�Q$�!@#           P}@������������������������       �����@�            0v@������������������������       �N�g�,@@            �\@                          �4@t��5E�@�           ��@                           �? ��Yt@�           |�@                          �2@ZnPˇ@q           `�@������������������������       ���{�=e@�            x@������������������������       ����@y            `i@                           @��>��@w           ��@������������������������       ��XB|VH@           �{@������������������������       ���8�L�@^            `c@                            �?�9�h0�@�           �@                           @#�b�@�            �q@������������������������       ���<'I@;             X@������������������������       ���
���@r            �g@                           @���ѡ@            �@������������������������       ��xkH�@D           P@������������������������       ��4r�ni@�            �r@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �a@     �Y@      v@      I@      }@      @     �l@      @@      {@     �Z@     �M@     �E@      S@      n@     �N@     �t@     t@     �{@     �U@     �`@     �P@     �P@     @b@      D@      b@      @     �]@      ,@     @c@      L@      A@      ;@     �G@     �V@      >@     �_@     `c@      c@      B@     �E@      .@     �A@     �C@      *@      N@      @      E@      @      F@      7@      @      $@      &@     �B@      @     �@@      H@      O@      "@      2@      *@      3@      2@      @      A@       @      8@      �?      A@      @      @      @      @      8@      @      6@      9@     �E@      @      @       @      @      @       @      4@       @      &@              9@      @      @      @       @      @       @      @      1@      1@      @      &@      @      *@      ,@      @      ,@              *@      �?      "@              �?       @       @      1@       @      1@       @      :@      @      9@       @      0@      5@       @      :@      �?      2@      @      $@      0@              @      @      *@      @      &@      7@      3@       @      4@      �?      (@       @      @      :@              ,@              @      (@                      @      &@      �?       @      0@      .@       @      @      �?      @      *@      �?              �?      @      @      @      @              @       @       @       @      @      @      @             @V@      J@      ?@     �Z@      ;@      U@      �?      S@      "@     �[@     �@@      =@      1@      B@      K@      7@     �W@     �Z@     �V@      ;@      M@      >@      *@     �R@      $@     �F@      �?     �H@      @     @Q@       @      3@      @      (@      <@      &@      G@     �K@     �Q@      0@      ,@      @      @      4@       @      @              @      �?      $@      @       @              �?      $@      �?              3@      <@      �?      F@      :@      @      K@       @      C@      �?      G@      @     �M@      @      &@      @      &@      2@      $@      G@      B@     �E@      .@      ?@      6@      2@     �@@      1@     �C@              ;@       @     �D@      9@      $@      &@      8@      :@      (@      H@      J@      4@      &@      7@      "@      (@      1@      1@     �C@              6@       @      A@      4@      @      $@      4@      2@      @      D@     �C@      *@      "@       @      *@      @      0@                              @              @      @      @      �?      @       @       @       @      *@      @       @     @i@     �R@      B@     �i@      $@      t@             �[@      2@     `q@      I@      9@      0@      =@     �b@      ?@      j@     �d@      r@      I@     �P@      =@      1@     �Y@       @      h@             �R@      �?     �f@      6@      (@      @      @     �M@      &@     �\@     @U@     �f@      4@      :@      .@      @      L@      �?     �V@              B@              W@      @      @      @              =@      �?      G@     �H@     �\@      &@      ,@      "@      @     �A@      �?     �L@              <@              P@      �?      @      @              <@      �?     �C@      8@      O@       @      (@      @              5@             �@@               @              <@      @      �?      @              �?              @      9@      J@      @      D@      ,@      (@     �G@      �?     �Y@             �C@      �?      V@      2@      @              @      >@      $@      Q@      B@     @Q@      "@     �A@       @      @      C@              R@              B@             �O@      1@      @              �?      7@      @      E@      ;@     �J@      @      @      @      @      "@      �?      ?@              @      �?      9@      �?                      @      @      @      :@      "@      0@       @      a@      G@      3@     �Y@       @      `@              B@      1@     �X@      <@      *@      $@      8@     �V@      4@     �W@     @T@     �Z@      >@      J@      .@      "@      2@      @      A@              @              2@      &@              @      @      ;@      @      5@      7@      ;@       @      3@      @               @      @      "@              @              $@      �?              @       @      .@       @      "@      @      @      �?     �@@      $@      "@      0@              9@                               @      $@               @      @      (@      @      (@      2@      4@      @      U@      ?@      $@     @U@      @     �W@             �@@      1@      T@      1@      *@      @      2@     �O@      .@     @R@      M@      T@      6@      D@      2@      @      J@      @     @Q@              =@      1@     �I@      &@      @      @      $@     �B@      *@      I@      >@      E@      *@      F@      *@      @     �@@       @      :@              @              =@      @      @       @       @      :@       @      7@      <@      C@      "@�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�FhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�0ը�@�	           ��@       	                   �;@�z�㥯@           ��@                           @�a�[f@f           L�@                          �2@m��88>@           ؉@������������������������       �P���c{@�            @j@������������������������       �]|׽h@|           H�@                          �3@{X�@c           ��@������������������������       �eț;�{@X            �_@������������������������       ��_	�>@           �y@
                           �?�k�N@�            �q@                            @�I���_@/            @T@������������������������       ��^G�<
@'            �P@������������������������       ���i���@             ,@                            �?���mQ@y            @i@������������������������       ��;ʜ�@?            �Y@������������������������       ��"��n@:             Y@                           @����K@�           ��@                            �?�&E�r&@_           ��@                           �?G�A�u�@�           �@������������������������       �������@L           �@������������������������       ��u�l�@<           @�@                           @;���@�           �@������������������������       �(��S�~@�           �@������������������������       ��s &��@             ?@                           @@�0�J3@P           0@                           @�����@�            �r@������������������������       �:���@�            @g@������������������������       ��R�9@D             \@                            �?M�S��$@�             i@������������������������       ����H@S            �]@������������������������       �-Y0sÒ@5            �T@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       pu@      a@      T@     �w@      C@     �}@      $@     `k@      8@     {@     �W@     �P@      C@      N@     Pp@     �K@      v@     �p@     @~@      V@     �a@     @Q@     �J@     @e@      7@     @a@      "@      ]@      1@     �`@     �I@      B@      5@      D@     @^@      7@      a@     �[@     @h@     �D@     @^@     �E@      F@      b@      6@      a@       @      W@      .@      ]@     �@@      ;@      ,@      ?@     �W@      .@     �]@     �W@     �c@     �B@     �R@      0@     �@@     @R@      (@     �W@       @     �L@      "@      T@      8@      1@      @      6@     �K@      @     �R@      K@      W@      7@      2@      @      @      .@      @      0@      @      .@      �?      3@      �?               @              <@              3@      0@     �C@      �?      L@      "@      ;@      M@       @     �S@      @      E@       @     �N@      7@      1@       @      6@      ;@      @     �K@      C@     �J@      6@     �G@      ;@      &@     �Q@      $@      E@             �A@      @      B@      "@      $@      $@      "@      D@      "@     �F@      D@     @P@      ,@      $@      @      @      7@      �?      (@              @              @      @      @                      @       @      @      2@      3@      @     �B@      8@       @      H@      "@      >@              <@      @      >@      @      @      $@      "@     �B@      @     �C@      6@      G@      @      4@      :@      "@      :@      �?       @      �?      8@       @      3@      2@      "@      @      "@      :@       @      2@      1@     �B@      @      @      &@              @              �?              @      �?      ,@       @      @       @      @      @              @       @      2@               @      @              @              �?              @              *@      �?      @       @      �?      @              @       @      1@              @      @                                                      �?      �?      �?                       @                                      �?              .@      .@      "@      5@      �?      �?      �?      5@      �?      @      0@      @      @      @      5@       @      *@      .@      3@      @      @      @      @      "@              �?      �?      1@      �?       @      *@      @       @      @       @      @      @      @       @      @      "@      $@      @      (@      �?                      @              @      @       @      @       @      *@      �?      "@      (@      &@             @i@      Q@      ;@     @j@      .@     Pu@      �?     �Y@      @     �r@      F@      >@      1@      4@     �a@      @@      k@     �c@      r@     �G@     �b@      F@      5@     `d@      *@     0q@      �?     �S@      @      o@      D@      ;@      *@      .@     �X@      4@     �b@     �]@     �n@      E@      Z@      =@      $@     �V@      @      b@              B@      @      d@      ;@      *@      @      @      K@      &@     �U@     @P@     �d@      *@      J@      1@      @     �D@      @     @Q@              3@       @     @X@      1@      @      @      �?      8@      @     �I@      >@     @Q@      @      J@      (@      @     �H@       @      S@              1@      �?     �O@      $@      $@      @      @      >@       @     �A@     �A@      X@      $@     �G@      .@      &@     @R@      @     @`@      �?     �E@       @      V@      *@      ,@      @      "@     �F@      "@      P@     �J@     �S@      =@      F@      .@      &@      P@      @      `@      �?     �E@       @      V@      *@      "@      @      @     �C@      "@      P@     �J@     �R@      =@      @                      "@               @                                              @               @      @                              @             �I@      8@      @     �G@       @     �P@              8@       @      I@      @      @      @      @     �D@      (@     �P@      D@      G@      @      ;@      0@      @     �@@       @     �A@              4@      �?      <@      @       @      @      @      5@      &@     �D@      2@      8@      @      .@       @       @      ?@      �?      3@              *@      �?      5@      �?               @      @      "@      @      9@      $@      1@      @      (@       @      @       @      �?      0@              @              @      @       @      �?              (@      @      0@       @      @              8@       @              ,@              ?@              @      �?      6@              �?      �?       @      4@      �?      :@      6@      6@       @      1@       @              @              (@              @      �?      &@              �?      �?              $@      �?      7@      ,@       @       @      @                       @              3@                              &@                               @      $@              @       @      ,@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�dihG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @P
w;9�@�	           ��@       	                   �3@�EC�@�           ƫ@                            @�����@,           $�@                            �?N� b��@Q           x�@������������������������       �ot��@�           ��@������������������������       �+	���
@|            �g@                           �?��z|`@�            �u@������������������������       �Q�
��@l            @e@������������������������       �y'��j�@o             f@
                          �<@7AI��o@�           ��@                           @��$˝@�           ��@������������������������       ����2^@�           ��@������������������������       ��2L'c+@           �x@                           @1�^K"Z@�            �r@������������������������       �Qr�<GY@�            �o@������������������������       �:G���@             G@                          �4@l5Fr��@�            `v@                            �?Ν<�Ѹ@T            ``@������������������������       �v0��<�	@             D@                          �2@n�	��,@;            �V@������������������������       �=>؀Sd
@            �G@������������������������       �6�����@             F@                          �9@$N�ݔ�@�            `l@                            �?��ˈ�@K            �`@������������������������       �4qR�yi@            �E@������������������������       �&�3<J@7            @V@                           @X�l<�@=            �W@������������������������       ���S,��@+             Q@������������������������       ����Lj�@             ;@�t�bh�h5h8K ��h:��R�(KKKK��h��B        @t@     `c@     �T@     u@     �G@     �|@      &@     �j@      7@     `{@     �[@      S@     �D@      P@      n@      Q@      x@     pt@     �{@      R@     �r@     @^@     �R@     Pt@     �D@     0z@      &@      h@      7@     `y@     �W@     �P@      C@     �N@     �j@     �K@     �u@      r@     �y@     �Q@     �Z@      =@      :@     �`@      @     `f@      �?     �R@      @     �d@      9@      ;@      @       @     �S@      "@     �\@     @X@     �f@      5@     �Q@      7@      0@     �W@       @     @a@             �J@      @     �`@      "@      8@      @      @     �J@      @      W@     @P@     @a@      0@     �M@      0@      .@     @U@       @      X@              C@      @     @\@      "@      *@      @      @     �E@      @      S@      M@     �Y@      ,@      &@      @      �?      "@              E@              .@              3@              &@      �?      @      $@              0@      @      B@       @      B@      @      $@     �D@       @     �D@      �?      5@              @@      0@      @      �?      �?      :@      @      6@      @@     �F@      @      2@      @      @      9@              ;@              @              1@       @              �?               @      �?      $@      &@      9@      @      2@      @      @      0@       @      ,@      �?      ,@              .@       @      @              �?      2@      @      (@      5@      4@              h@      W@     �H@     �g@     �B@      n@      $@     �]@      4@     @n@     �Q@      D@     �@@     �J@     �`@      G@      m@     �g@     �l@     �H@     `e@     �R@      A@     @f@      :@     @k@       @     �[@      2@     `j@     �H@      A@      6@     �D@     �\@      A@      k@      e@     `h@     �E@     ``@     �M@      ?@     `b@      9@      e@       @     �Y@      2@      e@     �B@      @@      2@     �@@     @R@      A@     `e@      a@     @a@     �D@      D@      .@      @      ?@      �?      I@              @             �E@      (@       @      @       @     �D@             �F@     �@@     �L@       @      5@      2@      .@      (@      &@      6@       @      "@       @      ?@      5@      @      &@      (@      3@      (@      0@      6@     �@@      @      3@      2@      *@      "@      &@      2@       @       @       @      4@      5@      @      $@      &@      0@      &@      0@      3@      9@       @       @               @      @              @              �?              &@               @      �?      �?      @      �?              @       @      @      :@      A@       @      (@      @     �B@              5@              @@      .@      "@      @      @      <@      *@      C@     �C@      @@       @      &@      "@      @      @              7@               @              $@      @       @              �?      @      �?      1@      ,@      ,@       @      @      @      �?      @               @              @                       @      �?                                      @      @      @              @      @      @      �?              5@              �?              $@       @      �?              �?      @      �?      ,@      $@       @       @      �?      @              �?              $@              �?              @       @                              @      �?       @      @      @       @      @              @                      &@                              @              �?              �?      �?              (@      @       @              .@      9@      @      @      @      ,@              *@              6@      &@      @      @       @      8@      (@      5@      9@      2@              "@      3@       @      �?      @      @              "@              0@       @      @       @       @      .@      &@      ,@      $@       @               @      *@                      @                                      @      @      @                      @      @              @                      @      @       @      �?              @              "@              &@      @      �?       @       @      "@      @      ,@      @       @              @      @      �?      @       @      $@              @              @      @      @      �?              "@      �?      @      .@      0@              @      @      �?      @       @      "@              @              @       @      @      �?              "@              @      *@      @               @       @                              �?              �?              @      �?                                      �?       @       @      (@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJz�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?E�7�2�@�	           ��@       	                   �@@>�O�)@           ��@                           @� �R@�           ԗ@                            @iU��)@�           X�@������������������������       �LQ��O�@�           ��@������������������������       �|��O�@"            |@                           �?e!g��X@           �y@������������������������       �5���z@P             ]@������������������������       ��믉� @�            �r@
                           �?&\���@              K@������������������������       � ���,2@
             5@                           @7��&[$
@            �@@������������������������       ��}ZG�@	             &@������������������������       ����F�@             6@                           �?����p@�           <�@                          �3@pu���@*           ؊@                           @�Q��	@�            Pv@������������������������       ���E��	@�            �k@������������������������       ��Q��v@Y            �`@                          �9@p��\9�@=           `@������������������������       �WΜ��@�            �x@������������������������       �$���Q@G            �Z@                           @���J�@�           �@                           �?�ܱ�ap@           ��@������������������������       ����@�             w@������������������������       �y��I@@7           �~@                          �5@��M���@v           (�@������������������������       ���L�X%@�            �w@������������������������       ����>��@�            �l@�t�bh�h5h8K ��h:��R�(KKKK��h��B        �r@     �`@     �U@     pu@     �E@      �@      $@     �l@      ;@     P{@     �\@      Q@      D@     �P@      n@      S@      v@     �r@     p{@     @W@     �^@      P@      L@     �_@      @@     �b@       @     @[@      3@     �`@     �K@      E@      7@      H@      X@      D@     @`@     �\@     @e@     �E@     �^@     �L@     �H@     @^@      @@     @b@       @     �Z@      3@      `@     �K@      C@      1@     �F@     @W@     �A@     @`@     @[@     @e@     �E@      V@     �B@     �C@     �V@      1@     �]@       @     �Q@      0@     �S@      J@      >@      (@      9@     �Q@      9@     �V@     �U@     �^@     �@@      G@      8@      0@     �M@       @      U@      @      C@      "@     �M@      <@      7@      "@      "@      H@      *@     �G@      E@      T@      3@      E@      *@      7@      @@      .@     �A@      �?      @@      @      3@      8@      @      @      0@      6@      (@      F@     �F@      E@      ,@     �A@      4@      $@      >@      .@      ;@              B@      @     �I@      @       @      @      4@      7@      $@     �C@      6@      H@      $@      (@      �?      @      *@      @      @              "@       @      1@      @               @      "@      @      @      $@      @      &@      �?      7@      3@      @      1@      &@      5@              ;@      �?      A@               @      @      &@      3@      @      =@      1@     �B@      "@              @      @      @               @              @              @              @      @      @      @      @              @                              �?      @       @                               @                                      �?               @      @              @                              @       @      @               @              �?              @              @      @      @      �?                       @                              @      �?      �?                              �?              �?              �?               @      �?                                                      @      �?      @               @                               @              @      @      �?                               @                     �e@     �Q@      ?@      k@      &@     �v@       @     @^@       @     s@      N@      :@      1@      3@      b@      B@      l@      g@     �p@      I@     �R@      &@      "@      S@      @     �b@             �H@      �?     �^@      0@      @              @      B@      @     �T@      O@     @^@      9@      2@       @       @      B@       @      R@              >@      �?      O@       @      @              �?      @       @      B@      *@     �N@      @      *@       @              :@      �?      G@              $@             �B@       @      @              �?      @       @      6@       @      C@      @      @               @      $@      �?      :@              4@      �?      9@                                       @              ,@      @      7@      �?     �L@      "@      @      D@       @     �S@              3@             �N@      ,@      @              @      =@      @      G@     �H@      N@      3@      G@      "@      @      ;@              O@              0@             �H@      ,@       @              �?      8@              A@     �F@      I@      $@      &@              �?      *@       @      1@              @              (@              �?              @      @      @      (@      @      $@      "@      Y@      N@      6@     �a@      @     �j@       @      R@      @     �f@      F@      3@      1@      ,@     @[@      >@     �a@     �^@     �b@      9@      I@      B@      ,@     �U@      @      \@              H@      @     �\@      B@      *@      ,@      @     �M@      =@     �T@      O@      S@      ,@      ,@      .@      @      B@      @      K@              *@      @      K@      0@      @      @      �?      8@       @      ;@      A@     �C@      @      B@      5@      @      I@              M@             �A@             �N@      4@       @      "@      @     �A@      5@     �K@      <@     �B@      @      I@      8@       @      K@      @     @Y@       @      8@      �?     �P@       @      @      @      @      I@      �?      N@      N@      R@      &@      4@      *@      �?      <@             @S@              5@              F@      @      @       @              ?@              G@     �C@     �F@      @      >@      &@      @      :@      @      8@       @      @      �?      7@      @              �?      @      3@      �?      ,@      5@      ;@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�o}hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @Ҷ�ؚ@�	           ��@       	                     @���o5@�           ��@                          �7@��>z*h@S           ��@                           �?����bs@           ��@������������������������       ���D��@y           �@������������������������       �����@�           P�@                           �?��k��@?           �@������������������������       �� *�Jp@�             m@������������������������       �4]X�T�@�            0q@
                           �?��S��@�           ��@                           �?�*�I@�            �p@������������������������       ����?�3@L            @^@������������������������       ��gO*3t@]            �a@                          �;@��Nc @            �x@������������������������       �q;��o�@�             u@������������������������       �����23@             �O@                           @��~-��@�           ,�@                           @.7F�E@�           �@                           �?Ly�3dn@2           ��@������������������������       �~��T��@�             l@������������������������       �c4��m�@�           ��@                            �?t�-��@T             b@������������������������       �)����@             A@������������������������       �U��L��
@<            �[@                          �6@�/{��r@(           �|@                          �3@"�U�u�@�            �r@������������������������       ����"��	@w            �f@������������������������       �t��Y��@H            �]@                           @n� V�@i             d@������������������������       �M{���7
@$             K@������������������������       �:q�.b@E            �Z@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       @t@     ``@     �U@     pv@     �F@     �|@       @     `m@      =@     0}@     �^@     �Q@      7@     �N@      o@     �P@      v@     �r@     �|@     �P@     @j@     �P@     �M@     �f@      8@      s@       @      c@      &@     �t@      R@      B@      .@      >@     �d@     �@@     `k@      f@     `r@     �F@      d@     �E@      B@     �`@       @     @l@      @     �V@      @     @p@     �F@      9@      ,@      1@     @_@      1@     �d@     �]@     `n@      ?@      Z@      4@      :@     @Z@      @      g@      �?     �F@       @      h@      ;@      1@      @      @      U@      "@      _@     �U@      h@      8@      E@       @       @     �F@      @     �X@      �?      =@              V@      &@      $@      @      @     �A@              O@     �D@     @[@      "@      O@      (@      2@      N@      �?     @U@              0@       @      Z@      0@      @              @     �H@      "@      O@     �F@     �T@      .@      L@      7@      $@      =@      @      E@      @     �F@       @      Q@      2@       @      "@      $@     �D@       @      E@     �@@     �I@      @      3@      &@       @      .@       @      @      @      ?@       @      >@      *@      @       @      @      8@      @      2@      *@      *@      @     �B@      (@       @      ,@      �?     �A@              ,@              C@      @      @      �?      @      1@      @      8@      4@      C@       @      I@      8@      7@      H@      0@     �S@      @     �O@      @      Q@      ;@      &@      �?      *@     �C@      0@     �J@     �L@     �I@      ,@      :@      @       @      6@      @      A@      �?      5@       @      @@      @      @               @      4@      @      2@      9@      9@      @      .@      �?      @      @      @      1@      �?       @      �?      @      @      �?               @      $@       @      ,@      "@      &@      �?      &@      @      �?      .@       @      1@              *@      �?      :@       @       @                      $@      @      @      0@      ,@      @      8@      4@      .@      :@      &@      F@      @      E@      @      B@      4@       @      �?      &@      3@      &@     �A@      @@      :@      $@      3@      $@      (@      3@      @      F@      @     �D@      @      B@      3@      @      �?      "@      *@      @      :@      <@      5@      $@      @      $@      @      @      @                      �?                      �?      �?               @      @      @      "@      @      @             �\@      P@      <@      f@      5@     �c@             �T@      2@     `a@      I@      A@       @      ?@     @U@      A@     �`@      ^@     �d@      5@     @T@     �G@      6@     @_@      .@      V@              Q@       @     �Z@     �D@      ?@      @      8@      K@      :@      V@     �T@     �W@      1@     @S@     �C@      6@      \@      .@     �Q@              M@       @     @T@     �A@      9@      @      5@      K@      8@     �Q@     @R@     @S@      *@      7@      .@      "@      @@      �?      :@              ,@              (@      @      �?      �?      @      $@      "@      5@      ,@      <@       @      K@      8@      *@      T@      ,@     �F@              F@       @     @Q@      @@      8@      @      1@      F@      .@     �H@     �M@     �H@      &@      @       @              *@              1@              $@              :@      @      @              @               @      2@      $@      1@      @      @      @              "@                                              @                                                      @      @      @      @      �?      @              @              1@              $@              6@      @      @              @               @      .@      @      *@             �@@      1@      @      J@      @      Q@              ,@      $@      @@      "@      @       @      @      ?@       @     �G@     �B@      R@      @      1@      ,@      @      A@      @     �M@              &@      $@      0@      @       @       @              ,@      @      8@      7@     �I@       @      &@      $@       @      0@             �C@               @              $@       @                              @      @      *@      1@     �D@              @      @      @      2@      @      4@              @      $@      @      @       @       @              @              &@      @      $@       @      0@      @              2@      @      "@              @              0@      @      �?              @      1@      @      7@      ,@      5@       @      @                      "@       @       @                              �?       @      �?              @      @              @       @      "@              &@      @              "@      �?      �?              @              .@      �?                       @      *@      @      1@      (@      (@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJh�VxhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@T�&�@�	           ��@       	                   �2@4rŦ�*@           <�@                           @{���@�           ��@                            �?Mhԑ�@*           �}@������������������������       ��g�~�@�            �l@������������������������       ���9�s@�            �n@                           �?���k�@v           ��@������������������������       ����0��
@�            �s@������������������������       �^Q>���@�            �q@
                           @m Z=�@�            0v@                           @�"5�@y            �h@������������������������       � ��M�N@C            �Z@������������������������       �󘀼�E@6            �V@                           @��G{��@f            �c@������������������������       �n�]U��@8            �T@������������������������       �֞�l/�@.            �R@                           �?E �d@(           t�@                            @2�7�T�@           ��@                          �;@t��X@x           `�@������������������������       �S�Y؀@?           �@������������������������       �S&��@9            �S@                          �:@�1w-�@�            @p@������������������������       �I�i=:@|            �h@������������������������       �v*�@%             P@                           �?)��]��@           ��@                           @hbRf@�            �@������������������������       ���ޛ��@K             `@������������������������       �f��?�@�            �@                           @�DZ�·@           0�@������������������������       �L���@�            `w@������������������������       ��:���f@            }@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �`@     �W@     �v@      F@     P~@      "@     �l@      :@     py@      X@     @Q@      @@      Q@     �o@      S@     @v@     �s@      |@     @S@     �V@      B@      ;@      c@      @     �k@      �?      X@      @     @f@     �B@      1@      @      "@     @S@      9@     �^@      Z@      h@      :@     @Q@      6@      5@      \@      @     �d@      �?     @R@       @     �b@      6@      ,@      @      "@      F@      6@     @V@     �T@     �b@      .@      ;@      "@       @     �L@      @      O@      �?      ?@       @      E@      .@      @      @      @      >@      .@     �F@      ?@      R@       @      2@              @      A@      �?      >@               @       @      2@       @      @      �?      @      (@      @      .@      .@      I@      @      "@      "@      @      7@      @      @@      �?      7@              8@      @       @       @       @      2@      (@      >@      0@      6@      @      E@      *@      *@     �K@             �Y@              E@             �Z@      @       @       @      @      ,@      @      F@     �I@      S@      @      3@      @      @      C@             �E@              8@             �L@      �?      @      �?      �?      "@              7@      <@      H@      @      7@      @      "@      1@             �M@              2@             �H@      @      @      �?      @      @      @      5@      7@      <@              5@      ,@      @      D@              L@              7@      �?      >@      .@      @                     �@@      @     �@@      6@      F@      &@      .@      @      @      2@              8@              $@              *@      (@      �?                      2@      �?      8@      *@      >@      "@      ,@      �?       @      (@              .@              @              $@      "@      �?                       @              @      @      .@              �?      @      @      @              "@              @              @      @                              $@      �?      2@      @      .@      "@      @      $@              6@              @@              *@      �?      1@      @       @                      .@       @      "@      "@      ,@       @       @                      0@              1@              @      �?      *@      �?       @                      $@              @      @       @              @      $@              @              .@               @              @       @                              @       @      @      @      @       @      n@     �X@     �P@     �j@      C@     �p@       @     �`@      7@     �l@     �M@      J@      ;@     �M@      f@     �I@     @m@      j@      p@     �I@      M@      2@      :@      M@      &@     @]@             �N@      @      V@      4@      *@      @      7@     �K@      .@     �S@     @S@     �X@      7@     �B@      &@      ,@     �E@      @     �X@             �C@              R@      (@      $@      @      @     �@@      @      P@     �F@     @R@      *@      A@       @      &@     �D@      @     �U@             �B@             @P@      "@      @              @      ;@      @      L@      D@      P@      *@      @      @      @       @       @      &@               @              @      @      @      @      �?      @       @       @      @      "@              5@      @      (@      .@      @      3@              6@      @      0@       @      @              0@      6@       @      .@      @@      9@      $@      4@      @      $@       @      @      1@              3@      @      0@      @      �?              ,@      *@      @      *@      6@      ,@       @      �?       @       @      @      @       @              @                       @       @               @      "@      @       @      $@      &@       @     �f@     @T@     �D@     @c@      ;@     �b@       @     �R@      4@     �a@     �C@     �C@      6@      B@     �^@      B@     `c@     ``@     �c@      <@     @R@     �H@      <@     @T@      2@      L@      @     �K@      "@      O@      4@      8@      $@      6@      N@      8@      O@      I@     �U@      "@      @               @      ,@      �?      0@      @       @      @      &@      @      (@                      @       @      0@      @      0@      �?     �P@     �H@      :@     �P@      1@      D@      @     �G@      @     �I@      1@      (@      $@      6@     �K@      0@      G@     �G@     �Q@       @     @[@      @@      *@     @R@      "@      W@       @      3@      &@     �S@      3@      .@      (@      ,@      O@      (@     @W@     @T@      R@      3@      H@      6@      @      >@      @      J@              @      �?     �C@       @      @      @      �?      :@      "@     �C@      @@      :@      &@     �N@      $@      @     �E@      @      D@       @      ,@      $@      D@      &@       @      @      *@      B@      @      K@     �H@      G@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�+�(hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @��ܶ^�@�	           ��@       	                   �4@Q�r�� @�           �@                           @7:a․@P           Д@                           �?YC�tG@Y           Ѐ@������������������������       ���5$0@�            u@������������������������       �ÜE�U�@�             i@                           �?x�LV_�@�           Ј@������������������������       ��Zm4`�@           pz@������������������������       �z�p�Qo@�            0w@
                           @���'@�           �@                           �?��T��@           0�@������������������������       �q{=di@�            Px@������������������������       ��
�X��@           |@                           @��68@�           ��@������������������������       �J��3=@7           �~@������������������������       ��T��S�@U             a@                           �?b�(�Q@�           d�@                          �9@W<6��E@(           �~@                           @�{���,@�            �y@������������������������       ���u�ޯ@�            �o@������������������������       ����*�
@Y            �c@                           �?��
��@3            @T@������������������������       �G���M
@             I@������������������������       �g`�f�	@             ?@                           @�i2�@�           x�@                           @{DX�@i            �@������������������������       ��%1���@           �{@������������������������       ����ʗ@J             Y@                           �?��h-�@,            �S@������������������������       ���g�@              L@������������������������       ��_X��@             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       @t@     @a@     �Q@      w@     �F@      @      @     0p@      @@     0z@      V@      O@      D@     �Q@     pp@     �O@     Pu@     �s@      |@     @P@      l@     @Y@     �@@     �q@      <@     x@      @     �d@      4@     �s@      H@      F@      <@      E@     �g@      H@      n@     �i@     �u@      G@     @V@      8@      .@     @b@      @     @k@              R@      "@     `d@      4@      :@       @      @     �V@      .@     @\@     �Y@      h@      6@     �B@       @       @     �U@             @R@              7@      @      J@      &@      &@      �?      @      F@      @     �B@     �H@     @P@      ,@      9@       @      @     �I@             �E@              .@      @     �B@      @      @              @      <@      @      ,@      :@      G@      (@      (@              @      B@              >@               @              .@      @      @      �?              0@      @      7@      7@      3@       @      J@      0@      @     �M@      @      b@             �H@       @     �[@      "@      .@      @      �?      G@       @      S@     �J@     �_@       @      ?@      &@      @      @@      @     @R@              >@              O@      @       @      @      �?      7@              ;@      <@     �R@      @      5@      @      @      ;@              R@              3@       @     �H@      @      @      �?              7@       @     �H@      9@     �J@      @     �`@     @S@      2@     `a@      9@     �d@      @     �W@      &@      c@      <@      2@      4@     �B@      Y@     �@@      `@      Z@      c@      8@     �T@      A@      &@     @Q@      &@     �\@      @      L@      @     �Y@      0@      "@      .@      7@      G@       @     @S@     �I@     �U@      0@     �A@      *@      @     �A@       @     @P@      @      ?@      �?      J@       @      @      @      @      0@      @      A@      ?@      B@       @      H@      5@       @      A@      "@      I@              9@      @      I@       @      @      "@      3@      >@       @     �E@      4@     �I@      ,@      J@     �E@      @     �Q@      ,@      J@              C@      @      I@      (@      "@      @      ,@      K@      9@     �I@     �J@     �P@       @      A@     �D@      @     �I@      @     �D@             �@@      @     �G@      &@      @      @      &@      B@      8@     �@@      @@     �M@       @      2@       @      �?      3@      @      &@              @              @      �?       @              @      2@      �?      2@      5@      @              Y@     �B@     �B@     �T@      1@     @\@      �?     @W@      (@      Z@      D@      2@      (@      <@     @R@      .@      Y@      [@     �Y@      3@     �L@      ,@      "@     �H@      @      H@      �?     �E@       @      B@      *@      @      @      @      <@      @      E@      L@      K@      @      D@       @      "@     �G@      @      H@             �B@      @      A@      "@      @              �?      4@      @      B@      J@     �F@      @      =@      @      @      <@      @      ?@              8@      @      (@      @       @              �?      $@      @      :@      A@      1@      @      &@      �?      @      3@              1@              *@              6@       @      �?                      $@              $@      2@      <@      �?      1@      @               @      �?              �?      @      �?       @      @      @      @      @       @      �?      @      @      "@      @      (@      @               @                      �?      @      �?              @              @      @      @                      @      @              @      �?                      �?                      @               @              @                      @      �?      @               @      @     �E@      7@      <@      A@      &@     @P@              I@      @      Q@      ;@      (@      "@      7@     �F@      $@      M@      J@     �H@      (@     �B@      4@      ;@     �@@       @      K@              I@      @     �O@      7@      (@      @      4@     �@@       @      H@     �G@      D@      (@      <@      .@      8@     �@@       @     �H@              D@      @      D@      6@      &@      @      3@      :@      @      D@     �@@      @@      "@      "@      @      @                      @              $@              7@      �?      �?      �?      �?      @      �?       @      ,@       @      @      @      @      �?      �?      @      &@                              @      @              @      @      (@       @      $@      @      "@              @      @              �?      @      @                              @                      @      @       @      �?      @       @      "@                              �?                      @                                      @                              @      �?      @      @                �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��'hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@��0?]�@�	           ��@       	                   �0@ak�Q�@�           ��@                           @72ӕë
@�            @m@                           �?�|�]�?
@            �h@������������������������       �l���}�
@F             [@������������������������       �):�TI@9            @V@                           �?����G�@            �B@������������������������       �W��*�@             8@������������������������       �� �P��?             *@
                           @cLޭ�@�           ��@                           �?":'��E@�           ؄@������������������������       �փ ��
@�            �p@������������������������       ����,�@           �x@                           @�;hv@B            ~@������������������������       ���XNR/@�            �r@������������������������       ��h*��@v            �f@                          �?@�!��ғ@>           ģ@                           �?wh� >a@�           ��@                          �4@����@]           Ѝ@������������������������       ��l8�?U@_            �b@������������������������       �N��?Ú@�           �@                          �7@	]؛9�@�           ��@������������������������       ��]ls�@�           ��@������������������������       ���	��@�           ��@                            @>_�SlD@R            �`@                           @�^��'@/            �Q@������������������������       ��'�
@            �G@������������������������       ��H��
@             8@                           @y���@#            �O@������������������������       ��AGM�	@             H@������������������������       �ߙ�(�b@             .@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �`@     �V@      u@      E@     �|@       @     `k@      3@     �|@     �\@     �M@      B@     @S@     @q@     @U@     @v@     @r@     0{@     �W@      W@      >@      6@     �]@      @     �j@             �R@      @      g@      A@      4@      @      $@     �Z@      4@      ]@     @V@      k@      5@      (@       @      �?      &@             �E@              3@             �@@      @      @              @      ;@      @      *@      1@      E@              (@       @              &@              A@              .@              >@      @      @               @      9@              *@      0@      ?@              @      �?              @              0@              $@              (@      @      @               @      $@              @      $@      8@              @      �?              @              2@              @              2@                                      .@              @      @      @                              �?                      "@              @              @                               @       @      @              �?      &@                                                      "@              @               @                               @              @              �?       @                              �?                                                      �?                                       @                              "@              T@      <@      5@     �Z@      @     @e@             �K@      @     �b@      ?@      1@      @      @      T@      0@     �Y@      R@     �e@      5@      ?@      &@      1@     �Q@      @      X@              8@      @     �U@      9@      (@              @     �K@      .@     �M@     �F@     @W@      ,@      0@      �?      @      3@      �?      K@              @       @      H@      @      @                      6@      �?      6@      .@      D@      @      .@      $@      $@      J@       @      E@              3@      �?     �C@      2@      @              @     �@@      ,@     �B@      >@     �J@      &@     �H@      1@      @      B@      @     �R@              ?@      �?      P@      @      @      @              9@      �?      F@      ;@     �T@      @      ?@      @      @      9@      @     �L@              (@              ?@      @      @      @              ,@      �?      =@      $@     �N@      @      2@      &@      �?      &@              1@              3@      �?     �@@               @       @              &@              .@      1@      5@      @     @l@      Z@      Q@     �k@     �A@      o@       @      b@      .@     0q@      T@     �C@      ?@     �P@      e@     @P@      n@     `i@     @k@     �R@     �j@     @T@     �L@     �j@      @@     �n@       @     �a@      .@     �p@     @S@     �B@      :@     �K@     �d@     �M@      m@     �h@     `j@     �Q@     �^@      5@      5@     �R@      $@      ]@      @     �L@      @     �X@     �A@      *@      $@      &@     �R@      0@      U@     @U@     �S@      4@      3@               @      (@       @      3@               @              ,@       @       @      @              &@      �?      @      2@      9@      @     �Y@      5@      3@      O@       @     @X@      @     �H@      @      U@     �@@      &@      @      &@      P@      .@     @S@     �P@     �J@      0@     @W@      N@      B@     @a@      6@      `@      @     �T@      &@     �d@      E@      8@      0@      F@     @V@     �E@     �b@     �[@     �`@     �I@      F@      :@      3@     �W@      $@      V@              A@       @     �V@      .@      ,@      @      1@      E@      7@      W@      G@     �K@      ?@     �H@      A@      1@     �E@      (@      D@      @     �H@      @      S@      ;@      $@      &@      ;@     �G@      4@      L@     @P@     �S@      4@      &@      7@      &@       @      @      @              @              &@      @       @      @      (@      @      @       @      @      @      @      @      .@      @       @              @              @              @      �?       @      @       @      @      @      @      �?      @      @              ,@      @      �?              @              @              @      �?                      �?      @      @      @      �?      @              @      �?              �?                              �?              �?               @      @      �?              �?      �?              @      @      @       @       @      @      @                      �?              @       @               @      $@      �?              @      @      �?              @      @      @      @      @                                      @                       @      $@      �?               @      @                               @       @                                      �?               @       @                                               @      @      �?        �t�bub��     hhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJa}chG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�r�
��@�	           ��@       	                     �?)�P�P4@�           ¥@                           @��A��{@�           �@                          �6@��|~:D@�           �@������������������������       �Kp�ɣ@�            �w@������������������������       ��~ǽ��@�            Pp@                           @g'���@           @|@������������������������       � m���@�             w@������������������������       ��%���4@5            �T@
                           @�x���@1           p�@                          �5@Y+�Bd^@�           P�@������������������������       �,}�k�@s           �@������������������������       ���ҕ�@M           ��@                           @���K@q           @�@������������������������       ��Vb<%@B            @Y@������������������������       �83J9f�@/           0~@                           �?Qi�ӭ@�           ��@                           @m����@�           ��@                          �6@dq|O�@            @y@������������������������       ��F��o�@�            �i@������������������������       ��1�&��@u            �h@                           �?�g^2A@�            �q@������������������������       �I7JK�
@)             P@������������������������       ��N��X�@�            �k@                          �7@;c~B�/@           P{@                           @�)V�M@�            �t@������������������������       �Z�O�k@�            �j@������������������������       ��>�� @G            @]@                          �;@��>zh@E            @Z@������������������������       ���A�P�@7             U@������������������������       �%pEh��@             5@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       Pt@      b@      X@     �v@      E@      ~@      @      k@      >@     p@     �V@     �Q@      D@     �R@      m@      Q@     `w@     r@     �w@     �U@     `l@     �W@      L@     q@      4@     pw@      @     �a@      3@     �w@     �K@      M@      8@      F@      d@      J@     0p@     �g@     �r@     �I@     �Q@      I@      ;@      `@      "@      a@       @     �N@      @     �b@      5@      6@      $@      4@     �P@      3@     �U@     @R@     �\@      5@      G@      >@      ,@     �Q@      "@     �L@       @      D@      @      Q@      (@      2@      @      *@     �C@      &@      K@      I@     @S@      1@      :@       @      &@     �H@       @     �C@              *@      @     �G@      @      ,@      @      @      0@      @     �A@      A@      I@      *@      4@      6@      @      6@      @      2@       @      ;@      �?      5@       @      @      @       @      7@      @      3@      0@      ;@      @      9@      4@      *@      M@             �S@              5@      �?      T@      "@      @      @      @      ;@       @      @@      7@      C@      @      5@      $@      &@      K@              R@              *@      �?      Q@      "@      @      @      @      9@      @      4@      0@      ?@       @      @      $@       @      @              @               @              (@              �?                       @      @      (@      @      @       @     �c@     �F@      =@      b@      &@     �m@      �?      T@      (@     @m@      A@      B@      ,@      8@     �W@     �@@     �e@     @]@     @g@      >@     @Y@      B@      6@     @Z@      @     ``@      �?      K@      "@     `c@      =@      ;@      (@      ,@     �M@     �@@      ]@      N@     �]@      5@     �E@      (@      @     �O@      @     �Q@              8@       @     �S@      $@      0@      @      @      5@      (@     @S@      D@     �S@      @      M@      8@      .@      E@      �?     �N@      �?      >@      @      S@      3@      &@      "@      @      C@      5@     �C@      4@     �D@      .@     �K@      "@      @     �C@      @      [@              :@      @     �S@      @      "@       @      $@     �A@             �L@     �L@     �P@      "@      @                      @              <@              �?      @      $@                                      @              $@      @      9@      �?      I@      "@      @      @@      @      T@              9@             @Q@      @      "@       @      $@      =@             �G@      J@      E@       @     �X@     �H@      D@     �V@      6@     �Z@      @      S@      &@     @^@     �A@      *@      0@      >@      R@      0@     �\@     �X@      T@     �A@      O@      :@      >@     �J@      1@     �G@      @      D@      &@      N@      7@      "@      *@      8@      E@      $@     �S@     @S@     �G@      2@     �@@      @      5@      =@      "@      =@      @      7@      @      9@      ,@      @      @      3@      6@       @     �K@     �F@      ?@      0@      7@      @       @      *@       @      6@      �?      *@              0@      @       @       @      @      (@      �?      =@      5@      4@      �?      $@      @      *@      0@      �?      @       @      $@      @      "@      &@      @      �?      (@      $@      @      :@      8@      &@      .@      =@      3@      "@      8@       @      2@              1@      @     �A@      "@      @      $@      @      4@       @      8@      @@      0@       @       @      @       @       @              "@              �?              "@       @                              @              @      @      @              5@      (@      @      6@       @      "@              0@      @      :@      @      @      $@      @      ,@       @      1@      ;@      $@       @      B@      7@      $@     �B@      @      N@              B@             �N@      (@      @      @      @      >@      @      B@      6@     �@@      1@      9@      (@      "@      ?@       @     �J@              8@             �G@      "@      �?              @      7@      @      ;@      6@      ;@      (@      5@      "@      @      0@       @      @@              3@              :@      "@                              ,@      @      4@      (@      ,@      $@      @      @       @      .@              5@              @              5@              �?              @      "@              @      $@      *@       @      &@      &@      �?      @      @      @              (@              ,@      @      @      @       @      @       @      "@              @      @      "@       @              @      �?      @              (@              "@       @      @      @       @      @      �?      @              @      @       @      @      �?               @                                      @      �?                              @      �?       @                      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��{hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @m��}@�	           ��@       	                    @E`M��@�           J�@                          �5@e �:`@e           l�@                           @�t���@�           ��@������������������������       ���'?\@k           ��@������������������������       ���1!@<
@6           �@                           �?�"�i�@�           `�@������������������������       �?6��.�@�             t@������������������������       ����3@�            �z@
                          �;@&,�E�@�           (�@                           @�;Ko(�@9           �@������������������������       �I#��>@�            �s@������������������������       ��n⪯�@x           8�@                           @ς�D��@]            �`@������������������������       ��H0Մ�@D            �V@������������������������       ��T���@             F@                           @�5M~�9@�           ��@                          @@@�����@            ��@                           �?p�$=�m@�           ��@������������������������       �\s>��@�           ��@������������������������       �S$7��C@Z             a@                           �? ���(
@            �@@������������������������       �+�%W�@
             0@������������������������       �ę�t+@	             1@                          �6@��DL�@�            Pp@                           @�}$��h@x            @g@������������������������       �� �}�
@n            @e@������������������������       �>��_�@
             0@                           @�U3�k�@1            �R@������������������������       ���.B̧@             D@������������������������       �[��Wu@            �A@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �r@     �^@      U@     �t@     �A@     `@       @      j@      6@     �|@     �[@     �O@      @@     �R@      p@      M@     �v@     pu@     �|@      U@     �i@     @U@     �G@     �n@      5@     �w@       @     `b@      *@     `w@     �Q@     �F@      9@      J@     �g@      E@      p@     `m@     �v@      H@      `@      O@      5@     �a@       @     �q@       @     @W@      @     �p@     �D@      9@      .@      7@     �^@      4@     �e@     �a@     @k@      A@     �P@      :@       @     �Y@              h@              K@      @     �c@      (@      .@      @      @     �P@      @     �X@     @W@      b@      1@     �D@      1@       @      O@             �S@              6@      @     �U@      @      $@              @      >@      @      O@      G@     �Q@      .@      :@      "@             �D@             @\@              @@              R@      @      @      @              B@      �?     �B@     �G@     �R@       @     �N@      B@      *@     �B@       @     �V@       @     �C@      @     �Z@      =@      $@      &@      3@     �L@      0@     @R@     �G@     @R@      1@      9@       @      @      3@       @      F@      �?      4@      @      M@      1@       @      @       @      :@      @      <@      .@      >@       @      B@      <@       @      2@      @      G@      �?      3@             �H@      (@       @      @      1@      ?@      *@     �F@      @@     �E@      "@     @S@      7@      :@     @Z@      *@     �X@      @      K@      @     @[@      =@      4@      $@      =@     �P@      6@     �U@     �W@      b@      ,@      P@      7@      1@     �W@      $@     �W@              G@      @     �W@      7@      3@      $@      :@     �O@      2@     @T@     �S@      ^@      $@      (@      @      @     �D@      @      B@              3@      �?      <@      *@      0@      @      $@      7@      "@      4@      9@     �@@       @      J@      3@      $@      K@      @      M@              ;@      @     �P@      $@      @      @      0@      D@      "@     �N@      K@     �U@       @      *@              "@      $@      @      @      @       @              ,@      @      �?              @      @      @      @      0@      9@      @      @              @       @       @      @               @              &@      @      �?              @      @      @      @      ,@      &@      @      @              @       @      �?      �?      @                      @      �?                              �?              �?       @      ,@              X@     �B@     �B@     �T@      ,@     �^@              O@      "@     �U@      D@      2@      @      7@     �P@      0@     �Z@      [@     �W@      B@      Q@      @@      B@     �J@      (@     �U@              H@      "@      L@      <@      ,@      @      3@      I@      .@     �U@     @V@     �M@      ?@     @P@      @@      @@     �I@       @     �U@             �G@      "@      L@      ;@      ,@      @      .@      I@      .@     �T@      U@      L@      ?@     �G@      8@      ;@      E@       @      P@             �D@       @      E@      6@      ,@      @      .@      F@      $@     �Q@     @R@      I@      7@      2@       @      @      "@              7@              @      �?      ,@      @                              @      @      &@      &@      @       @      @              @       @      @                      �?                      �?              �?      @                      @      @      @               @              �?      �?                              �?                      �?              �?                              @      �?      @              �?              @      �?      @                                                                      @                              @                      <@      @      �?      >@       @     �A@              ,@              >@      (@      @      �?      @      0@      �?      3@      3@     �A@      @      2@      �?      �?      8@       @     �A@              ,@              9@      @      @               @       @              $@      ,@      6@       @      2@      �?      �?      8@       @     �@@              (@              8@      @      �?               @      @              @      ,@      4@       @                                               @               @              �?               @                      @              @               @              $@      @              @                                              @      @      �?      �?       @       @      �?      "@      @      *@      @      @                      @                                              �?      @                              @      �?      @      �?      $@              @      @              �?                                              @       @      �?      �?       @      @              @      @      @      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��"hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?Gc`�`�@�	           ��@       	                     @ۏ�	�@�           ��@                          �5@�s�~�9@U           ��@                          �1@��kz�@           �z@������������������������       �!��In�
@>            �V@������������������������       ��O�7@�             u@                           @c����@?           �~@������������������������       �AJ'��@�            `u@������������������������       �$���@i             c@
                          �4@}0,B��@�           (�@                           �?�ew�@�            `m@������������������������       ���_9@?            �Y@������������������������       ��N|@W            �`@                           @����[@           �{@������������������������       ���x�&@�            �t@������������������������       �DtԤ.�@G             [@                           @X֭<�_@�           �@                           @(��!�@           �@                            @T�qt#@s           ��@������������������������       ����i@           �z@������������������������       ���QXj@f            `e@                            �?Εv��@�           H�@������������������������       �)��"+$@�            `x@������������������������       ����6�4@�            0r@                           @K�wX�@w           @�@                           @�U�Ӎ@�           ��@������������������������       �oYw��	@�            �q@������������������������       �kW�F@�            `w@                           @oZ�`�@�            �w@������������������������       ��j��J�@=            @X@������������������������       �	��ݎ	@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �r@     �`@     @U@     �w@     �B@      |@      (@     �n@      6@     �~@      W@     �H@      >@     �V@     �k@     �Q@     �v@     �r@     �|@     �S@     �]@     @R@     �H@     �d@      6@     �_@      &@     �\@      1@     �c@     �C@      :@      (@      N@      R@      C@     �c@     `b@     �c@     �A@     @P@     �C@      8@      Y@      "@     �P@      @      P@       @     �\@      2@      3@      @      ;@     �D@      <@     @V@     �N@      \@      4@      >@      ,@      @     �N@      �?      E@              ;@      @     �G@      @      $@      �?      @      5@      @     �F@      =@      N@      $@      &@              @      "@      �?      $@              @              $@                      �?       @      @      �?      �?       @      4@              3@      ,@       @      J@              @@              5@      @     �B@      @      $@              @      0@      @      F@      5@      D@      $@     �A@      9@      1@     �C@       @      9@      @     �B@       @      Q@      ,@      "@      @      5@      4@      7@      F@      @@      J@      $@      ;@      2@      *@      8@      @      5@      @      ?@             �H@      ,@       @      @       @      0@      ,@      @@      6@      8@      @       @      @      @      .@      @      @              @       @      3@              �?      @      *@      @      "@      (@      $@      <@      @      K@      A@      9@      P@      *@      N@      @     �I@      "@     �E@      5@      @      @     �@@      ?@      $@      Q@     �U@      F@      .@      5@       @      $@      .@      "@      :@       @      *@       @      &@      "@       @      @      @      *@      @      A@      <@      8@      @      ,@      �?      @       @              1@              @              @      @              @      �?       @       @      1@      &@      @      �?      @      �?      @      @      "@      "@       @      @       @      @      @       @              @      &@      �?      1@      1@      4@      @     �@@      @@      .@     �H@      @      A@       @      C@      @      @@      (@      @       @      =@      2@      @      A@      M@      4@      &@      <@      5@      .@      C@      �?      2@       @      <@      @      2@      $@      @      �?      5@      ,@      @      >@      H@      0@      &@      @      &@              &@      @      0@              $@      �?      ,@       @       @      �?       @      @       @      @      $@      @             �f@      N@      B@     @k@      .@     0t@      �?      `@      @     �t@     �J@      7@      2@      >@     �b@      @@     @j@     �b@     0s@      F@     �X@      F@      5@      _@      &@     `d@             �S@      �?      g@     �B@      ,@      $@      (@     �T@      =@     �^@     �R@      b@      8@     �L@      6@      "@      L@      @     �Q@             �A@             �R@      4@      @      @      @      L@      *@      J@      F@     �H@      *@      H@      &@      @     �E@      @      G@              1@              K@      ,@       @      @      @     �E@      @     �C@     �A@     �D@      @      "@      &@      @      *@      �?      9@              2@              4@      @       @      �?      �?      *@      "@      *@      "@       @      @     �D@      6@      (@      Q@      @      W@             �E@      �?     �[@      1@      $@      @      @      :@      0@     �Q@      ?@      X@      &@      4@      (@       @     �I@      �?     �J@              &@              O@      @      @      @      @      .@      @     �B@      2@     @Q@       @      5@      $@      @      1@      @     �C@              @@      �?     �H@      &@      @      �?      �?      &@      "@      A@      *@      ;@      @     �T@      0@      .@     �W@      @      d@      �?     �I@      @      b@      0@      "@       @      2@      Q@      @     �U@      S@     @d@      4@     �H@      $@      @      J@             �X@             �B@      �?     @Z@      $@      @      @      @      E@      �?     �L@      G@     �\@      (@      4@              @      ;@              L@              3@      �?     �E@      @      �?      �?               @              5@      2@     �L@      @      =@      $@      @      9@             �E@              2@              O@      @      @      @      @      A@      �?      B@      <@      M@       @      A@      @       @      E@      @     �N@      �?      ,@      @      D@      @      @      @      (@      :@       @      >@      >@     �G@       @      @              @      (@       @      0@      �?      @      �?      @      @      �?       @      @      @              @      @      1@              ;@      @      �?      >@       @     �F@              &@       @     �B@      @      @       @      @      3@       @      8@      ;@      >@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�L0�@�	           ��@       	                    �?ɸ �e@           ,�@                          �:@����=@o           ��@                            �?��yŴ:@*           �|@������������������������       ���'�"�@V            �a@������������������������       �a��'��@�            �s@                           �?(F��^�@E             Z@������������������������       �,  �}�	@             7@������������������������       �≮��?@3            @T@
                          �5@"�%�@�           l�@                           �?�'`$@           @}@������������������������       �z�/B�u@R             b@������������������������       ��2%"@�            @t@                           �?豟�s?@�           8�@������������������������       ����Wi@x             i@������������������������       ��5d�C@           �{@                           @���즨@t           |�@                           @�F�_k@]           ��@                            �?Bh�\�@v            �@������������������������       �$ڐ��@�            pv@������������������������       �m��3@�             k@                           @S�t͇@�            py@������������������������       �ntӛO}@�             p@������������������������       ������@[            �b@                          �3@!/�1��@           ��@                            @�%<h@o           p�@������������������������       ��r�>�
@3           P~@������������������������       ����"J@<            @Z@                          �<@�l�4�C@�           Ȅ@������������������������       ��:`ǵ@�           �@������������������������       �'�Iݭ
@&             N@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �b@      U@     �u@     �D@     P}@      @      k@      A@     {@     @[@     @T@      F@     @P@      l@      T@     �x@     �s@     z@     �U@     �^@      P@     �M@     �c@      ;@      a@      @      ]@      9@     �a@      G@     �I@      8@      F@     @V@     �F@     `f@     �a@     �c@     �E@      D@      &@      9@      A@       @      N@      �?     �D@       @      N@      0@      &@      @      $@      7@      (@     �K@     �J@     @Q@      0@      ?@      "@      0@      >@      @      M@              ;@      @     �K@      &@      &@       @      @      1@      @      G@     �H@      M@      ,@      &@      @       @      (@       @      1@              "@              8@              @      �?      @      @              @      ,@      1@      "@      4@      @      ,@      2@      @     �D@              2@      @      ?@      &@      @      �?       @      &@      @      E@     �A@     �D@      @      "@       @      "@      @       @       @      �?      ,@      @      @      @              @      @      @      @      "@      @      &@       @       @              �?                       @              @       @      @                      �?      �?              �?              �?      @              @       @       @      @       @              �?      &@      @      �?      @              @      @      @      @      "@      @      @       @     �T@     �J@      A@     @_@      3@      S@      @     �R@      1@     �T@      >@      D@      1@      A@     �P@     �@@      _@     �U@      V@      ;@     �E@      $@      ,@     �P@      $@      C@              <@      (@     �B@       @      1@      �?      &@      5@      *@      N@     �C@      ;@      *@      5@      @      @      ?@       @      @               @      @      ,@      �?      @              @      @      @      .@      @      @      @      6@      @      &@     �A@       @     �@@              4@       @      7@      @      (@      �?      @      .@      @     �F@     �A@      6@      $@      D@     �E@      4@     �M@      "@      C@      @     �G@      @      G@      6@      7@      0@      7@     �F@      4@      P@      H@     �N@      ,@      ,@      "@      $@      5@      �?      0@      �?      5@              0@      $@      @      @      @      &@      @      .@      "@      7@      �?      :@      A@      $@      C@       @      6@      @      :@      @      >@      (@      1@      $@      3@      A@      *@     �H@     �C@      C@      *@     @h@      U@      9@     �g@      ,@     �t@      �?      Y@      "@      r@     �O@      >@      4@      5@      a@     �A@     �j@     �e@     @p@      F@     �S@     �D@      .@      R@      $@      `@             �D@       @     �_@      >@      2@      .@      "@      Q@      7@     �[@      S@     �V@      <@     �L@      4@      @      G@      @     �R@              =@       @      M@      9@      $@      "@      @     �H@      .@     �N@     �D@     �H@      *@      >@      *@      �?      ?@      @     �E@              ,@              ?@      3@      @      @      @     �@@      "@      B@      ;@      G@      @      ;@      @      @      .@       @      ?@              .@       @      ;@      @      @      @      @      0@      @      9@      ,@      @      @      5@      5@      "@      :@      @      K@              (@             @Q@      @       @      @      @      3@       @      I@     �A@      E@      .@      @      *@      @      .@      @     �B@              @             �D@      �?      @       @      �?      3@       @      D@      7@      8@      (@      1@       @      @      &@              1@              @              <@      @       @      @       @              @      $@      (@      2@      @      ]@     �E@      $@     �]@      @     �i@      �?     �M@      @     `d@     �@@      (@      @      (@      Q@      (@      Z@     @X@      e@      0@      H@      5@      @      G@       @     @\@              C@             @U@      @       @      @      @      @@      @      D@      A@     �X@      �?      A@      .@      @      D@       @     @W@              8@             �R@       @      @      @              ;@      @      B@     �@@      V@              ,@      @       @      @              4@              ,@              $@       @       @              @      @      @      @      �?      &@      �?      Q@      6@      @     @R@       @      W@      �?      5@      @     �S@      =@      @      �?      "@      B@      @      P@     �O@     �Q@      .@     �N@      1@       @     @R@             �U@              5@      @      S@      9@      @              @     �A@      @     �O@     �I@      M@      .@      @      @      @               @      @      �?                       @      @              �?      @      �?              �?      (@      (@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ���~hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?F���_�@�	           ��@       	                    @U�xg @�           �@                            @��@�           |�@                          �?@M^>�'w@           ��@������������������������       ������E@           ��@������������������������       �P�����@             ;@                          �:@��K@~           `�@������������������������       �N"���@@4           �~@������������������������       ��đp�@J            @`@
                            �?۟{�OR@b            @c@                           �?j�ɾ��	@             D@������������������������       �TY�	�@
             *@������������������������       ���пT@             ;@                           �?�U#!�@F            �\@������������������������       ����&
i@             B@������������������������       �6�fe�@1            �S@                          �4@v���@�            �@                           @o׾���@           �@                            @�I����@g            �@������������������������       �75�e@�           `�@������������������������       �Q���%@o            �f@                          �3@;vU��6@�            �q@������������������������       ������V
@�            �j@������������������������       ��5J�	@)            �P@                          �9@�?�@�           X�@                          �6@Pm04[\@�           ��@������������������������       �Fn[�@�            �t@������������������������       �Q�u^6@�            �x@                           �?�cT@�            �s@������������������������       �
�K��@a            �a@������������������������       �s���@l             f@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@     @`@     �U@     �t@     �I@     �@      @     `k@      =@      }@     �]@      L@      D@     �R@     �m@      K@     �u@     s@     �z@     �U@     @_@      Q@     �K@     �^@      C@     `b@      @      W@      4@     �b@      L@     �B@      <@     �M@      V@      >@     �_@     @`@     @e@     �H@      [@     �L@      K@     �\@      <@      ^@      @     �U@      3@     �`@     �J@      B@      9@     �J@     @T@      9@     �[@     �^@      d@      H@      I@     �A@      3@     @U@      $@     �R@       @      D@      @      V@      ;@      3@      1@      3@      K@      ,@     �M@     @P@     �Z@      >@     �H@      <@      2@     @U@      $@      R@       @     �A@      @      V@      ;@      2@      1@      2@      K@      $@     �M@     @P@      Z@      <@      �?      @      �?                      @              @                              �?              �?              @                       @       @      M@      6@     �A@      >@      2@     �F@      �?      G@      ,@     �G@      :@      1@       @      A@      ;@      &@     �I@      M@      K@      2@     �F@      ,@      3@      <@      2@     �F@      �?      >@      $@     �C@      6@      0@      @      :@      4@       @      I@     �E@     �@@      2@      *@       @      0@       @                              0@      @       @      @      �?      @       @      @      @      �?      .@      5@              1@      &@      �?       @      $@      ;@              @      �?      *@      @      �?      @      @      @      @      1@      @      $@      �?      @      @                      @       @               @              "@                       @      @               @              �?      �?      �?       @      �?                              @              �?              �?                                                              �?      �?               @      @                      @       @              �?               @                       @      @               @                              �?      *@      @      �?       @      @      3@              @      �?      @      @      �?      �?      @      @      @      1@      @      "@              @              �?      @      @      @               @      �?      �?      @                              @       @       @      �?                      @      @              @      @      .@               @              @              �?      �?      @      @      �?      .@      @      "@             `k@      O@      @@      j@      *@     Pv@      �?     �_@      "@     �s@      O@      3@      (@      0@     �b@      8@     `k@     �e@     @p@      C@     �V@      4@      *@      `@       @     @k@             �T@       @     �g@      ,@      (@      "@      @     �S@      (@     @^@     @W@     �e@      *@     @R@      0@      $@     @\@      �?      e@             �R@      �?     �c@      *@       @       @       @      K@       @     �S@     �L@     `a@      (@      K@      ,@      $@     �U@             `a@              L@      �?     ``@      $@       @       @      �?     �E@      @     @R@      H@     �]@      @      3@       @              :@      �?      =@              2@              9@      @                      �?      &@       @      @      "@      5@      @      2@      @      @      0@      �?      I@               @      �?     �@@      �?      @      �?      �?      8@      @      E@      B@      A@      �?      .@      @      �?      (@             �E@              @              =@      �?      �?              �?      7@      @      8@      7@      ;@              @               @      @      �?      @              �?      �?      @              @      �?              �?              2@      *@      @      �?      `@      E@      3@      T@      &@     `a@      �?     �F@      @      `@      H@      @      @      *@     �Q@      (@     �X@     �T@     �U@      9@      V@      A@      *@     �O@      @      Z@              <@      @     @X@     �B@       @               @      J@      $@     �Q@      N@      C@      ,@      7@      ,@      @      7@      @     �P@              *@      @      H@      ,@       @              @      5@       @     �C@      8@      3@      @     @P@      4@      @      D@              C@              .@      @     �H@      7@                      @      ?@       @      ?@      B@      3@      "@      D@       @      @      1@       @     �A@      �?      1@      �?      @@      &@      @      @      @      2@       @      <@      6@     �H@      &@      .@      @       @      @      @      $@      �?      $@      �?      4@      @      @      �?              @       @      &@      &@      2@      $@      9@      @      @      $@      @      9@              @              (@      @       @       @      @      (@              1@      &@      ?@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��KhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?h!���@�	           ��@       	                    �?���@           ��@                          �8@�:-w�@J           @�@                          �7@~7�%�J@�             w@������������������������       �kY?.@�            �t@������������������������       ����Р@             B@                           �?�n���@_             c@������������������������       ��X�x@             E@������������������������       ��V��@D            �[@
                          @@@�^;�@�           ��@                           �?�ƣ���@�           ��@������������������������       �`;�{�@0            �R@������������������������       �2�y���@i           (�@                           �?pC��'
@!            �K@������������������������       �l�u5x@             4@������������������������       ������@            �A@                           @�)J��O@�           ��@                           @��f���@,           ��@                          �5@a�8���@e           H�@������������������������       ���F��@`           X�@������������������������       �k��X@           �y@                            @��4.�@�            ps@������������������������       �<�N@�            �o@������������������������       ���f��@(            �M@                            @C�J��8@g           ؍@                           @'����@           ��@������������������������       ���d�@�            Py@������������������������       �_�:P/@           �y@                           �?-�u.4=@_            �`@������������������������       �I�[���	@,             Q@������������������������       �]��|@@3            �P@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@      `@     �S@     �v@     �A@      }@      @     @m@      :@      {@     �]@     �O@     �C@     �O@      m@     �Q@     px@     �r@      |@     �N@     `b@      Q@      L@     �c@      7@     �b@      @     @]@      0@     �a@     �I@     �A@      8@     �D@     @V@     �E@     �b@     �`@     `e@      9@      F@      *@      6@     �D@      @     �H@             �E@      �?     �O@      2@      0@       @      @      >@      *@      E@     �B@     �P@      @     �A@       @       @      ?@      �?     �B@              @@              K@       @      @      @      @      2@       @      ;@      ;@      L@      @     �A@       @      @      ?@      �?     �B@              ;@             �G@      @      @      �?      @      2@      @      7@      7@     �G@      @                      �?                                      @              @       @               @                      �?      @      @      "@      �?      "@      @      ,@      $@       @      (@              &@      �?      "@      $@      &@      @      �?      (@      @      .@      $@      $@              @      �?      @       @              @               @              �?      @      @      @              @      �?      �?       @      @              @      @       @       @       @       @              "@      �?       @      @      @       @      �?      @      @      ,@       @      @             �Y@     �K@      A@     �\@      4@      Y@      @     �R@      .@      T@     �@@      3@      0@     �A@     �M@      >@     @[@     �X@     @Z@      4@     �Y@     �F@      @@     �[@      1@      Y@      @     �P@      .@      T@      ?@      3@      (@     �A@     �M@      :@     �Z@     �U@     �Y@      4@      @      @               @              ,@              @       @       @              @              @       @      �?      @      ,@       @       @     �X@      C@      @@     �Y@      1@     �U@      @     �O@      *@     �S@      ?@      0@      (@      =@     �L@      9@     �Y@      R@      Y@      2@      �?      $@       @      @      @                      @                       @              @                      @      @      (@      @                      @      �?      �?                              @                       @              �?                      @      �?              �?              �?      @      �?      @      @                      �?                                      @                               @      (@       @             �i@      N@      6@      j@      (@     �s@             @]@      $@     0r@      Q@      <@      .@      6@      b@      ;@      n@      e@     pq@      B@     �Z@     �B@      *@     �a@      "@     �d@             �Q@      @      e@      H@      3@      &@      *@     @R@      ;@     @a@     �W@      b@      :@     @U@      A@      &@      \@      @      Z@              F@      @     @a@      D@      *@      @      (@      O@      2@     �Z@      R@      \@      7@      =@      5@      @      Q@             �K@              7@             �U@      6@      $@      @      @      @@      (@     @S@      E@     �T@      $@      L@      *@      @      F@      @     �H@              5@      @     �I@      2@      @      @      @      >@      @      >@      >@      =@      *@      6@      @       @      <@      @     �O@              :@       @      ?@       @      @      @      �?      &@      "@      ?@      7@     �@@      @      ,@      @      �?      ;@      �?      L@              4@       @      9@       @      @      @      �?       @      @      7@      3@      <@      �?       @              �?      �?      @      @              @              @                                      @      @       @      @      @       @     @X@      7@      "@     @Q@      @     �b@             �G@      @     �^@      4@      "@      @      "@     �Q@             �Y@     @R@     �`@      $@     @V@      2@      "@     �I@      @     ``@              C@      @     @Z@      3@      @       @      @      O@             �W@      L@     @]@      @     �F@       @       @      9@       @     �S@              5@      @     �J@       @      @      �?      �?      >@              C@      ?@      M@      @      F@      0@      @      :@      �?      J@              1@      �?      J@      1@       @      �?      @      @@             �L@      9@     �M@      �?       @      @              2@              1@              "@              1@      �?       @       @      @      "@              @      1@      1@      @      @      @              ,@              &@              @              @                                      @               @      @      $@       @      �?       @              @              @              @              (@      �?       @       @      @      @              @      &@      @      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��}?hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?�
p��@�	           ��@       	                   �@@��I�@           ��@                           @�|e@�           ��@                           �?C�v���@V           h�@������������������������       �x�h@�            �t@������������������������       �O�F�@~           ��@                           �?��]��@�           �@������������������������       �yE����@z             h@������������������������       ��E<`��@            |@
                            @PK���@"            �J@                          @A@>��_@             @@������������������������       �����@             0@������������������������       �����@
             0@������������������������       ���3�@             5@                           �?؋F�	@�           ̡@                          �3@.M�,�@(           ��@                            @������	@           �z@������������������������       ��OJ��	@�             u@������������������������       �*����	@/            @V@                            @��A��0@!           �|@������������������������       ��Le@�            �w@������������������������       �?ӿ��@1            �T@                            �?�<E��u@c           ȕ@                          �5@Y�pw�@           Њ@������������������������       �/��>�@=           @�@������������������������       �O�9��@�             u@                          �6@��
�Y�@U           ��@������������������������       �y{��
@�            Pu@������������������������       �ĝ�ؖ#@x            `h@�t�bh�h5h8K ��h:��R�(KKKK��h��B        �r@     �`@     @W@     �v@     �J@     �~@      (@     �n@      =@     P{@     �W@      L@      D@     �P@     �j@      O@      y@     0s@      {@     �R@      \@     �P@     �M@     �c@      A@     @_@      $@     �`@      5@      ^@      K@      >@      7@      H@      W@      A@     �d@     �c@      c@      F@      \@     �K@     �L@     �b@      A@     @_@      $@      _@      5@     �]@     �H@      <@      3@      G@      V@      @@     `d@     �c@     �b@      F@      L@      4@     �B@     �U@      5@      V@      $@     �Q@      "@     @S@      D@      0@      *@      <@     �F@      .@     �W@     @Z@     �U@      8@      6@      @      3@      <@             �B@      @      7@      @      9@      ,@       @       @      @      2@      @      <@     �B@      D@      $@      A@      ,@      2@      M@      5@     �I@      @      H@      @      J@      :@       @      &@      8@      ;@       @     �P@      Q@      G@      ,@      L@     �A@      4@     �O@      *@     �B@             �J@      (@     �D@      "@      (@      @      2@     �E@      1@     @Q@     �J@      P@      4@      ?@      @      $@      .@      @      @              1@       @      "@      @               @       @      1@      @      9@      3@      3@      �?      9@      ?@      $@      H@       @      ?@              B@      $@      @@      @      (@      @      0@      :@      (@      F@      A@     �F@      3@              &@       @      @                               @               @      @       @      @       @      @       @      �?      �?       @                       @              @                               @              �?               @                      @       @      �?                                       @              @                              @              �?                                       @       @                                              @              @                               @                               @                       @              �?                                      @       @      �?                                              �?      @              @       @                              �?       @             @g@     @Q@      A@     @j@      3@      w@       @     �\@       @     �s@      D@      :@      1@      2@     �^@      <@     �m@     �b@     �q@      >@     �R@      3@      0@     @P@      @     @d@             �H@       @     @^@      &@       @      �?      @     �E@      @     �W@     �I@     ``@      3@     �B@       @      @     �@@      @     �Y@              5@       @      P@      @      �?               @      0@       @      F@      5@      P@      @      <@      �?      �?      <@      �?     �T@              3@       @     �F@              �?                      0@       @     �D@      (@      K@      @      "@      �?      @      @      @      4@               @              3@      @                       @                      @      "@      $@              C@      1@      (@      @@      @      N@              <@             �L@       @      @      �?       @      ;@      @     �I@      >@     �P@      0@      =@      (@      (@      ;@       @      L@              4@              H@      @      @      �?       @      .@       @      G@      >@      M@      "@      "@      @              @      �?      @               @              "@      @      @                      (@      �?      @              "@      @     �[@      I@      2@      b@      (@      j@       @     �P@      @     �h@      =@      2@      0@      ,@      T@      7@     �a@     @X@     �b@      &@     �R@      9@      *@     @S@      $@     @\@              A@      @     @_@      8@      $@      ,@      @     �J@      (@     �V@     @Q@      X@      "@      =@      ,@      @      C@             @S@              9@             �U@      "@       @      *@      @      9@       @     �O@      I@      N@      @      G@      &@      @     �C@      $@      B@              "@      @      C@      .@       @      �?       @      <@      @      ;@      3@      B@      @      B@      9@      @      Q@       @     �W@       @      @@       @     �Q@      @       @       @      "@      ;@      &@     �I@      <@     �K@       @      3@      (@       @     �B@      �?     �R@              5@              I@      @       @              @      ,@      �?     �C@      2@     �B@      �?      1@      *@      @      ?@      �?      4@       @      &@       @      5@       @               @      @      *@      $@      (@      $@      2@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJW��WhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B                             @������@�	           ��@       	                     @����|@�	           �@                            �?]��#@�           ��@                          �3@t�Wm?p@\           ��@������������������������       �9����q@           �@������������������������       ��s�,@Z           Д@                          �6@o����@�            �@������������������������       ��p�o�@�            Py@������������������������       �ؔ��>@�            `m@
                           @�t�3@�           �@                           @�:Ă@           `�@������������������������       �)�
!H4@�           (�@������������������������       ��Pm�7x@*            �Q@                          �5@��2�O�@�            �p@������������������������       ��3���W@r             f@������������������������       ����^J@6            @W@                          �6@�*�8i
@)            �O@                          �3@�u�	3�@            �A@������������������������       ���	M�1@	             0@������������������������       �I���}f@             3@                           �?��i���@             <@������������������������       �7�nt@
             ,@������������������������       �;%Ͳ�� @	             ,@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     ``@     �U@     @w@      A@     �@      *@      m@      8@      |@     �X@     �I@      @@     �R@     `m@      O@     �v@     ps@     pz@     �S@     �t@     @`@     �U@      w@      =@     �@      *@      l@      8@     �{@     �X@     �I@      >@     �R@     �l@      N@      v@      s@     �y@     �S@     �l@     �T@     �I@      q@      3@      x@      &@     �a@      *@     �t@      P@     �D@      4@      H@     �e@      D@     �o@      j@      t@     �M@     `e@     @Q@      C@     @k@      .@     pp@      $@     @\@      $@     `n@      N@      >@      3@     �B@     �`@     �A@      i@     �c@     @p@     �H@     �@@      1@      $@     �X@       @     @Y@             �F@      @      ^@      1@      (@      @      @      L@      @     @R@     �K@     @_@      ,@     @a@      J@      <@     �]@      *@     @d@      $@      Q@      @     �^@     �E@      2@      0@      ?@     @S@      =@     �_@     @Y@     �`@     �A@     �L@      ,@      *@      L@      @     �^@      �?      ;@      @      W@      @      &@      �?      &@     �D@      @     �J@      J@      O@      $@      =@      @      @      B@       @     �U@              6@              L@      @       @              $@      9@             �D@      ;@      F@      @      <@      &@      @      4@       @      B@      �?      @      @      B@      �?      @      �?      �?      0@      @      (@      9@      2@      @      Y@     �G@      B@      X@      $@     @_@       @     @U@      &@     @[@     �A@      $@      $@      :@     �L@      4@     �X@      X@      V@      3@     @T@      C@      A@      Q@      "@     �V@       @      O@      &@     @R@      =@       @      $@      7@     �G@      1@     @Q@     @S@      J@      (@     �R@      >@      ?@      O@      @     @T@       @      N@      $@     �Q@      7@       @      @      4@     �E@      (@     �P@     �R@      I@      &@      @       @      @      @      @      "@               @      �?       @      @              @      @      @      @      @      @       @      �?      3@      "@       @      <@      �?     �A@              7@              B@      @       @              @      $@      @      >@      3@      B@      @      "@      @      �?      1@              ;@              4@              ?@      @      �?               @       @      @      (@      $@      ;@      @      $@      @      �?      &@      �?       @              @              @       @      �?              �?       @              2@      "@      "@      @      �?      �?               @      @       @              @              @                       @              @       @      &@      @      *@              �?                       @      �?       @              @              @                       @                               @       @       @                                       @              �?               @                                                                      @       @      @              �?                              �?      �?              @              @                       @                              @              @                      �?                      @                      �?              @                                      @       @      @      @      @                      �?                      @                      �?              �?                                      @              @              �?                                                                                       @                                      �?       @              @      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ?�rhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �? ;�[�@�	           ��@       	                     @ ��@           �@                           �?��	C@a           P�@                           �?>��;�@           �z@������������������������       �����G@X            @b@������������������������       ��x.��)@�            �q@                           �?9;��B�@^           �@������������������������       ������@|            `g@������������������������       ��<-�ށ@�            t@
                           @�'>`@�           ��@                          �?@�|���@3           0�@������������������������       ���>	�@%           �~@������������������������       �h2|wO�@             <@                          �3@�v��:@�            @j@������������������������       �LD��v@"             F@������������������������       ����
�@b            �d@                            @�?��3=@�           ��@                          �6@8�$1�@{           ��@                            �?Q\�r��@            ��@������������������������       �~o�/a@4           ��@������������������������       �_X�9�	@�            `r@                           �?�d̵�@{           (�@������������������������       �26��-�@�            �q@������������������������       ������@�            `t@                           �?#����@	           @z@                          �7@3h:&�@�            �l@������������������������       �0G�	q@i             e@������������������������       ��b ��"
@$            �O@                           @��g@|            �g@������������������������       �}˶�0�@R            @_@������������������������       �����p+
@*             P@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       t@      `@     @V@     �u@      F@     @@      (@     �l@      C@     �{@     �Y@     �L@      G@     �O@     `o@     �J@     0x@     �q@     �{@      R@     �]@     �P@      L@     �`@      <@     �b@      &@     @_@      =@      c@      E@     �B@      8@      H@     �Z@      9@     �c@     �`@     �f@      E@     �Q@     �E@      :@      X@      @      V@      @      I@      &@      \@      *@      ,@      3@      6@     �I@      1@     �U@     �L@     @^@      @@     �B@      .@      .@     �F@              I@              .@      �?     �F@      @      @      @      $@      <@       @      C@      3@     �P@      6@      .@      @       @      @              0@              �?              1@              �?              @      (@              "@      (@     �@@      @      6@      &@      @      C@              A@              ,@      �?      <@      @      @      @      @      0@       @      =@      @     �@@      1@     �@@      <@      &@     �I@      @      C@      @     �A@      $@     �P@       @      "@      *@      (@      7@      "@      H@      C@     �K@      $@      "@      @      @      1@      �?      9@       @      2@              :@      @      @      @      �?      "@      @      9@      @      1@      �?      8@      6@      @      A@      @      *@      @      1@      $@     �D@      @      @      @      &@      ,@      @      7@      ?@      C@      "@      H@      7@      >@      B@      8@     �O@      @     �R@      2@      D@      =@      7@      @      :@     �K@       @     @R@     �R@      O@      $@      8@      (@      6@      :@      3@     �F@      @     �L@      ,@      4@      :@      ,@      @      5@     �C@      @     �L@     �J@     �H@      @      8@       @      0@      :@      1@     �F@      @     �L@      ,@      4@      7@      ,@      @      1@     �C@      @      L@      G@     �H@      @              @      @               @                                              @              �?      @                      �?      @                      8@      &@       @      $@      @      2@              2@      @      4@      @      "@              @      0@      �?      0@      6@      *@      @       @       @      @      @              "@              �?               @       @                              @              @      @      �?      @      6@      "@      @      @      @      "@              1@      @      2@      �?      "@              @      *@      �?      (@      0@      (@      @     `i@     �O@     �@@     @k@      0@     �u@      �?     �Z@      "@     r@      N@      4@      6@      .@      b@      <@     �l@     �b@     pp@      >@     �c@      H@      7@     �g@      ,@     �r@      �?     �S@       @      l@      G@      ,@      5@      "@     @_@      2@     �h@     @]@     @k@      5@      S@      7@      $@     @_@      @     `m@             �O@      @     �b@      7@      (@      0@       @      S@       @     �a@     �P@     @d@      1@      O@      6@       @     �Y@      @     �c@              G@      @     �Z@      4@      "@      .@             �K@       @     @[@      K@     �^@      ,@      ,@      �?       @      7@      �?      S@              1@             �D@      @      @      �?       @      5@              A@      *@     �C@      @      T@      9@      *@     �O@      "@     �O@      �?      0@      @      S@      7@       @      @      @     �H@      $@      L@      I@      L@      @     �E@      (@      @      B@      "@     �@@      �?      "@      @      =@       @              @      �?      9@      @      1@      6@      4@      @     �B@      *@      @      ;@              >@              @             �G@      .@       @       @      @      8@      @     �C@      <@      B@             �G@      .@      $@      >@       @     �I@              ;@      �?     @P@      ,@      @      �?      @      4@      $@      =@      @@     �F@      "@      9@      @      @      6@      �?      ?@              2@      �?     �F@      @      @                       @      @      *@      2@      4@      @      3@      @      @      2@      �?      ?@              &@      �?      ;@      �?                              @      �?      "@      0@      ,@      @      @      @              @                              @              2@       @      @                      �?      @      @       @      @      �?      6@      "@      @       @      �?      4@              "@              4@      &@              �?      @      (@      @      0@      ,@      9@      @      3@      @      @       @      �?      0@              @              @      &@              �?      @      @      @      $@      @      1@      @      @       @      �?      @              @              @              .@                               @      @              @       @       @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJj;�yhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�2����@�	           ��@       	                   �7@�����@*           ��@                           �?�Ȯ��/@c           ��@                            @l>��9!@�            v@������������������������       ����ʿ@y            @h@������������������������       ��]��;�@f            �c@                            @a9JюU@�           ��@������������������������       ���F�&�@�            x@������������������������       �]7�mL&@�             n@
                           @Oi��f@�           ��@                          �9@�7�j'T@@           @@������������������������       ����ӻ�@u            �g@������������������������       �%{�ϩ�@�            `s@                           �?�M���@�            `l@������������������������       �/��.��@!             K@������������������������       �r��,E�@f            �e@                          �6@K�f�9S@t           >�@                           @I��T�@�           ��@                          �2@fR���@x           H�@������������������������       ���tZ�
@�            �o@������������������������       �hL�W[x@�            �t@                          �5@���_� @6           ،@������������������������       �	N�2��@           �@������������������������       ��=Ը�O
@4            @V@                           @�o�@�           ؅@                           �?�,����@�           ��@������������������������       ���E
��@�            0s@������������������������       ��a��ޭ@�            @t@                          �<@�V9�.�
@,             Q@������������������������       ���u�n	@"            �I@������������������������       �X�SZ@
             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       Pu@     �]@     �V@      u@      C@     �{@      @     �n@     �B@     0|@      [@     �P@      F@     @Q@     `o@      P@     Pu@     �s@     P|@      X@     @b@     �Q@      M@     @c@      ;@     �[@      @     �a@      ?@     `c@      M@      E@      6@      G@     �[@      @@     @a@     �b@     �d@     �G@     @W@      B@      :@      \@      0@     �R@       @     @Q@      1@     �W@      @@      *@      @      1@     @Q@      0@     �S@     �U@     @Y@      7@     �B@      @      "@     �A@       @      C@      �?      ?@              ;@      &@      @       @      @      4@       @      <@      B@      F@      @      3@      @       @      5@       @      ;@      �?      0@              5@      �?      �?                      (@      @      *@      2@      >@      @      2@      @      @      ,@      @      &@              .@              @      $@       @       @      @       @      @      .@      2@      ,@       @      L@      >@      1@     @S@       @      B@      �?      C@      1@      Q@      5@      $@       @      ,@     �H@       @      I@      I@     �L@      1@     �D@      1@       @     �L@      @      ,@              2@      "@      F@      $@      @              &@      7@      @     �@@      ;@     �C@      0@      .@      *@      "@      4@      @      6@      �?      4@       @      8@      &@      @       @      @      :@      �?      1@      7@      2@      �?     �J@      A@      @@      E@      &@     �B@      @      R@      ,@      N@      :@      =@      2@      =@      E@      0@      N@      O@     �O@      8@     �B@      0@      <@      8@       @      7@      @      N@      &@     �B@      :@      6@       @      1@      ?@      "@     �C@      F@      C@      3@      "@       @      .@      @      @      (@       @      1@      @      7@      &@      @      @      "@      $@              ,@      1@      "@      2@      <@      ,@      *@      3@      @      &@      �?     �E@      @      ,@      .@      2@      @       @      5@      "@      9@      ;@      =@      �?      0@      2@      @      2@      @      ,@              (@      @      7@              @      $@      (@      &@      @      5@      2@      9@      @      @      @       @                       @               @              @                               @                      &@      @      "@              *@      &@       @      2@      @      @              $@      @      1@              @      $@      $@      &@      @      $@      ,@      0@      @     `h@      H@      @@      g@      &@     �t@      �?     �Y@      @     �r@      I@      8@      6@      7@     �a@      @@     `i@     @e@     r@     �H@     @]@      ;@      8@      _@       @      p@             @S@      @     �h@      <@      6@      .@      @     �T@      0@     `b@      ]@      k@      ;@      F@      (@      @     �M@             �U@              5@             @U@      *@      $@       @      @     �A@      *@     �P@      A@     @R@      2@      .@      �?      �?      >@             �D@               @             �F@       @      �?              @       @      @      ;@      *@     �C@      @      =@      &@      @      =@             �F@              *@              D@      @      "@       @              ;@      @     �C@      5@      A@      &@     @R@      .@      3@     @P@       @     @e@              L@      @     @\@      .@      (@      @      @     �G@      @     @T@     �T@      b@      "@      Q@      .@      $@     �L@      �?     �b@             �G@      @     �Y@      ,@      (@      @      @      F@      @     �Q@     �T@      a@      @      @              "@       @      �?      4@              "@       @      &@      �?                              @              &@              @       @     �S@      5@       @      N@      "@     @R@      �?      :@             �X@      6@       @      @      0@      M@      0@      L@      K@      R@      6@      Q@      4@       @     �M@      "@     �P@      �?      6@             �W@      .@       @      @      0@     �F@      *@      I@     �F@     @Q@      6@     �A@       @      @      9@       @     �B@      �?      $@              K@      @       @      �?      �?      3@      @      1@      ?@      >@      2@     �@@      2@      @      A@      �?      >@              (@              D@      "@              @      .@      :@      @     �@@      ,@     �C@      @      $@      �?              �?              @              @              @      @              �?              *@      @      @      "@      @              "@      �?              �?              @               @              @      @              �?              *@      @      �?      @      �?              �?                                                       @                      @                                              @      @       @        �t�bub��     hhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ-�bhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �6@o��:�@�	           ��@                           @�>|��j@�           ʢ@                           @�\�2S�@�           ��@                            �?JS1��@�           @�@������������������������       �i=*��@�           �@������������������������       ��7@�0p@M           p�@������������������������       �rW`�q�@             9@                           �?��e�I�@           �@	       
                   �3@mF ��=@           z@������������������������       �۬�ߞ%
@�            �r@������������������������       ��|9���
@V            @]@                          �5@�[R�@�           ؈@������������������������       �5��]@d@�           ��@������������������������       ��I\h��	@B             Z@                            @BX�E@�           ��@                          �>@{�J�3Y@�           ��@                           �?�TQ�@7           ��@������������������������       ��d��6�@�            �u@������������������������       �ϰ���@N           �@                           �?�Oc]�+@N            �]@������������������������       ���U+V@-            �P@������������������������       ��ӿ#ء	@!             J@                           @[�ґp@*            @                           �?�K�L9_@�            �u@������������������������       ��xk�c@�            `o@������������������������       �ID�N\@?            �X@                          �<@1o��آ@Y            �b@������������������������       ��h`L@@            �Z@������������������������       ��	�.`@             E@�t�bh�h5h8K ��h:��R�(KKKK��h��B        �t@     �`@     �T@      u@     �I@     �}@       @     `i@     �F@     �z@     �X@      J@      B@     �Q@      m@     �Q@     @y@      s@     �|@     �U@      e@     �N@     �G@     �h@      3@      x@      @     �_@      9@     @r@     �C@      ?@      .@      1@     �a@      ?@     `p@     `h@     `s@     �C@      Y@     �B@      C@     @Z@      1@     `b@      @      P@      .@     �^@      8@      3@       @      *@     @Q@      7@     �`@     @Z@     �`@      3@     �X@      B@      C@     @Z@      ,@     `b@      @     �K@      .@      ^@      8@      3@      @      *@     @Q@      7@     �_@     @Z@     �`@      3@      H@      *@      7@     �P@      @      R@              8@      .@     @Q@       @      ,@      @      @      B@      "@     �P@      M@     �W@      (@     �I@      7@      .@     �C@      &@     �R@      @      ?@             �I@      0@      @      �?      @     �@@      ,@     �M@     �G@      C@      @      �?      �?                      @                      "@               @                       @                              @                             @Q@      8@      "@      W@       @     �m@             �O@      $@     @e@      .@      (@      @      @     @R@       @      `@     �V@     @f@      4@      B@      @      @      9@      �?      Y@              <@      @     �E@      "@       @              @      <@       @     �C@      8@     �M@      @      >@              �?      3@      �?     @R@              :@      @     �B@       @       @              @      ,@       @      3@      0@     �H@      @      @      @      @      @              ;@               @              @      @                      �?      ,@              4@       @      $@      @     �@@      5@      @     �P@      �?      a@             �A@      @     �_@      @      $@      @             �F@      @     �V@     �P@     �]@      ,@      >@      4@       @      M@              [@              =@       @     �[@      @      $@      @              C@      @     @S@      O@     �\@      *@      @      �?       @      "@      �?      =@              @      @      1@      �?                              @              *@      @      @      �?      d@     �R@      B@     `a@      @@     �W@      @      S@      4@      a@     �M@      5@      5@     �J@     �V@      D@     �a@     �[@     �b@      H@      \@      G@      8@      W@      .@      Q@      @     �F@      @     �X@      A@      &@      (@      A@     �Q@      9@     �Z@     @Q@     �[@      <@     @Y@      A@      0@     �V@      .@      N@       @     �D@      @     �U@     �@@       @      (@      7@      Q@      4@      X@     �P@      W@      8@      8@      .@      &@      C@      "@      (@       @      :@              ?@      ,@      @      @      (@      <@      @      A@      4@     �B@      *@     @S@      3@      @     �J@      @      H@              .@      @      L@      3@      �?      @      &@      D@      *@      O@      G@     �K@      &@      &@      (@       @      �?               @      �?      @       @      (@      �?      @              &@      @      @      &@      @      2@      @      @      (@      @                       @              @       @      @              @              @      @      @      @       @      "@       @       @              @      �?              @      �?                      @      �?                       @                      @      �?      "@       @     �H@      <@      (@     �G@      1@      :@       @      ?@      .@      C@      9@      $@      "@      3@      3@      .@     �A@      E@     �C@      4@     �B@      1@      $@      B@      &@      2@       @      8@      *@      ,@      6@      @      @      *@      0@       @      >@      >@      2@      4@      4@      "@      @      @@       @      $@       @      .@      (@      @      1@      @      @      (@      ,@      @      2@      7@      .@      .@      1@       @      @      @      @       @              "@      �?      "@      @      �?              �?       @      �?      (@      @      @      @      (@      &@       @      &@      @       @              @       @      8@      @      @      @      @      @      @      @      (@      5@              &@      @      �?      @      @       @              @       @      5@      �?      @       @       @      �?      @      @      @      1@              �?       @      �?      @       @                      �?              @       @              �?      @       @              �?       @      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJөWhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�nY�.�@�	           ��@       	                    @������@           @�@                          �;@iAy�i�@�           �@                          �:@��u��1@�           ��@������������������������       �2+�;6@e           ��@������������������������       �	�A�n8@              I@                          �@@~"+_@i            @e@������������������������       ����z�@Z            �b@������������������������       ���l}@             6@
                           �?=�Lb�@,           P}@                           @���@_             b@������������������������       �=5���@:            @W@������������������������       ����v��
@%             J@                            �?2����@�            @t@������������������������       ����s�s@D            �Z@������������������������       �J���@�             k@                           �?�Hj�@�           �@                            @��\{\@�           ��@                            �?�]����@�           h�@������������������������       �1����@t            @e@������������������������       �8 �F0�
@           0|@                          �2@w,|%��@^             b@������������������������       ���@%             M@������������������������       �����@9            �U@                           @�;��E@�           �@                          �3@������@/           Ћ@������������������������       �ʴ�8�@�            �t@������������������������       �����U@Y           ��@                            �?��C,@�           �@������������������������       ��
�(:�@�            �w@������������������������       ��S��_@�            `p@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@     �]@     @V@     @u@      C@      ~@      $@     @i@     �@@     P|@      \@      R@      H@     �T@     �n@     �M@     �w@      s@     �z@      Q@     �`@      N@     �G@     �b@      7@     �b@       @      Y@      8@     @e@      H@      C@      <@     �I@     @Z@      3@      b@      `@     �c@      ?@     �W@      B@      ?@      \@      $@     �\@       @     �R@      5@     �Z@     �C@      6@      1@      @@     @P@      .@     �[@     @V@     �^@      :@      T@      2@      7@     �W@      "@     @[@       @      M@      1@     @Y@      <@      4@      $@      :@     �K@      .@     @X@     �R@      \@      6@      T@      2@      5@     @V@      "@     �Z@       @     �K@      0@     @Y@      <@      2@      $@      :@     �J@      (@     @X@     �O@     �W@      6@                       @      @              @              @      �?                       @                       @      @              &@      1@              .@      2@       @      1@      �?      @              1@      @      @      &@       @      @      @      $@              *@      .@      &@      @      .@      (@      @      .@      �?      @              .@      @      @      "@      �?      @       @      $@              *@      .@      &@      @              @       @       @                               @                       @      �?      @      @                                                      C@      8@      0@     �B@      *@     �A@              9@      @      P@      "@      0@      &@      3@      D@      @     �A@     �C@      B@      @      $@      $@      @      &@      �?      ,@              �?              6@      @              �?      @      0@      �?      .@      .@      &@      �?      @      @       @       @              $@                              .@      @              �?      @      ,@              ,@      @      @      �?      @      @       @      "@      �?      @              �?              @                                       @      �?      �?      "@      @              <@      ,@      (@      :@      (@      5@              8@      @      E@      @      0@      $@      *@      8@      @      4@      8@      9@      @      @      $@       @      *@      @       @              @      �?      "@               @      @      @       @      @      @      @      $@       @      6@      @      $@      *@      @      3@              3@       @     �@@      @       @      @      @      0@              1@      1@      .@       @     `j@     �M@      E@     �g@      .@     �t@       @     �Y@      "@     �q@      P@      A@      4@      @@     �a@      D@     @m@     @f@     �p@     �B@      K@      @      0@     �P@      @     `a@              F@      �?     �V@      5@      @      �?      @      K@      @     �R@     �L@     �Y@      1@      E@      @      $@     �M@      �?      ^@             �A@      �?     �S@      &@      @      �?      @      D@      @      N@     �D@      W@      (@      "@              @      2@      �?      :@              *@      �?      <@      @                      �?      *@      @      $@      .@      3@       @     �@@      @      @     �D@             �W@              6@             �I@      @      @      �?      @      ;@      �?      I@      :@     @R@      $@      (@      @      @       @       @      3@              "@              &@      $@                      @      ,@      �?      .@      0@      &@      @      "@              @      @      �?       @              @              @      @                      @      �?              @      $@      �?              @      @      @      @      �?      &@              @              @      @                              *@      �?      "@      @      $@      @     �c@      J@      :@      _@      (@      h@       @      M@       @      h@     �E@      >@      3@      9@     �U@      A@     �c@     @^@      e@      4@     �U@      9@      .@      U@      "@     �[@             �F@      @     �\@      @@      ,@      &@      1@      J@     �@@     �U@     �N@     @S@      (@      .@      �?      @      E@              G@              6@              J@      @      @      �?      �?      3@      $@      E@      8@     �A@       @     �Q@      8@      &@      E@      "@      P@              7@      @     �O@      9@      @      $@      0@     �@@      7@     �F@     �B@      E@      $@     �Q@      ;@      &@      D@      @     �T@       @      *@      @     �S@      &@      0@       @       @     �A@      �?      R@      N@     �V@       @      I@      6@      @      4@      �?     �F@              "@              F@       @      @      @      @      0@      �?     �J@      A@      I@      @      5@      @       @      4@       @      C@       @      @      @      A@      @      $@      �?       @      3@              3@      :@     �D@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�-�9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?ҿ��U�@�	           ��@       	                     @�iL���@?           ��@                           �?k����@X           �@                            �?t�ooMX@�            �s@������������������������       ���
�S@`            �b@������������������������       �����"@g            `d@                           @08��.a@�           P�@������������������������       �`P#/�
@1           �}@������������������������       �J�`�1@`             b@
                           �?���n@�            px@                           �?{"�?��@�             k@������������������������       �gC<�n@/             S@������������������������       �fs�@��@S            �a@                           @C��4M@e            �e@������������������������       ��"9��i@'            �P@������������������������       ��lb�@>            @[@                          �6@fv���@m           @�@                          �5@>:��Y�@�           \�@                           �?�;CM`�@;           ̓@������������������������       ��g�5�@)           P}@������������������������       ��p���@           ��@                           �?�/r�ӂ@�            �l@������������������������       ������@A             [@������������������������       �ԫaE<6@I             ^@                           @���O�@�           $�@                           �?�燞�@�           ؄@������������������������       ��w,S��@�             o@������������������������       ���zs��@            z@                           �?��t��@           �z@������������������������       �����@k            `c@������������������������       ��C��
@�            0q@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@      a@     �T@     @w@      D@     0|@      "@     @m@      >@     0|@     @[@     �M@      >@     @T@     �l@      L@     `u@     ps@     �}@     @U@     �Z@      =@     �A@      Z@      $@     �e@      �?     �T@      @     �c@      D@      (@      $@      4@     @U@      $@     �_@      ]@      d@     �B@     �M@      5@      7@     @T@      @     �a@             �K@      �?     @^@      2@      @      "@      "@     �M@      @      X@      T@      `@      .@      7@      "@      &@      3@      @      <@              1@             �B@      .@      @      "@      @      7@      �?     �@@      <@     �D@       @      (@      @      @      ,@      �?      0@              ,@              5@      @      �?      @       @      &@      �?       @      &@      *@      @      &@      @      @      @       @      (@              @              0@      $@      @      @      �?      (@              9@      1@      <@      @      B@      (@      (@      O@      �?     @\@              C@      �?      U@      @      @              @      B@       @     �O@      J@     �U@      @      7@      @      @     �G@      �?      W@              ?@             @P@      �?      @              @      ?@       @     �J@     �D@      N@      @      *@      @       @      .@              5@              @      �?      3@       @                      �?      @              $@      &@      ;@             �G@       @      (@      7@      @      A@      �?      ;@      @      B@      6@      @      �?      &@      :@      @      >@      B@     �@@      6@      4@      @      $@      *@      @      .@      �?      6@      @      0@      (@      @      �?      $@      ,@      @      4@      4@      2@      @       @      @      �?      @              @      �?      "@      �?      @      @              �?      @      $@              @      (@      @              (@      @      "@      $@      @      &@              *@      @      "@      @      @              @      @      @      .@       @      .@      @      ;@       @       @      $@      @      3@              @              4@      $@       @              �?      (@      @      $@      0@      .@      2@      $@      �?       @      @              @              �?              $@       @       @                      @      �?               @      @      $@      1@      �?              @      @      *@              @              $@       @                      �?       @       @      $@       @      &@       @     `l@     �Z@      H@     �p@      >@     @q@       @      c@      9@     `r@     @Q@     �G@      4@     �N@      b@      G@      k@     `h@     ps@      H@     �^@     �J@      =@     @c@      (@     `h@      �?     �R@      "@     �i@     �A@      >@       @      .@      R@      7@      b@      [@     �f@      9@     �Y@      H@      9@      `@      @     �c@             @Q@      @     �c@      <@      <@       @      *@      L@      0@      _@      Z@     �d@      8@      E@      ,@      &@     �F@      @     �I@             �@@      @     �A@      1@      &@      @       @      =@      @      B@      G@      L@      *@     �N@      A@      ,@     �T@             �Z@              B@              _@      &@      1@      @      @      ;@      $@      V@      M@      [@      &@      3@      @      @      :@      @      C@      �?      @       @     �F@      @       @               @      0@      @      4@      @      1@      �?      &@               @      "@      @      5@      �?      �?      �?      5@      @      �?               @      @      @      @       @       @               @      @       @      1@              1@              @      �?      8@      �?      �?                      "@      @      .@       @      "@      �?     @Z@      K@      3@     �\@      2@     @T@      @     @S@      0@     �V@      A@      1@      (@      G@      R@      7@      R@     �U@     @`@      7@     @P@      =@      $@     �R@      $@      N@      @      K@      (@      D@      8@      ,@       @      <@     �B@      $@     �C@      M@      Q@      4@      6@      @      �?      6@      @      >@      @      6@      (@      4@       @      @      @      @      &@      �?      1@      7@      @@      �?     �E@      7@      "@      J@      @      >@      @      @@              4@      0@      &@      @      6@      :@      "@      6@     �A@      B@      3@      D@      9@      "@      D@       @      5@              7@      @      I@      $@      @      @      2@     �A@      *@     �@@      =@      O@      @      1@      "@      @      0@      @      @              @      @      1@                      �?              6@       @      ,@      &@      *@      �?      7@      0@      @      8@      @      0@              0@             �@@      $@      @      @      2@      *@      @      3@      2@     �H@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ 6jhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@Xd�e��@�	           ��@       	                   �0@oa_�B0@p           �@                            @�<0/
@z            @h@                           �? �}ן	@]            �a@������������������������       �>��_�@
             0@������������������������       ����Y��@S            �_@                           @v���j�	@            �I@������������������������       �pL�/�@            �B@������������������������       ���`��� @	             ,@
                            �?P��b�j@�           �@                           �?m���@�           ��@������������������������       �jѮ���
@�            �s@������������������������       ��2<�I�@�            `w@                          �2@�dV>�@H           `�@������������������������       �%��DL@�             w@������������������������       ��z��h@_            @c@                          �9@ ����b@-           ��@                           �?���@9           ��@                           @XO3L�@�           ��@������������������������       ��׹��@           �|@������������������������       �E�)�7@�             s@                           @f�e�d@N           H�@������������������������       ��XP��I@a           ��@������������������������       �nl&�<&@�             w@                            �?M�R�@�           ��@                           �?mh:#�%@�            `l@������������������������       �s�I��@5            @U@������������������������       �s�|���@R            �a@                          �?@��6a��@m           ��@������������������������       �(��E@-           �|@������������������������       �g���@@            @[@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       u@      _@     �Y@     @t@     �A@     @~@      .@     �j@      >@     �{@     @Y@     �P@     �B@     �O@     �n@     �Q@     �x@     �s@     �z@      V@      V@      6@      B@     �_@      "@     �k@      @      S@      @     �g@      ?@      <@      @      "@     �T@      3@     @b@     @X@     `h@      5@      *@              @      1@             �D@      @      (@              =@       @                      �?      *@              ,@      (@      @@              "@               @      ,@              >@              "@              2@                              �?      &@              (@      &@      :@              @                      �?              �?              �?              @                              �?      �?                              @              @               @      *@              =@               @              .@                                      $@              (@      &@      6@              @               @      @              &@      @      @              &@       @                               @               @      �?      @               @                       @              @      @       @              &@       @                               @               @      �?      @               @               @      �?              @              �?                                                                                      �?             �R@      6@      @@     @[@      "@     �f@              P@      @     �c@      =@      <@      @       @     @Q@      3@     �`@     @U@     `d@      5@      =@      0@      3@     �Q@      �?      X@              6@      @      ]@      ,@      3@      @      @     �B@      $@     �S@     �D@      Y@      *@      ,@       @      @      <@      �?      I@              @              R@      @      @      �?              1@       @      C@      1@     �F@      @      .@       @      (@      E@              G@              .@      @      F@      &@      0@       @      @      4@       @      D@      8@     �K@      @      G@      @      *@     �C@       @     �U@              E@             �E@      .@      "@      @      @      @@      "@      K@      F@     �O@       @      @@      @      "@      ;@       @     �O@              >@             �A@       @      @      @       @      4@       @      A@      @@      G@       @      ,@      �?      @      (@              7@              (@               @      *@      @               @      (@      �?      4@      (@      1@              o@     �Y@     �P@     �h@      :@     Pp@      &@     `a@      9@     �o@     �Q@      C@      ?@      K@     `d@     �I@     �n@      k@     `m@     �P@     `d@     @Q@      J@      a@      *@     @g@       @     @S@      3@      h@     �I@      4@      .@     �C@     @Y@      @@     @g@     �c@     �b@     �E@      M@      @@      ?@     �M@      &@      P@       @     �L@      *@     @T@      6@      .@      "@      =@     �B@      0@      Q@     @R@      O@      ;@      ;@      *@      4@     �D@      @     �H@       @      E@      @     �G@      3@      $@      �?      6@      5@      (@      A@      D@      <@      5@      ?@      3@      &@      2@      @      .@              .@      @      A@      @      @       @      @      0@      @      A@     �@@      A@      @     @Z@     �B@      5@     @S@       @     �^@              4@      @      \@      =@      @      @      $@      P@      0@     �]@      U@     �U@      0@     �R@      4@      (@      B@       @     @T@              .@       @      T@      0@      �?       @       @     �@@       @     @S@     �G@      J@      *@      ?@      1@      "@     �D@             �D@              @      @      @@      *@      @      @       @      ?@      ,@     �D@     �B@     �A@      @     �U@     �@@      ,@      O@      *@     �R@      "@      O@      @     �N@      3@      2@      0@      .@      O@      3@      N@     �M@     �U@      8@      0@      @      @      3@      @      @@              5@              3@      �?              @      @      2@      @      2@      4@      7@      "@      @              �?       @      @      *@              @              &@                      @      @      *@      @      @      @      @       @      "@      @      @      &@              3@              1@               @      �?              @      @      @              ,@      .@      4@      @     �Q@      <@      "@     �E@      "@     �E@      "@     �D@      @      E@      2@      2@      $@       @      F@      .@      E@     �C@     �O@      .@      N@      2@      @     �D@      @     �A@      @     �C@      @     �A@      .@      ,@      @      @      D@      *@      <@      :@      M@       @      $@      $@      @       @       @       @      @       @              @      @      @      @      @      @       @      ,@      *@      @      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�z5hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����@�	           ��@       	                    �?���e��@           ��@                          �:@} ���@h           @�@                           @�?��|@1           @}@������������������������       ���y�@�            �v@������������������������       ��\zo:@I            �Z@                           �?q@��@7             U@������������������������       ��un�@             9@������������������������       �0��U_@(            �M@
                           �?c��q�@�           �@                            �?pJ:��1@�            �v@������������������������       �� �|	�@B             [@������������������������       ��W{�H�@�            �o@                          �?@DxyT,&@�           ��@������������������������       �����@�           p�@������������������������       ��R�Y@&            �P@                           �?��S>B@�           ʡ@                          �;@�z�k?@/           Ћ@                            @-�oa��@           p�@������������������������       �H�KyL)@�           ��@������������������������       �x�)?Y�@i             f@                            �?e$L�@             F@������������������������       ���w��@             @@������������������������       �	4%'V@
             (@                           @|���b�@n           ��@                          �3@�K�rc�@�           ��@������������������������       ��x���/@�            �i@������������������������       �� 8�o(@           y@                           @���3�#@�           `�@������������������������       �mt�@�            �q@������������������������       �Gw-@<           �~@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@     �`@      S@     �v@      G@     �~@      @     �m@      1@     }@     �X@     �Q@     �C@      P@     �k@     �S@     �u@     �q@     �z@     �V@     �a@     �Q@      K@     �b@     �@@     �b@      @     �`@      &@      b@     �G@     �E@      2@      C@      V@     �B@     �_@     �a@     @c@      I@      H@      6@      3@     �M@      @     �P@      �?     �E@      @     �G@      *@      &@      @      $@      ;@      *@      <@      C@      S@      3@      D@      .@      1@     �M@      @      K@             �A@      @      D@      "@      @      �?       @      :@      (@      7@      A@      P@      .@      @@      @      *@     �H@      @     �H@              =@      @      >@       @      @              @      1@      $@      1@      1@     �I@      .@       @      $@      @      $@      �?      @              @              $@      �?              �?      @      "@       @      @      1@      *@               @      @       @                      (@      �?       @              @      @      @       @       @      �?      �?      @      @      (@      @      @               @                      @              @              @                      �?       @              �?                      @              @      @                              "@      �?      @              @      @      @      �?              �?              @      @      "@      @      W@      H@     �A@     �V@      =@      U@      @      W@      @     �X@      A@      @@      .@      <@     �N@      8@     �X@     �Y@     �S@      ?@     �B@      @      "@      .@      $@     �@@       @     �E@       @      ?@      (@      @      @      @      2@       @     �G@     �@@      ;@      "@      @      @       @      @      @      *@       @      9@              ,@                       @       @       @       @       @      @      @      @     �@@      �?      @      (@      @      4@              2@       @      1@      (@      @      @      @      $@      @     �C@      <@      5@      @     �K@     �D@      :@     �R@      3@     �I@      @     �H@      @     �P@      6@      :@       @      5@     �E@      0@     �I@     �Q@     �I@      6@     �F@      >@      6@     �P@      1@     �H@      @      G@      @      M@      5@      :@      @      4@      E@      .@     �I@     �O@      I@      5@      $@      &@      @       @       @       @              @              "@      �?              @      �?      �?      �?              @      �?      �?     `j@      P@      6@     @k@      *@      u@             �Y@      @      t@      J@      ;@      5@      :@     �`@      E@     �k@      b@     0q@      D@     �T@      "@      $@      R@      @     �b@              E@      �?     @`@      .@      @       @      $@      F@      (@     �V@     �M@     @_@      9@     �R@      "@      @      R@      @     @b@              E@      �?      _@      .@      @               @     �D@       @     @V@     �L@     �]@      7@      N@      "@      @     �J@      @     �]@              @@      �?     �X@      @      @              @      ?@      @     �R@     �H@     �Z@      (@      .@               @      3@      @      ;@              $@              :@      $@                      @      $@      @      .@       @      *@      &@      @              @                      @                              @               @       @       @      @      @      �?       @      @       @      @              @                      @                              @               @               @      �?      @                      @                                                                                                               @               @      �?      �?       @       @       @      `@     �K@      (@     @b@      @     �g@              N@      @     �g@     �B@      6@      3@      0@     �V@      >@     ``@     @U@     �b@      .@      I@      =@       @     �O@       @      Q@             �@@              Y@      3@      @      $@      $@     �D@      2@     �N@     �C@      F@      @      $@      @      @      ;@              (@               @              F@      @                      @      .@      @      =@      0@      8@      �?      D@      :@      @      B@       @      L@              9@              L@      .@      @      $@      @      :@      .@      @@      7@      4@      @     �S@      :@      @     �T@      @      ^@              ;@      @     �V@      2@      1@      "@      @      I@      (@     �Q@      G@     �Z@       @      0@      @      �?      C@      �?     @P@              $@      @      3@      @       @       @              ,@      &@      9@      0@      G@       @     �O@      5@      @     �F@      @     �K@              1@      �?     �Q@      ,@      "@      @      @      B@      �?     �F@      >@      N@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ(�ohG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?B�.�@�	           ��@       	                    �?e���@�           0�@                           @��I�:@W           ��@                           @ퟬ�?A@           �z@������������������������       ����m*@�            �p@������������������������       �I� @k            �d@                           �?��1%�@B            @X@������������������������       ��a�1�@             :@������������������������       �D�+g@2            �Q@
                           �?n�.v:@�           �@                          �9@�2 �e�@�             x@������������������������       ��C9�j�@�            �r@������������������������       �Iæ��@:             U@                          �:@~��K@�           ��@������������������������       �'�.'K@G           H�@������������������������       ���[�@q            `f@                           @w�5̜7@�           ��@                          �2@�Ș33@!           f�@                           @�1�L
U@�           ��@������������������������       �hgG���
@           P|@������������������������       ��o�B@�
@�            �p@                           �?������@\           ��@������������������������       � b����@�           �@������������������������       ���B�Ȉ@�           ��@                          �4@K��D�@�            @i@                          �3@�I��)�	@>             X@������������������������       ���Y�<$	@/            @Q@������������������������       �?��w�@             ;@                           @�B���Z@F            �Z@������������������������       �Ū�h@,            @R@������������������������       ���X��@            �@@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       0t@     `a@     �T@     v@     �@@     @~@       @     �n@     �@@     �|@     �W@      O@     �A@      O@     �n@     �R@     w@     @r@     �{@     �S@     �^@      Q@      M@     �a@      5@     �a@      @     �`@      9@     `a@      G@      C@      2@      G@     �Y@      C@     �`@      _@     �e@      B@     �F@      2@      <@     �G@      @      L@      �?      ?@      "@     �I@      1@      "@      @      @     �A@      (@     �F@      @@     �P@      $@     �D@      (@      5@     �E@      @      G@      �?      ;@      "@     �C@      0@      "@      @       @      @@      (@      @@      7@     �H@      $@      :@      "@      ,@      9@      �?     �@@              1@      "@      6@      *@      @      @       @      1@      $@      0@      $@      =@       @      .@      @      @      2@       @      *@      �?      $@              1@      @      @                      .@       @      0@      *@      4@       @      @      @      @      @              $@              @              (@      �?               @      @      @              *@      "@      1@                      �?      @      �?              @                               @                              �?       @              @      @      �?              @      @      �?      @              @              @              $@      �?               @      @      �?              $@      @      0@             @S@      I@      >@      X@      2@     �U@      @     @Y@      0@      V@      =@      =@      (@     �C@     �P@      :@     �V@      W@     �Z@      :@      =@      ,@      (@     �@@       @      @@              F@      @      C@      &@      &@       @      &@      .@      @      B@      F@      B@      @      <@      &@      @      8@      �?      =@              D@              A@      @      @              &@      &@      @      =@      ;@      =@      @      �?      @      @      "@      �?      @              @      @      @      @      @       @              @       @      @      1@      @              H@      B@      2@     �O@      0@      K@      @     �L@      (@      I@      2@      2@      $@      <@      J@      5@      K@      H@     �Q@      5@     �A@      3@      $@      F@      .@      J@      @     �A@      (@     �B@      1@      ,@      @      8@      A@      &@      G@      B@      I@      4@      *@      1@       @      3@      �?       @              6@              *@      �?      @      @      @      2@      $@       @      (@      5@      �?      i@     �Q@      8@     @j@      (@     `u@       @     @\@       @      t@      H@      8@      1@      0@      b@      B@     @m@      e@     �p@     �E@      f@     @P@      7@      i@      (@     �s@       @     @Z@       @     �r@     �C@      7@      &@      0@     �^@     �A@      j@     �b@     @o@     �E@     �H@      4@      @     @R@      �?     �Z@             �G@             �`@      @       @      @      @      9@      @      R@      J@     @Z@      $@      @@      @      �?     �L@      �?     �Q@              9@              S@      @      @      �?      @      (@      @      J@      4@      R@      @      1@      *@      @      0@              B@              6@              L@       @      �?       @              *@              4@      @@     �@@      @     �_@     �F@      3@      `@      &@     �i@       @      M@       @     �d@      A@      .@       @      *@     @X@      =@      a@     �X@      b@     �@@     �P@      2@      @      P@      $@     �\@       @     �A@      @      U@      6@      @      @      @      H@      (@     �E@     �F@     @Q@      1@      N@      ;@      .@      P@      �?      W@              7@       @      T@      (@      &@      @      @     �H@      1@     �W@     �J@      S@      0@      9@      @      �?      "@              =@               @              8@      "@      �?      @              7@      �?      9@      2@      1@              @                      @              2@              @              $@              �?      @               @      �?      4@      $@       @              @                      @              ,@              @              "@                                       @      �?      "@      @      @              �?                                      @                              �?              �?      @                              &@      @      �?              2@      @      �?      @              &@              @              ,@      "@              @              .@              @       @      "@              ,@      @      �?                       @              @              @      "@              @               @              @      @      @              @      �?              @              @                               @                                      @              �?       @      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJuPp!hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@����@�	           ��@       	                    @�*,���@           �@                           �?��hw�@           ܒ@                           �?�Vaʔ@           �y@������������������������       �t����d@�            �q@������������������������       �����	@Y            @`@                            �?��ڬ�@            Ј@������������������������       �N?"��c@           �z@������������������������       �R��·@�            �v@
                           �?�*_l��@            @�@                          �1@�Eb @&            ~@������������������������       ��D+ �@`            �c@������������������������       ����@�            @t@                           @#	���@�           p�@������������������������       ����;G@*           �}@������������������������       ��ܻX��
@�             q@                            @H	뭻@�           �@                          �?@ʀ��0@�           �@                           �?p���@f           ��@������������������������       �;�T�o@            x@������������������������       ��ɝ�Pv@b           ��@                           �?�}"�m@3             U@������������������������       �~w`�!�@             K@������������������������       ���Kv>�@             >@                           @�j_�A@'           �{@                           �?F�7���@           `x@������������������������       ��EgRI@V            �`@������������������������       ��jN�j@�             p@                          �<@#�ۅ&@$             L@������������������������       �H�~���@            �E@������������������������       �XL��J@             *@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �^@     �S@     �u@      F@     p@      "@     `o@      <@     pz@     �\@     �O@      ;@     �S@      j@     �O@     �w@      t@     `{@      S@     `g@      K@     �B@      m@      7@     �x@      @      c@      ,@     pp@      I@     �F@      $@      B@     @_@      =@     �n@      h@     s@     �B@     �X@      =@      <@      [@      3@     @b@      @     �T@       @     �_@      B@      :@      @      =@      N@      9@      ^@     �Z@     @^@      9@      B@      $@      @     �@@      @     �N@             �@@      �?     �L@      @      @       @      (@      3@      �?     �B@      >@     �J@      @      =@      "@      @      2@      @     �D@              :@      �?      @@      @      @       @      (@      0@      �?      :@      0@     �A@              @      �?              .@              4@              @              9@       @                              @              &@      ,@      2@      @     �O@      3@      5@     �R@      .@     @U@      @      I@      @     �Q@      =@      7@      @      1@     �D@      8@     �T@     @S@      Q@      2@      9@      "@      *@     �H@             �D@      @      6@      @     �A@      "@      .@      @      &@      2@      3@     �H@      D@     �E@      .@      C@      $@       @      :@      .@      F@      �?      <@             �A@      4@       @              @      7@      @      A@     �B@      9@      @      V@      9@      "@      _@      @     `o@             �Q@      @      a@      ,@      3@      @      @     @P@      @     @_@     �U@      g@      (@      A@      @       @      E@      @      [@             �A@       @      H@       @      @              @      @@              D@     �C@      R@      @                      �?       @      @      D@              "@              ;@              �?              @      $@              $@      *@      >@      @      A@      @      �?      A@              Q@              :@       @      5@       @      @              @      6@              >@      :@      E@      @      K@      3@      @     �T@      �?     �a@             �A@      @      V@      (@      .@      @             �@@      @     @U@     �G@      \@      @      <@      "@      @      P@      �?     �R@              8@             �N@      $@      $@      @              2@      @     �I@      8@     @V@      @      :@      $@       @      2@             @Q@              &@      @      ;@       @      @                      .@      �?      A@      7@      7@       @     �a@     @Q@     �D@     �]@      5@     �Z@      @     �X@      ,@      d@     @P@      2@      1@     �E@      U@      A@     @a@      `@     �`@     �C@     �Y@     �H@      8@     �V@      .@      V@      @     �L@      @     �^@     �C@      "@       @      8@     �O@      8@     �Y@     �S@     �Y@      5@     �X@      C@      5@     �U@      .@     �T@       @     �J@      @     �]@      B@       @      @      2@     �N@      6@     �W@      S@     �U@      .@      D@      (@       @      D@      (@     �@@       @      1@      @      M@      3@      �?       @      @      >@      @      @@     �@@      9@      "@     �M@      :@      *@      G@      @     �H@              B@             �N@      1@      @      @      .@      ?@      3@      O@     �E@      O@      @      @      &@      @      @              @      �?      @              @      @      �?      �?      @       @       @       @      @      .@      @              &@      @      @              @              @               @              �?      �?      @       @       @       @       @      @      @      @                                      �?      �?                       @      @                      @                      @      �?       @      �?     �C@      4@      1@      <@      @      2@       @     �D@      "@     �B@      :@      "@      "@      3@      5@      $@      B@      I@      ?@      2@     �@@      ,@      0@      :@              .@       @      D@      "@      A@      6@      @      @      .@      1@      @      ?@      H@      >@      2@      2@       @      @      "@              �?              (@              *@       @      @       @       @      @      @      (@      6@      (@      @      .@      @      (@      1@              ,@       @      <@      "@      5@      4@      @      @      *@      ,@      @      3@      :@      2@      (@      @      @      �?       @      @      @              �?              @      @      @       @      @      @      @      @       @      �?              @      @      �?       @      @      @              �?              @              @       @      @       @      @       @      �?                               @                                                                      @                               @              @      �?      �?        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�'?hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @F^衖�@�	           ��@       	                    �?\�=e�@           "�@                          �6@�N��@*           ș@                          �4@��1v�@*           �@������������������������       �x���ǁ@�           @�@������������������������       ��nx+`�@�             o@                           @��c�tW@            ��@������������������������       ��/>�r@^           ��@������������������������       ��e��@�            �o@
                          �5@g$�2�^@U           ��@                           �?�ҟA@�            @r@������������������������       �(�t!�@S            �`@������������������������       ���x>�@b             d@                            �?yX|�ג@�            `o@������������������������       ����@]             c@������������������������       �Whf��T@C            �X@                           @�'�L�@1           ��@                           @nn��@�            �x@                          �5@U[�sU;@�            Pv@������������������������       ���K�ӛ@�            @k@������������������������       �C��6@W            `a@                          �9@���R��@             B@������������������������       ���q�@             <@������������������������       �      @              @                           �?�x��r@2           ��@                          �2@_3]�@�           @�@������������������������       �1W�`}o
@�            �p@������������������������       ��� �b�@�             x@                          �7@X���@�           8�@������������������������       ��<s,�@3           �@������������������������       �x�e�j�@e             e@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       `r@     �`@     �R@     `u@      C@     x�@      "@     �i@     �@@     �|@     �Z@      N@     �C@     @R@     pp@     @P@     �w@     `s@     @y@     @X@     @e@      V@     �L@     @h@      @@     �j@      "@     �`@      ;@     �l@      R@     �B@     �@@      I@     �b@     �H@     �h@     @g@     `h@     �P@     @]@     @P@     �J@     �a@      >@      c@      "@     �Y@      9@     �d@     �H@      @@      5@      G@     @[@     �@@      c@     �a@     �b@     �K@     @Q@      ?@      <@      U@      &@     �\@      @      B@      &@     �V@      5@      2@      @      (@     �E@      .@     @S@     �S@      W@      ;@     �L@      .@      6@     @P@      "@     �R@      �?      :@      @      M@      (@      &@      @      @     �A@      "@      G@     �L@     �S@      9@      (@      0@      @      3@       @     �C@       @      $@      @     �@@      "@      @              @       @      @      ?@      5@      *@       @      H@      A@      9@     �M@      3@      C@      @     �P@      ,@     �R@      <@      ,@      1@      A@     �P@      2@      S@     �O@     �L@      <@     �A@      4@      5@      C@      $@      6@      @     �G@      ,@     �E@      ;@      (@      *@      3@      F@      &@      I@      I@     �@@      2@      *@      ,@      @      5@      "@      0@              4@              ?@      �?       @      @      .@      6@      @      :@      *@      8@      $@     �J@      7@      @     �I@       @     �O@              @@       @     @P@      7@      @      (@      @     �D@      0@      F@     �F@      G@      (@      .@      "@      �?     �@@              ?@              4@              D@      $@      @      @      �?      7@      @      A@      A@      5@      @      @      @              "@              (@              (@              9@       @              @               @       @      3@      ,@      "@       @       @      @      �?      8@              3@               @              .@       @      @       @      �?      .@      @      .@      4@      (@      �?      C@      ,@      @      2@       @      @@              (@       @      9@      *@       @      @      @      2@      "@      $@      &@      9@      "@      8@      "@              "@      �?      1@              @       @      1@      $@               @       @      *@      @      @      "@      8@      �?      ,@      @      @      "@      �?      .@              @               @      @       @      @      �?      @      @      @       @      �?       @      _@      G@      2@     �b@      @     �s@             �Q@      @     �l@      A@      7@      @      7@     @\@      0@     �f@      _@      j@      >@      9@      ,@      @      >@       @      P@              $@             @P@      @      @       @      @      3@       @     �N@      2@      C@      0@      7@      (@      @      >@       @      K@              @              P@       @      @      �?      @      2@      @      L@      2@      @@      0@       @      @      @      3@              A@              @              E@      �?      @      �?      �?      @      @      ?@      &@      9@      ,@      .@      @      @      &@       @      4@              �?              6@      �?                      @      *@              9@      @      @       @       @       @                              $@              @              �?      @      �?      �?              �?      �?      @              @               @      �?                              $@              �?              �?      �?      �?      �?              �?              @              @                      �?                                               @                       @                                      �?                       @             �X@      @@      (@     �]@      @      o@             �N@      @     �d@      =@      3@      @      1@     �W@       @      ^@     �Z@     `e@      ,@     �J@      0@      @     �O@      @      `@              9@       @     �S@      2@      @       @             �E@      �?      K@     �I@     �V@      "@      ,@      @              ;@       @      E@              .@             �B@      �?      @      �?              3@              >@      .@      I@      @     �C@      &@      @      B@       @     �U@              $@       @     �D@      1@      �?      �?              8@      �?      8@      B@     �D@      @      G@      0@      @     �K@             �]@              B@      @     �U@      &@      .@       @      1@     �I@      @     �P@     �K@      T@      @     �@@      "@       @     �E@             �X@              A@      @      T@      @      ,@       @       @      A@      @      H@      F@      I@      @      *@      @      @      (@              5@               @              @      @      �?              .@      1@       @      2@      &@      >@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��YhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @����h@�	           ��@       	                   �5@��1��@           X�@                           �?����@�           h�@                          �4@�����
@           �{@������������������������       ���3=46@�            �u@������������������������       ���t�
@4             W@                           @N1 �@u            �@������������������������       ��H�܃3@�             y@������������������������       ��Rww�3@}           p�@
                           �?o�mɲ@�           H�@                           @I�K���@           �z@������������������������       ������@�            0q@������������������������       �=��9
;@a             c@                           �?$�Ĳ�@�           8�@������������������������       �c�X>>�@�            w@������������������������       �eej;��@�            �n@                           @����@�           t�@                           @����a@"           �@                           �?�^��t>@           ��@������������������������       ��Mpxx�@�            �p@������������������������       �=y�=s@Y           p�@                           �?�<��
@             F@������������������������       ��� 8��@             &@������������������������       ��aK�)	@            �@@                            @��=�@           ؂@                          �6@r}�Լ@8           �~@������������������������       �8�� @�            pr@������������������������       �:|�`,�@y             h@                           @�W�
@G            �\@������������������������       ����0��	@&            �M@������������������������       �<b��N�	@!             L@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �[@      T@     �v@      B@      @      @      p@      8@     �{@      [@     @Q@      D@      L@     `m@      L@     �w@     Pt@      |@      Q@     �g@      O@      J@      j@      5@     v@      @     �d@      .@     @s@     �P@      ;@      2@      9@      c@      6@     �l@     �i@     pr@     �J@     @Y@      <@      ,@     `a@      $@     �k@       @     �V@      &@     @g@      9@      2@      (@      "@     �Q@      @     `b@     �Z@     �i@      @@      E@      @       @     �L@      "@      J@       @     �A@      $@      :@       @      @       @      @      7@       @     �H@     �A@     �K@       @      ;@      @       @      E@      "@     �G@       @      8@      @      6@       @      @       @      @      6@       @      =@      <@     �I@      @      .@      @              .@              @              &@      @      @              �?              �?      �?              4@      @      @       @     �M@      5@      @     �T@      �?      e@              L@      �?      d@      1@      &@      $@      @      H@      @     �X@      R@     �b@      8@      4@      "@      @      F@             �O@              0@              O@      &@      @       @       @      1@      @     �H@      =@      H@      2@     �C@      (@      @      C@      �?     @Z@              D@      �?     �X@      @      @       @       @      ?@       @     �H@     �E@     @Y@      @      V@      A@      C@     @Q@      &@     �`@      @      S@      @     �^@      E@      "@      @      0@     @T@      .@     @T@      Y@     �V@      5@     �B@      $@      "@      3@      @     �P@      @      C@      @     �N@      1@      @       @      @      :@      @      <@      G@      B@      @      9@      @      @      *@      @      E@      @      7@      @      B@      &@      @       @      @      0@              *@      B@      8@      @      (@      @      @      @              9@              .@      �?      9@      @                              $@      @      .@      $@      (@      �?     �I@      8@      =@      I@      @     �P@       @      C@             �N@      9@      @      @      (@     �K@      &@     �J@      K@     �K@      .@      8@      .@      ;@      A@      @     �@@       @      >@              @@      7@      @      @      $@      8@      &@      =@     �@@      7@       @      ;@      "@       @      0@       @     �@@               @              =@       @              �?       @      ?@              8@      5@      @@      @      _@     �H@      <@     �c@      .@     �a@             @V@      "@     �`@     �D@      E@      6@      ?@     �T@      A@     �b@     �]@      c@      .@     @R@      >@      3@      X@      .@      M@             �L@      @      T@      7@      9@      0@      ,@     �L@      5@     �T@     �R@     �R@      (@     �Q@      ;@      3@     �W@       @      M@             �I@      @     @S@      6@      9@      ,@      ,@      K@      4@     �R@     �Q@     @R@      (@     �C@      @      (@      ?@      @      1@              1@       @      2@      "@      @      @      @      3@      @      3@      7@      <@      @      ?@      6@      @      P@      @     �D@              A@      @     �M@      *@      5@      &@      &@     �A@      *@     �K@     �G@     �F@       @      @      @              �?      @                      @              @      �?               @              @      �?      "@      @      �?              @                                                       @                      �?                               @              @                                      @              �?      @                      @              @                       @              �?      �?      @      @      �?             �I@      3@      "@     �N@             @U@              @@       @     �K@      2@      1@      @      1@      :@      *@     �P@      F@     �S@      @     �C@      3@      @     �I@              R@              ;@       @     �A@      .@      &@      @      0@      9@      &@     �I@      C@      P@       @      1@      ,@      @      ?@             �M@              ,@      �?      7@       @      &@      �?      �?      *@              ?@      8@     �D@       @      6@      @      @      4@              *@              *@      �?      (@      @               @      .@      (@      &@      4@      ,@      7@              (@               @      $@              *@              @              4@      @      @      @      �?      �?       @      .@      @      .@      �?       @               @       @              $@              @              "@      @      �?                               @      &@       @      @              @                       @              @                              &@              @      @      �?      �?              @      @      &@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJwB$hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�� 3��@�	           ��@       	                     @�q�d��@�           �@                           �?L{C�$@b           ��@                          �5@��h�N@=           �}@������������������������       �{�����@            y@������������������������       ��~4m@0            �R@                           �?~�B�D@%           ,�@������������������������       �����Q�	@+            @������������������������       �����5@�           ؈@
                          �4@�*|
=<@�           ��@                           @�n�&@-           �@������������������������       �VO��`@�            �z@������������������������       ���s	@4            �T@                           �?f.�Z�@d             c@������������������������       �O#Q��@,            �P@������������������������       �4QQ4�@8            �U@                           �?�� 轋@�           D�@                          �:@�i6?@�           �@                           �?��&�
T@           �{@������������������������       ���l��@U            @`@������������������������       ��iF�A@�            `s@                            @��7`�/@�            Pt@������������������������       ����o{�@}             i@������������������������       �z��?A�@O            @_@                           @|�k˨@�           ��@                          �<@��@;Y@B           �@������������������������       �|�G*��@           0z@������������������������       ��mI�@:            �W@                            @a>k���@�            @j@������������������������       ��
��z2@n            �f@������������������������       ���Pa>�@             >@�t�b��     h�h5h8K ��h:��R�(KKKK��h��B`       �t@      [@     �U@     �t@      B@     P~@      @     �l@      >@     �}@     �\@     �N@     �C@     @P@     `l@     @R@     �v@     �t@     �{@     @T@     �f@     �L@     �E@     �j@      ;@     �v@             �`@      .@     �s@      L@      C@      1@      7@     @`@      @@     @n@      g@     @s@     �F@     @]@     �B@      7@     �e@      .@     @q@              V@      *@     �m@     �C@      >@      .@      *@      W@      6@     �e@     �\@     �o@      >@     �G@      $@       @     �O@      @     �K@              5@      $@      F@      @      .@      �?      &@      8@       @     �A@      <@     @P@      2@      C@       @      @      N@      @     �C@              3@      @     �D@      @      ,@              @      8@      �?      @@      <@      I@      2@      "@       @       @      @      �?      0@               @      @      @       @      �?      �?      @              @      @              .@             �Q@      ;@      .@      \@      &@     �k@             �P@      @     `h@      @@      .@      ,@       @      Q@      ,@      a@     �U@     �g@      (@      =@      �?      �?      F@       @     @Y@              ;@       @      T@       @       @      �?              :@      @      K@      <@     @U@      @     �D@      :@      ,@      Q@      "@      ^@              D@      �?     �\@      >@      *@      *@       @      E@      $@     �T@      M@     @Z@      @     �O@      4@      4@     �C@      (@      V@             �F@       @     @S@      1@       @       @      $@      C@      $@     �Q@     �Q@     �J@      .@     �J@      &@      ,@      =@      $@     �Q@              =@       @     �O@      *@      @       @      @      =@      $@     �F@      J@     �H@      ,@      I@      $@      *@      7@      $@      J@              0@       @     �H@      *@      @       @      @      <@      $@      E@     �F@      C@      *@      @      �?      �?      @              2@              *@              ,@                              @      �?              @      @      &@      �?      $@      "@      @      $@       @      2@              0@              ,@      @      @              @      "@              9@      2@      @      �?      @               @      @       @      @               @              @       @      @              �?      @              @      &@      @              @      "@      @      @              &@               @              "@       @                       @      @              4@      @      �?      �?     �b@     �I@      F@     �\@      "@     @^@      @     �W@      .@     �c@     �M@      7@      6@      E@     @X@     �D@     @_@     `b@      a@      B@     �I@      =@      @@      N@      @     �J@       @     @P@      (@      K@      =@      1@      2@      :@     �E@      ;@     �S@     @Q@      P@      =@      >@       @      1@      =@      @      C@              >@      @     �E@      2@      @      @      5@      ?@      "@     �N@      @@     �A@      5@      @              @      $@      @      &@              @       @      .@      @      @              �?      ,@      �?      1@      *@      *@      @      7@       @      $@      3@      �?      ;@              7@      @      <@      .@      �?      @      4@      1@       @      F@      3@      6@      2@      5@      5@      .@      ?@      @      .@       @     �A@      @      &@      &@      *@      .@      @      (@      2@      1@     �B@      =@       @      &@      ,@      @      1@              ,@       @      8@              $@      @      "@      "@      �?       @      (@      *@      2@      4@      @      $@      @       @      ,@      @      �?              &@      @      �?      @      @      @      @      @      @      @      3@      "@      @     �X@      6@      (@     �K@       @      Q@      �?      >@      @      Z@      >@      @      @      0@      K@      ,@     �G@     �S@     @R@      @     @Q@      @      "@      E@      �?     �O@      �?      1@       @     @S@      7@      @      @      *@     �B@      @      A@      I@     �G@      @      M@      @      @      B@             �M@              1@       @     �L@      1@      @      �?      (@      =@      �?      :@      F@      C@      @      &@      �?      @      @      �?      @      �?                      4@      @               @      �?       @      @       @      @      "@       @      =@      .@      @      *@      �?      @              *@      �?      ;@      @              �?      @      1@       @      *@      <@      :@              <@      ,@              &@      �?      @              (@      �?      .@      @                      @      0@      @      *@      ;@      6@              �?      �?      @       @              �?              �?              (@      �?              �?              �?      �?              �?      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�LthG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�c_��@�	           ��@       	                     @�σ1@           Й@                          �6@�O8J�k@e           ��@                          �4@]����@M           Ȁ@������������������������       �aF |.h@�            �w@������������������������       �w5�J@d            �c@                           �?n��P@           �{@������������������������       ��5jU��@U            �_@������������������������       ��^�2>N@�            �s@
                          �3@ν�]�@�           �@                           �?))ԥ%@~             j@������������������������       ��aM�=@A            @[@������������������������       �z�5�N@=            �X@                           �?҉�)<@1            }@������������������������       ��;u1��@@            �V@������������������������       �R�m�d=@�            �w@                           @��[I��@�           ��@                           �?�ь���@�           ��@                           @<
sZ?/@+           P�@������������������������       �d�:�M@�             n@������������������������       ��[G ��@�           Ѓ@                          �6@vc_��@t           ��@������������������������       ��֦U9@           py@������������������������       �Fi2~�@q             e@                            @���p�@           `�@                          �<@��T=�@�           (�@������������������������       ��`��@@w           �@������������������������       ��P1�@)             Q@                          �0@8����-@d            �d@������������������������       ��U��@             .@������������������������       ����S�@]             c@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@      b@      T@     `u@      F@     `}@      @     �l@     �@@      |@     @\@     �M@      @@      Q@      p@     �S@     �v@     �r@     @z@     �U@     �^@     �Q@     �K@     �b@      ?@      d@      @     @]@      6@     `a@      K@      =@      4@      E@      \@     �F@     `a@      b@      c@     �E@     �R@     �J@      8@     �[@      &@      Z@       @      L@      &@     �W@      3@      2@      $@      3@     @P@     �@@      S@     �Q@      Y@      <@     �G@      4@      *@     �R@      �?      S@              4@       @     �G@      "@      @       @       @      A@      $@      E@      B@      O@      5@     �@@       @      (@      L@             �G@              .@      �?      B@      "@      @      �?       @      ;@      @      8@      <@     �H@      2@      ,@      (@      �?      3@      �?      =@              @      @      &@                      �?      @      @      @      2@       @      *@      @      ;@     �@@      &@     �A@      $@      <@       @      B@      @      H@      $@      (@       @      &@      ?@      7@      A@      A@      C@      @      @      @      @      @      @      &@              @              5@      "@      @      @              @      @      &@      &@      &@      @      8@      :@      @      @@      @      1@       @      =@      @      ;@      �?      @      �?      &@      9@      4@      7@      7@      ;@       @     �H@      2@      ?@     �C@      4@      L@      @     �N@      &@      F@     �A@      &@      $@      7@     �G@      (@     �O@     �R@      J@      .@      (@      @      &@      *@      @      :@       @      2@              &@      "@      @      @              :@      @      6@      8@      .@      �?       @       @      @      "@              ,@              @              @      @              @              0@      �?      1@      (@      @              @       @      @      @      @      (@       @      *@              @      @      @                      $@       @      @      (@       @      �?     �B@      ,@      4@      :@      1@      >@      �?     �E@      &@     �@@      :@      @      @      7@      5@      "@     �D@      I@     �B@      ,@       @      @      @      �?       @      &@      �?      &@      @      @      �?      �?              �?       @      �?      .@      @       @      @      =@      &@      .@      9@      .@      3@              @@       @      ;@      9@      @      @      6@      3@       @      :@     �E@      =@      &@     @j@     �R@      9@      h@      *@     `s@      �?     �\@      &@     ps@     �M@      >@      (@      :@     @b@      A@      l@     �c@     �p@      F@     �a@     �B@      &@     @[@      @      k@             �S@      @      m@      B@      $@      @      *@     @X@      ,@      a@     @X@     �e@      =@     �U@      ,@      "@     �N@      @      b@             �D@       @     �`@      2@      @       @      $@      P@      @     �U@     �L@      \@      2@      8@      @              6@       @     �@@              ,@              F@       @      �?       @              1@      @      4@      &@      8@       @     �O@      @      "@     �C@       @     �[@              ;@       @     �V@      $@      @              $@     �G@       @     �P@      G@      V@      $@     �J@      7@       @      H@      �?     @R@              C@       @     �X@      2@      @      @      @     �@@      "@      I@      D@     �O@      &@      9@      &@       @      @@      �?      M@              ?@              R@       @      @      @              8@      @      F@      :@      I@       @      <@      (@              0@              .@              @       @      :@      $@       @              @      "@       @      @      ,@      *@      @     �Q@     �B@      ,@      U@       @     @W@      �?     �A@      @     �S@      7@      4@      @      *@     �H@      4@     �U@     �M@     @W@      .@      J@      <@      &@      R@       @     @S@      �?      8@      @      M@      5@      ,@      �?      &@      C@      ,@      L@      J@     @U@      .@     �F@      <@       @     �Q@      @      R@              4@      @      L@      0@      ,@      �?      @      C@      *@     �H@      H@     @Q@      (@      @              @       @      �?      @      �?      @               @      @                      @              �?      @      @      0@      @      2@      "@      @      (@              0@              &@              5@       @      @      @       @      &@      @      ?@      @       @              @      @       @      �?                              @                                                      �?                                              ,@      @      �?      &@              0@              @              5@       @      @      @       @      $@      @      ?@      @       @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ���ahG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @W���ӂ@�	           ��@       	                   �6@�0���@�            �@                          �4@%o�m��@h           `�@                            �?m�X��@H           $�@������������������������       �����:@�           `�@������������������������       �֘pb��
@�            s@                           �?Wύc2t@            �|@������������������������       ��Y���@,            �R@������������������������       ��0D��@�            @x@
                           @��$��@�           @�@                           �?"����@�           Ȅ@������������������������       �#U���@�            pq@������������������������       ���*B/V@�             x@                           �?����n�@�            �t@������������������������       �Z)k�@O            �^@������������������������       ��+�،@�            �j@                          �6@4Ɖ�m�@�           $�@                          �5@ �s�l�@�           ��@                           @����@T           �@������������������������       �
B��5�@           `|@������������������������       ��>�v��	@:             W@                           �?VK}��C@8             W@������������������������       ��ڇ+��@             &@������������������������       ��A����
@1            @T@                          @@@٧)p@'           �|@                           �?J����H@           �z@������������������������       ��,�|a,@N            �]@������������������������       �[ZH�$@�             s@                           @�,��Y
@            �A@������������������������       ��׋�@             7@������������������������       ��[���@
             (@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �]@     �V@     �u@     �I@     �@      @     �h@      A@     �|@     �Z@     �M@      B@     �N@      n@      K@     �y@     `r@     �z@      S@     �l@     @S@      I@     �p@      7@      y@      @     ``@      5@     @u@     �L@      F@      7@     �D@      g@     �B@     pr@     �j@     �t@      I@     @Z@      F@      9@     �e@      @     �s@      @     �T@      *@     �n@      ?@     �@@      $@      3@     @Z@      1@     `h@     @`@     `m@      :@     �T@      6@      3@     �`@      @     @m@             �M@      @      i@      6@      3@      @       @     �R@      &@     �a@     �X@     `h@      4@     �P@      1@      1@      \@       @     `c@             �D@      @     �d@      2@      ,@      @      @      K@      &@      \@     �U@     `b@      .@      .@      @       @      6@       @     �S@              2@              B@      @      @              @      5@              <@      (@      H@      @      7@      6@      @     �C@      @     �T@      @      8@      "@     �F@      "@      ,@      @      &@      >@      @     �K@      @@      D@      @      @      @      �?      @              .@      @      �?      @      @       @              �?      @              @      @       @      &@              2@      3@      @      @@      @     �P@              7@      @      E@      @      ,@      @       @      >@      �?     �I@      8@      =@      @     �_@     �@@      9@     �V@      0@      U@       @      H@       @     �W@      :@      &@      *@      6@     �S@      4@      Y@      U@     �W@      8@     �W@      7@      4@      J@      "@     @S@       @      ?@      @     �P@      0@       @      $@      @      I@      @     �Q@      H@     �J@      .@      <@      @      @      1@      @     �@@              (@              >@      "@      @      @      �?      ;@      �?     �C@      3@      7@      &@     �P@      0@      ,@     �A@      @      F@       @      3@      @      B@      @      @      @      @      7@      @      ?@      =@      >@      @      ?@      $@      @     �C@      @      @              1@       @      <@      $@      @      @      .@      =@      *@      >@      B@     �D@      "@      ,@              @      (@      @      @               @       @      &@      @              �?      �?      5@      @      (@      &@      @      @      1@      $@              ;@      @      @              .@              1@      @      @       @      ,@       @      @      2@      9@      A@      @     �X@      E@     �D@      U@      <@     �\@       @     �P@      *@      ^@     �H@      .@      *@      4@      L@      1@     �\@      T@     @X@      :@     �L@      9@      2@     �E@      .@     �U@              A@      @      V@      ;@      @      @       @     �A@       @     �T@     �F@     �K@      @     �I@      3@      .@     �B@      *@      S@              ?@      @      Q@      3@      @      @       @      <@      @     �Q@      E@     �K@       @     �G@      0@      &@      @@      *@     �M@              9@      @      H@      3@      @      @       @      3@      @      Q@      @@     �F@       @      @      @      @      @              1@              @              4@              �?                      "@              @      $@      $@              @      @      @      @       @      $@              @              4@       @       @                      @       @      (@      @               @               @              �?              �?                                               @                      @       @                                      @      @      @      @       @      "@              @              4@       @                              @              (@      @               @     �D@      1@      7@     �D@      *@      =@       @     �@@      $@      @@      6@       @      $@      2@      5@      "@      ?@     �A@      E@      6@     �D@      .@      2@      C@       @      =@       @      ?@      $@      @@      0@       @      @      .@      5@      "@      =@     �@@     �D@      6@      &@      @      "@       @      @      @              "@      @      ,@       @      @               @      �?      �?      @      (@      (@      @      >@      &@      "@      >@      @      7@       @      6@      @      2@      ,@      @      @      *@      4@       @      7@      5@      =@      1@               @      @      @      @                       @                      @              @      @                       @       @      �?                              @      �?      @                                              @              @      @                       @      �?                               @      �?       @                               @                      @                                                      �?      �?        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�g�qhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@jO9fH�@�	           ��@       	                     @ w�.�@n           ,�@                           @�Z���@D           ��@                           �?��e��@d           �@������������������������       �l��%@            �j@������������������������       ����5@�            �v@                          �0@k��m�
@�           ��@������������������������       ���� z@C             Z@������������������������       ����H:@�           ��@
                           �?Tr�7I�@*           �~@                           @���X@�            �p@������������������������       ��\g��@�            �n@������������������������       �� ���	@             6@                           @��8�{d@�            �k@������������������������       ��i��,P
@m            `f@������������������������       ��/g�B
@            �E@                          �6@Q�̥��@=           |�@                           �?�`X�r@�           �@                          �5@̂ə��@�            @m@������������������������       ����@�@N             a@������������������������       ���.�M@?            �X@                           @��AE��@           �w@������������������������       �5���@�            �i@������������������������       ��d#h@u            �e@                           @�����@�           p�@                           �?�eZ)X@�           �@������������������������       �!N�m}"@            �z@������������������������       ����d%@�           ؈@                          �8@IqP��@�            pq@������������������������       ��9-���@J            @^@������������������������       �a��rm�@l            �c@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       Ps@     �`@     �V@     �u@     �D@     �~@      @     �k@      B@     �|@     @[@      N@      =@      S@      k@      Q@     w@     `s@     0|@      T@     ``@      >@     �@@     �e@      0@     Pq@             @V@      0@     �o@      E@      <@      @      ,@     @T@      2@      g@     �a@     �m@     �@@     �T@      5@      4@      b@      @     �i@             �O@      (@      i@      6@      5@      @      "@      M@      "@     @a@     @X@     `e@      ?@     �H@      $@      0@     �U@      @     �O@              9@      $@     �Q@      (@      $@       @       @      6@      @     �H@     �I@      P@      4@      4@       @      @      :@       @      >@              &@              >@       @       @       @       @      @              .@      6@      >@      @      =@       @      "@      N@       @     �@@              ,@      $@     �D@      $@       @              @      0@      @      A@      =@      A@      .@      A@      &@      @      M@             �a@              C@       @      `@      $@      &@       @      �?      B@      @     @V@      G@     �Z@      &@      @      �?              @              8@                              8@               @                      @              "@      @      9@              >@      $@      @     �J@             �]@              C@       @     @Z@      $@      "@       @      �?      =@      @      T@     �E@     �T@      &@      H@      "@      *@      <@      (@      R@              :@      @     �J@      4@      @      �?      @      7@      "@     �G@      G@     �P@       @      9@      @      "@      *@      &@      >@              &@      @      2@      "@      @      �?      @      1@      @     �@@      >@     �B@      �?      5@       @      "@      $@      &@      ;@              $@      @      1@       @      @      �?      @      0@      @      =@      >@     �B@              @       @              @              @              �?              �?      �?                      �?      �?              @                      �?      7@      @      @      .@      �?      E@              .@             �A@      &@                              @      @      ,@      0@      =@      �?      3@       @      �?      (@      �?      E@              (@              =@      &@                              @       @      "@      *@      4@      �?      @      @      @      @                              @              @                                      �?      @      @      @      "@             @f@      Z@      M@     `f@      9@     �j@      @     �`@      4@     �i@     �P@      @@      8@      O@      a@      I@      g@     �d@     �j@     �G@     �I@      @@      5@      K@      @     �V@      �?      ?@      @     @P@      ,@      *@      @      1@     �D@       @     �Q@      D@      F@      @      7@      (@      "@      6@      �?      ?@      �?      0@              ,@      @       @              ,@      .@              :@      (@      8@      @      3@      @      @      5@              &@              @              @       @       @              @      @              1@      $@      2@      @      @       @      @      �?      �?      4@      �?      $@              "@      @                      @      "@              "@       @      @              <@      4@      (@      @@       @     �M@              .@      @     �I@      @      &@      @      @      :@       @     �F@      <@      4@              .@      @      $@      1@       @      ?@              $@      �?      :@      @       @      @      �?      .@      @      5@      2@      (@              *@      *@       @      .@              <@              @      @      9@      �?      "@               @      &@      �?      8@      $@       @             �_@      R@     �B@     @_@      6@     @_@      @     �Y@      ,@     �a@     �J@      3@      5@     �F@     �W@      E@     @\@     �_@     @e@      E@      V@     �N@      >@     �X@      5@     @X@      @     �Y@      ,@     �[@     �H@      .@      2@     �A@      S@     �D@      W@     �X@      `@      C@      9@      @      $@      @@      @     �E@             �D@      @      F@      0@      @      $@      $@      >@      "@      ?@     �G@      D@      4@     �O@      K@      4@     �P@      1@      K@      @     �N@      $@     �P@     �@@      (@       @      9@      G@      @@     �N@      J@     @V@      2@     �C@      &@      @      :@      �?      <@              �?              ?@      @      @      @      $@      3@      �?      5@      <@     �D@      @      $@      @      @      4@              ,@                              0@       @                       @      &@              @       @      *@      @      =@      @      @      @      �?      ,@              �?              .@       @      @      @       @       @      �?      ,@      4@      <@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��PhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���ּ@�	           ��@       	                    �?�`!�@           ��@                            �?��@_           ��@                           �?�"#V�@�            �u@������������������������       ��#�W�@J            @^@������������������������       �O]�}�@�            �k@                          �1@4S9P=�@�            �k@������������������������       ��Ү��X
@             ?@������������������������       �Ur@��@y            �g@
                            @C���-@�           ��@                           @J6&@h           ��@������������������������       ����)�@            Pz@������������������������       �'�e�H@h             f@                           �?�QN���@@           ��@������������������������       ��[�&v@y            @i@������������������������       ���"�@�            �t@                           �?���L@�           P�@                           @I&
@��@�           �@                          �4@� ��[�
@           �{@������������������������       � 0G>s�@�            �o@������������������������       ��K���@v            `g@                          �2@�Sg��@�            �r@������������������������       �w����	@H            �\@������������������������       �.&S-�x@{            �f@                           @ν���@�           �@                           @(HB��@;           �@������������������������       �`N���@�           `�@������������������������       �&��;�@�            Pq@                           �?�<k�#@j           (�@������������������������       ����$�@�            �q@������������������������       �Ǳ �C@�            �r@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       @u@      ]@     �\@     �t@     �G@     �}@      @     �n@      A@     �z@     �Z@     �P@     �J@      N@     @m@      J@     @w@     @t@      |@     �N@      c@     @Q@      R@     �a@      @@     @_@      @     @_@      9@     �d@      K@     �E@      >@      C@     �Y@      @@     �a@     �b@     �d@      =@      F@      0@      ;@      N@      @      H@       @      3@      @      N@      1@      &@      @      "@     �D@      ,@      C@      J@      S@      *@      9@      &@      5@      C@              <@      �?      ,@      �?      @@      @      @      @      @      =@      $@      ,@     �@@     �J@      "@      $@      �?      .@      $@              "@      �?      @              ,@      �?       @               @      $@      �?       @      ,@      4@      @      .@      $@      @      <@              3@               @      �?      2@      @      @      @      @      3@      "@      (@      3@     �@@      @      3@      @      @      6@      @      4@      �?      @      @      <@      $@      @              @      (@      @      8@      3@      7@      @                               @      �?      @                              @      @      �?              @      @      @               @       @              3@      @      @      4@       @      .@      �?      @      @      9@      @      @                      @      �?      8@      1@      5@      @      [@     �J@     �F@     �T@      =@     @S@      @     �Z@      2@     @Z@     �B@      @@      7@      =@      O@      2@      Z@     @X@      V@      0@      K@      D@      7@      J@      *@      D@       @      G@      &@      N@      .@      2@       @      *@     �B@      (@     �G@      H@      H@      $@      D@      ?@       @      B@      "@     �B@       @     �@@      "@      E@      .@      "@      @      @      =@      @      ?@      C@      <@       @      ,@      "@      .@      0@      @      @              *@       @      2@              "@      @      @       @      @      0@      $@      4@       @      K@      *@      6@      ?@      0@     �B@      �?      N@      @     �F@      6@      ,@      .@      0@      9@      @     �L@     �H@      D@      @      ,@      @      @      $@      @      2@              @@              ,@       @      @      @      $@       @      @      6@      5@      3@      @      D@      @      0@      5@      *@      3@      �?      <@      @      ?@      4@      "@      (@      @      1@      �?     �A@      <@      5@      @     �g@     �G@      E@      h@      .@     �u@      �?      ^@      "@     @p@      J@      8@      7@      6@     ``@      4@     �l@     �e@     �q@      @@      O@      @      &@      K@      &@     @`@             �G@             �V@      &@      @              @     �H@              U@      G@     �\@      (@     �@@      @       @      @@       @      W@              2@             �P@      @      @              �?      @@             �F@      8@     �O@      @      .@      @              6@      �?      O@              @              F@      @                      �?      0@              2@      .@     �E@      �?      2@               @      $@      @      >@              &@              7@      @      @                      0@              ;@      "@      4@      @      =@       @      "@      6@      @      C@              =@              7@      @                      @      1@             �C@      6@     �I@      @      @              @       @      @      1@              4@              $@                              @       @              0@      "@      6@       @      8@       @      @      4@              5@              "@              *@      @                      �?      .@              7@      *@      =@      @     �_@      D@      ?@     @a@      @      k@      �?     @R@      "@     @e@     �D@      3@      7@      1@     �T@      4@     @b@      `@     �e@      4@     �M@      <@      0@     �U@       @     �b@             �H@      "@     �V@      >@      &@      *@      $@     �F@      4@     @U@      S@     �Z@      $@      E@      :@      .@     @Q@      �?     @V@              <@             @Q@      5@      @       @      @      B@      &@     �N@      L@     �P@      $@      1@       @      �?      1@      �?      O@              5@      "@      5@      "@      @      @      @      "@      "@      8@      4@     �D@             �P@      (@      .@      J@       @     �P@      �?      8@              T@      &@       @      $@      @     �B@             �N@     �J@     @P@      $@      B@      @      @      C@       @     �@@      �?      3@              B@       @               @              2@              =@      <@      <@      �?      ?@      "@      (@      ,@             �@@              @              F@      @       @       @      @      3@              @@      9@     �B@      "@�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJG0� hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?E�C�@�	           ��@       	                    �?w�DL�@�           4�@                          �:@๑�_@d           �@                          �5@	t��@/           �|@������������������������       ��ʴտ@�            @q@������������������������       ��k�t�@w            @g@                           @XU�kU�@5             U@������������������������       ��u�D7@              J@������������������������       �nܯO�@             @@
                           �?�Wn�%@�           ��@                          �;@g�[�.@�            �w@������������������������       ��F���@�            �r@������������������������       ���0a��@+            @S@                          �:@�q��vJ@�           ��@������������������������       ��`�z$U@@            @������������������������       �V�v��@u             h@                           @�|���F@�           ��@                          �8@�6�S�@8           d�@                           @����@�           \�@������������������������       �w�@�           ��@������������������������       �|yx�~4@�             p@                           �?g-�`��@�             p@������������������������       ��� Np@2            �V@������������������������       �z�	\E@k             e@                           @ۥ��j@a           �@                          �2@]U��b�@W            `a@������������������������       ��[�Q@1            �R@������������������������       �H�@
@&             P@                          �3@�%2U]�@
           ��@������������������������       ����y&�
@�            �x@������������������������       ���e~�f@           �|@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       t@      `@     @Y@     `v@     �H@     �|@      @     @k@      :@     �{@     �[@     �M@      K@      P@     �l@     �S@     �v@     �s@     �|@     @S@     @_@     @P@     @P@     �^@      A@     @`@      @     @_@      5@     �`@     �N@      ?@     �@@      E@      W@     �@@      c@      b@     @c@      G@      H@      7@      :@      B@      @     �N@      �?      @@      @     �F@      5@      @      @      @      @@      .@     �E@      D@     @Q@      ;@     �D@      2@      5@      B@      @     �J@              7@      @     �@@      3@      @      @      @      ?@      ,@     �D@     �C@      K@      3@      @@      "@      @      9@      @      ?@              @       @      :@      "@      @               @      (@      @      4@      ;@      D@      *@      "@      "@      ,@      &@      �?      6@              0@      �?      @      $@      �?      @       @      3@       @      5@      (@      ,@      @      @      @      @                       @      �?      "@              (@       @      �?      @      @      �?      �?       @      �?      .@       @      @       @      @                       @      �?       @               @       @      �?      @              �?      �?       @              @       @      �?      @       @                      @              �?              @                              @                              �?      &@             @S@      E@     �C@     �U@      =@     @Q@       @     @W@      2@     �V@      D@      9@      ;@     �A@      N@      2@     @[@      Z@     @U@      3@      @@      @      *@      <@       @      6@             �E@      @      ?@      0@      @      *@      @      3@      @     �G@      @@      C@      @      =@      @      @      7@      @      6@             �A@      @      >@      $@      @       @      @      *@             �D@      8@      B@      @      @       @       @      @       @                       @      �?      �?      @              &@              @      @      @       @       @      @     �F@     �B@      :@      M@      5@     �G@       @      I@      ,@     �M@      8@      3@      ,@      <@     �D@      *@      O@      R@     �G@      (@      =@      0@      3@      A@      2@     �F@       @     �@@      ,@     �I@      6@      *@      $@      9@     �@@      @      G@     �C@     �@@      "@      0@      5@      @      8@      @       @              1@               @       @      @      @      @       @      @      0@     �@@      ,@      @     �h@     �O@      B@     �m@      .@     �t@             @W@      @     Ps@      I@      <@      5@      6@      a@      G@      j@      e@     �r@      ?@     �Z@     �E@      0@     �a@      &@      f@              L@       @     @e@      :@      2@      ,@      ,@     �R@      D@     �a@     @X@     @a@      2@     @U@      >@      *@      ]@       @     @b@             �G@      �?     �a@      6@      2@      @      $@      M@      9@     �]@     �T@     �[@      ,@      Q@      7@      (@     @U@      �?     �W@              <@             �\@      1@      (@       @      "@      I@      3@      Y@      O@     �S@      ,@      1@      @      �?      ?@      �?     �I@              3@      �?      ;@      @      @      @      �?       @      @      3@      5@      @@              6@      *@      @      9@      "@      ?@              "@      �?      <@      @              "@      @      1@      .@      7@      ,@      ;@      @      �?       @      �?       @      @       @               @              ,@                      @              @      &@      "@      @      (@      @      5@      &@       @      1@      @      7@              @      �?      ,@      @              @      @      $@      @      ,@      &@      .@      �?     @V@      4@      4@     �W@      @     �c@             �B@      @     `a@      8@      $@      @       @      O@      @     �P@     �Q@     �d@      *@       @                      0@              9@                      @      9@                                      @              "@      &@     �B@       @      @                      &@              ,@                               @                                       @              @      @      9@              @                      @              &@                      @      1@                                      �?               @       @      (@       @     @T@      4@      4@     �S@      @     ``@             �B@             �\@      8@      $@      @       @     �M@      @      M@      N@     �_@      &@      <@      "@      @      ?@       @     �S@              <@             �O@      �?      �?      @      �?      1@      @      9@      ;@     �P@      @     �J@      &@      .@      H@       @     �J@              "@             �I@      7@      "@      @      @      E@       @     �@@     �@@     �N@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�
hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @CK�;�@�	           ��@       	                    �?>BG�@�           j�@                          �:@!mS*�@�           ��@                           @1ڀHE�@�           (�@������������������������       �����@.           ��@������������������������       �8��
@n            �e@                          �?@�����@a            �b@������������������������       ������X@P            �^@������������������������       ����#
@             <@
                           �?�b:G5@�           T�@                           �?�d��@�           X�@������������������������       �����k@t             h@������������������������       ��P�@@!           �|@                            �?F��%j@F           P�@������������������������       ���`�_g@�           `�@������������������������       �X�m	�_@�            �q@                           @��QVr@�           P�@                           �?������@           ��@                           @��1��@�           8�@������������������������       ��Ӌ���@�            �s@������������������������       ���#�}�@           �z@                           @Fyd�!�@V             a@������������������������       ��h��@D            @\@������������������������       ��@w�B	@             8@                           @c'%8��@�            @r@                          �1@9�P?�@M            �_@������������������������       �3�U�nu@             =@������������������������       ��$��N>@<            �X@                           @�禒�
@`            �d@������������������������       ���Ip@6            �V@������������������������       ���g��@*            �R@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       Pv@     �_@     �T@     v@     �G@     @|@      @     `m@      B@     @|@     @V@      M@      B@     �Q@      p@     �O@      w@     Ps@     �{@     @Q@     �m@      V@     �G@     @q@      1@     �t@      @     �a@      :@     �t@      K@      D@      8@     �B@     �e@      F@     �p@      i@     �u@     �G@      W@      4@      4@     @^@      &@     �a@      @     �N@      (@     �b@      <@      (@      (@      "@     �S@      $@      ]@     @Z@     `d@      4@      T@      4@      *@     @\@      @     `a@       @      K@      @     ``@      ,@      (@       @       @     @R@      @      Y@     @W@      b@      2@     �Q@      ,@      *@     �X@      @     @\@       @     �F@      @     �W@      "@      (@      @      @      P@      @     @T@      S@      `@      2@      "@      @              ,@      �?      :@              "@             �B@      @              @      �?      "@              3@      1@      0@              (@              @       @      @       @      �?      @       @      3@      ,@              @      �?      @      @      0@      (@      3@       @      @              @       @      @       @      �?      @       @      0@      &@              @              @       @      0@      $@      2@              @               @                                      @              @      @                      �?      �?      @               @      �?       @      b@      Q@      ;@     `c@      @      h@      �?      T@      ,@      g@      :@      <@      (@      <@      X@      A@     �b@     �W@     �g@      ;@      K@      C@      (@      T@      @      I@      �?     �A@      $@      Q@       @      &@       @      (@     �F@      4@      J@     �E@     �S@      3@      8@       @      @      @@      �?      1@              "@              0@       @       @      @      @      3@              0@      *@      2@      �?      >@      >@      "@      H@      @     �@@      �?      :@      $@      J@      @      "@       @      @      :@      4@      B@      >@     �N@      2@     �V@      >@      .@     �R@             �a@             �F@      @      ]@      2@      1@      @      0@     �I@      ,@     �X@      J@     @[@       @     �P@      7@      @     �G@             @V@              @@      @     �Q@      1@      *@      @      *@      <@      *@     �M@      E@     @V@      @      8@      @      "@      <@              K@              *@      �?      G@      �?      @      �?      @      7@      �?      D@      $@      4@      �?     @^@     �C@     �A@     @S@      >@     �]@       @     �W@      $@     �]@     �A@      2@      (@      A@     �T@      3@     @Y@     @[@      X@      6@     �U@      @@     �A@     �J@      9@     �S@       @      S@      $@     �Q@      =@      ,@      &@      >@      K@      3@      T@     @U@      R@      0@     @R@      5@      =@     �E@      9@      O@       @     �P@      "@      L@      :@      *@      "@      =@     �H@      &@     @Q@     @R@     @P@      *@      6@       @      *@      5@       @      :@      �?     �@@      @      2@      &@      @       @      .@      :@       @      =@      C@      8@      @     �I@      *@      0@      6@      7@      B@      �?     �@@      @      C@      .@      @      @      ,@      7@      @      D@     �A@     �D@       @      ,@      &@      @      $@              1@              $@      �?      .@      @      �?       @      �?      @       @      &@      (@      @      @      &@      @      @      "@              0@               @      �?      &@      @      �?              �?      @      @      $@      (@      @      @      @      @      @      �?              �?               @              @                       @                      @      �?                              A@      @              8@      @     �C@              2@             �G@      @      @      �?      @      <@              5@      8@      8@      @      *@      @              @      @      3@              $@              ,@      @                      @      (@               @      @      .@      @                              @       @      $@              @              @                              @       @                                      �?      *@      @              @      @      "@              @              &@      @                              $@               @      @      .@      @      5@      �?              1@              4@               @             �@@      �?      @      �?      �?      0@              *@      2@      "@       @      (@                      @              0@              @              7@      �?                              @               @      "@      @      �?      "@      �?              &@              @               @              $@              @      �?      �?      (@              @      "@      @      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ���4hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�bSf�@�	           ��@       	                   �?@t�@�&�@           ��@                           �?ܶ�;]@�           ؘ@                            @=ْm�@U           P�@������������������������       �{`�S<\@�            Px@������������������������       �:��Jv@`            �d@                          �:@|Eg�5�@�           0�@������������������������       �5�v�$�@           x�@������������������������       � �?!�t@v            �g@
                           �?���=@E            @\@                           �?�ׯ���	@             B@������������������������       �p�y	O�@             4@������������������������       �+�%W�@
             0@                            �?�VR��@/            @S@������������������������       �ˣS���@             @@������������������������       ���Mc�
@            �F@                          �3@lS��<@�           D�@                            �?P��#/@H           (�@                           @��9�W
@T           Ȁ@������������������������       ���50�	@�            q@������������������������       �zX2��	@�            �p@                           �?zl6Ӕ*@�            �v@������������������������       �uߣ%S�	@{            �f@������������������������       �6��De�
@y             g@                           @T�G�6@A           t�@                           @���t@�           �@������������������������       �\�7?U@�           ��@������������������������       ����!�@k            �e@                          �8@L?�� @C           �@������������������������       �	�9 �@�            u@������������������������       �E�|��@l             e@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@     �]@     �U@     �u@     �@@     }@      @     �l@     �C@     �}@      W@     �M@      F@      N@     �k@      Q@     �w@     �s@     �{@     �T@      b@     �M@     �N@     �b@      :@     �a@      @     @\@      :@     @d@     �D@      @@      <@     �F@     @W@     �A@     �b@     �b@     �h@     �E@     �a@      D@     �G@     @b@      8@     `a@      @     @Z@      :@     �c@      C@      ?@      1@      D@     �V@      =@     @b@      a@      h@      D@     �K@       @      4@     �L@      @      N@              <@       @     �K@      *@      @      @      @     �@@      (@     �A@     �I@     @W@      *@      E@      @      "@     �E@             �G@              1@             �D@       @      @      @      @      :@      (@      8@      9@     �O@      &@      *@       @      &@      ,@      @      *@              &@       @      ,@      @      �?                      @              &@      :@      >@       @     @U@      @@      ;@     @V@      5@     �S@      @     @S@      8@      Z@      9@      8@      *@     �A@      M@      1@     �[@     �U@     �X@      ;@     �R@      8@      8@     �N@      4@      S@       @      K@      4@     �X@      4@      6@      @      >@     �G@      $@      W@     �P@     �R@      9@      &@       @      @      <@      �?      @      �?      7@      @      @      @       @      @      @      &@      @      3@      3@      8@       @      @      3@      ,@      @       @      @               @              @      @      �?      &@      @       @      @      @      ,@      @      @      �?      @      "@      �?       @      �?                              �?      @      �?              @      �?       @              @                      �?       @       @      �?              �?                              �?              �?               @      �?       @                                              @      �?               @                                              @                      �?                              @                      @      *@      @      @               @               @               @                      &@       @      �?      @      @      "@      @      @       @       @                               @              @                                      @                      @              @       @       @       @      &@      @      @                              �?               @                      @       @      �?              @      @      @      �?     �h@      N@      :@     `h@      @     0t@      �?     �\@      *@     �s@     �I@      ;@      0@      .@      `@     �@@      m@     �d@      o@      D@     �K@      2@      @     �T@      �?     �c@             �O@      �?     �d@      "@      @       @      @      I@      (@     �X@     �G@      ^@      @      @@      (@      @      G@             �R@             �@@      �?     �]@      @      �?       @             �B@      @     �M@      8@     @T@      @      $@      @      @      =@              <@              @             �P@      @      �?                      8@      @     �B@      $@     �E@       @      6@      @              1@              G@              :@      �?     �J@                       @              *@      �?      6@      ,@      C@      @      7@      @       @      B@      �?     �T@              >@              G@      @      @              @      *@      @      D@      7@     �C@      �?       @      @              >@      �?      C@              1@              ,@              �?              �?      @       @      0@      (@      ?@      �?      .@      @       @      @             �F@              *@              @@      @      @               @       @      @      8@      &@       @              b@      E@      5@     @\@      @     �d@      �?      J@      (@     �b@      E@      5@      ,@      (@     �S@      5@     �`@     �]@      `@      A@     @S@      :@      $@     �S@      @      Z@              F@      @     �Y@      ;@      0@      (@      @     �A@      4@     �Q@     @R@      P@      ;@      Q@      9@       @      P@      @     �S@              =@      @     �U@      5@      *@      $@      @      =@      *@     �I@     �L@      F@      6@      "@      �?       @      ,@              :@              .@       @      .@      @      @       @      @      @      @      4@      0@      4@      @     �P@      0@      &@     �A@       @      O@      �?       @      @     �G@      .@      @       @      @      F@      �?     �O@     �F@      P@      @     �C@      "@      @      :@             �G@              @      @     �A@      $@       @       @      @      =@      �?      H@      @@      >@      @      <@      @      @      "@       @      .@      �?      �?              (@      @      @                      .@              .@      *@      A@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�HqhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��4d�@�	           ��@       	                    �?��AK#@:           �@                          �9@%�A��@�           ؃@                            @e��E��@V           Ѐ@������������������������       �-利�@           0y@������������������������       �XB���;@P            �`@                            �?�ؑț�@@            @X@������������������������       ����՗@)            �P@������������������������       �O����o@             ?@
                            @R��^+ @�           ��@                           @�"�(a�@+           �@������������������������       �Mѣ��w@�            �p@������������������������       ���mp�%
@�            �n@                          �:@7�.�S@y            �g@������������������������       �j�i�@i            @c@������������������������       ����qOY@            �A@                            @6H|��@^            �@                          �5@J-�:�q@y           �@                            �?إ�[��@^           p�@������������������������       �7�p� �@�           H�@������������������������       ��m3�@�            �l@                           @6�g���@           ��@������������������������       ��VY�"T@�            �t@������������������������       ��2�ܩ@F           8�@                           @��Xut@�           `�@                          �;@�H���@n           �@������������������������       ���A#��@/           �{@������������������������       �F!�{@?            �X@                           @��B�@w            @e@������������������������       �Y �Ym�
@K            @[@������������������������       �\��o@,            �N@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       @u@     �b@     �X@     �v@     �B@     }@      @     �j@      <@     �y@     �\@     �N@      B@     @P@     �o@     @Q@     `x@      s@     �z@     @R@     �Z@     �@@     �B@     �^@       @     @d@      �?     @U@      @     @d@     �J@      0@       @      2@      X@      .@      _@     �S@     `e@      A@      K@      0@      3@     �E@      @     �T@      �?     �C@      �?     �U@      7@      $@      @      @     �G@      @     �E@     �E@     �U@      4@      I@      *@      ,@     �A@      @     �S@             �B@             �Q@      4@      @      �?      @     �B@              D@     �B@     @S@      ,@      A@      *@      @      ;@       @      N@              6@              L@      *@      @               @      :@             �A@      <@     �P@      &@      0@              $@       @      @      2@              .@              .@      @              �?      @      &@              @      "@      $@      @      @      @      @       @      �?      @      �?       @      �?      .@      @      @       @       @      $@      @      @      @      $@      @      @      �?      @      @              @              �?              ,@       @      @      �?       @       @       @       @      @       @      @               @               @      �?      �?      �?      �?      �?      �?      �?      @      �?               @      �?      �?      �?       @      @     �J@      1@      2@     �S@      �?     �S@              G@      @      S@      >@      @      @      &@     �H@      (@     @T@      B@      U@      ,@      B@      $@      (@     �K@             @Q@              >@       @     �M@      .@      @      @      @     �B@      �?     �P@      >@     �Q@      @      3@      $@      @     �@@              7@              ,@      �?      >@      .@      �?      @      @      8@              >@      .@      @@      @      1@              "@      6@              G@              0@      �?      =@               @              �?      *@      �?     �B@      .@      C@              1@      @      @      8@      �?      $@              0@      @      1@      .@      @              @      (@      &@      ,@      @      ,@      "@      1@      @      @      (@      �?      $@              ,@      @      1@      (@      �?              @      @      @      ,@      @      (@      "@                              (@                               @                      @       @              �?      @      @              @       @              m@     �\@      O@     `n@      =@     �r@       @     �_@      6@     �o@      O@     �F@      <@     �G@     �c@      K@     �p@     `l@     @p@     �C@     @e@     @T@      A@     �g@      (@     @m@      �?     @S@      (@     `f@     �E@      B@      5@      ?@     �_@      A@     �h@     �c@      h@      @@      Q@      >@      4@     �Z@             @a@              B@      @     @Y@      5@      7@      .@      "@     �O@      ,@     @\@     @Z@      ^@      3@     �H@      9@      3@     �T@             �X@              5@      @     �R@      .@      1@      .@      @     �E@      ,@      V@     �W@     @W@      1@      3@      @      �?      8@              D@              .@              :@      @      @               @      4@              9@      &@      ;@       @     �Y@     �I@      ,@     @T@      (@      X@      �?     �D@       @     �S@      6@      *@      @      6@     �O@      4@      U@      K@     @R@      *@     �F@      2@      @      8@      @     �J@      �?      3@       @      D@      .@      "@      @      @      6@      @      ;@      $@      6@      @     �L@     �@@      "@     �L@      "@     �E@              6@      @      C@      @      @       @      .@     �D@      .@     �L@      F@     �I@      "@     �O@      A@      <@     �K@      1@     @Q@      �?      I@      $@     �R@      3@      "@      @      0@     �@@      4@     @Q@      Q@     �P@      @      J@      ;@      9@     �@@      1@      K@      �?      C@      $@     �D@      ,@       @      @      .@      9@      1@      L@     �J@     �H@      @      G@      1@      4@      :@      *@     �J@      �?      =@      "@      ?@      *@       @       @      &@      4@      .@     �K@     �B@      B@      @      @      $@      @      @      @      �?              "@      �?      $@      �?              @      @      @       @      �?      0@      *@              &@      @      @      6@              .@              (@             �@@      @      �?      �?      �?       @      @      *@      .@      2@       @      @       @       @      (@              (@              "@              7@      @                               @      @      $@      &@      *@              @      @      �?      $@              @              @              $@              �?      �?      �?      @              @      @      @       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�n�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �3@������@�	           ��@       	                     @�:��Q	@y           ��@                           @�	0�P@�           ��@                           �?9m���@�            �x@������������������������       �Fѝ�C�@�            �p@������������������������       ����T�	@P             `@                           @(��!"6@�           X�@������������������������       ��Ц]��
@�            �s@������������������������       ���,�z�
@�            �r@
                          �1@�<G@�            w@                           @N(b�1�@l            �c@������������������������       �(Ɓ1�^@G             Z@������������������������       �u�����
@%            �K@                           @b+_�u�@�            @j@������������������������       ��8���@x            �f@������������������������       �$މ�q@             =@                           �?nɎJ�(@6           ȣ@                           @;:�q@�           �@                            @L/�@�           ��@������������������������       ��B��a)@�           ؅@������������������������       ����G}N@0           �~@������������������������       �|�K-�@             5@                           @3�jN�@7           ��@                          �5@b� ��@Y           ��@������������������������       �JT^/�Y@�            �u@������������������������       �K%q]�E@}           ��@                           �?Z�,��@�            pw@������������������������       ��Z�v�@j            `e@������������������������       �k�L:eG@t            �i@�t�bh�h5h8K ��h:��R�(KKKK��h��B        �v@     `b@      S@     Pt@      B@     P{@      @      q@      5@     P|@     �Y@     �L@      @@     �P@     �l@      R@     x@     �r@     �{@     �V@     @W@      ?@      6@     �_@       @      i@      �?      X@      @     �h@      =@      6@      @      @     @T@      7@     @_@     �V@     @h@      9@      L@      6@      &@     @Y@      @     @b@              O@      @     �c@      .@      3@      @      @      L@      &@     @Y@     �P@     �c@      1@      3@      @      @     �L@       @     �A@              8@      @      G@      (@      @              @      :@      @     �C@      ?@      O@      "@      0@      @      @     �@@       @      8@              .@      @      :@       @      @               @      4@      @      .@      8@     �G@      @      @              �?      8@              &@              "@              4@      @                       @      @              8@      @      .@      @     �B@      .@      @      F@      �?     �[@              C@      �?     �[@      @      (@      @              >@      @      O@     �A@     @X@       @      (@       @      @      <@             �N@              ,@             �J@      �?      (@      �?              2@      @     �B@      "@      J@      @      9@      @       @      0@      �?      I@              8@      �?     �L@       @               @              (@      �?      9@      :@     �F@      @     �B@      "@      &@      :@      @      K@      �?      A@             �E@      ,@      @      �?       @      9@      (@      8@      9@     �A@       @      0@      @       @      &@       @      8@      �?      (@              >@      @      @               @      "@      @      @      @      @      @      &@      @      @      @              $@      �?       @              6@      @       @                      @      @      @       @      @      @      @              @      @       @      ,@              @               @              �?               @      @               @      @      �?              5@       @      @      .@      @      >@              6@              *@       @              �?              0@      @      3@      3@      <@      @      2@       @      @      $@      @      >@              .@              &@       @              �?              .@      @      3@      0@      4@      @      @                      @                              @               @                                      �?                      @       @             �p@      ]@      K@     �h@      <@     �m@      @      f@      1@     �o@     �R@     �A@      <@      N@     `b@     �H@     @p@     �j@      o@     @P@     �X@     �Q@      C@     �X@      3@      U@      @     @Z@      .@     �[@     �A@      7@      1@     �E@     �Q@      =@     �]@      V@     �Z@     �B@     �X@     �O@      C@     @X@      .@      U@      @     �Y@      .@     �[@     �@@      7@      1@     �E@      Q@      =@     �\@      V@     �Z@     �B@      G@      C@      3@     �P@      @      K@       @     �N@      @     @U@      2@      @      &@      0@      F@      4@     @R@     �B@      R@      6@      J@      9@      3@      >@      &@      >@      @      E@      &@      :@      .@      1@      @      ;@      8@      "@      E@     �I@      A@      .@              @              �?      @                       @                       @                               @              @                             `e@      G@      0@      Y@      "@      c@             �Q@       @     �a@     �C@      (@      &@      1@     @S@      4@     �a@      _@     �a@      <@     �^@      8@       @      S@       @     �^@              P@       @     �X@      5@      $@      "@      @     �L@      1@     �X@     �W@     @U@      8@     �@@       @      @      >@      @      G@              3@             �B@      @      @       @       @      .@      @     �D@     �J@      :@      "@     @V@      0@      @      G@      @     @S@             �F@       @      O@      .@      @      �?      @      E@      (@     �L@     �D@     �M@      .@     �H@      6@       @      8@      �?      >@              @              F@      2@       @       @      $@      4@      @      F@      >@     �L@      @      5@      &@      @      "@      �?      2@              @              8@      $@               @      �?       @       @      *@      .@      9@       @      <@      &@      @      .@              (@              �?              4@       @       @              "@      (@      �?      ?@      .@      @@       @�t�bub�s     hhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�9RhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���Y�@z	           ��@       	                     @`���@7           p�@                          �:@+��M@`           ؍@                           �?�xU@            �@������������������������       �W�E8v>@&           �|@������������������������       � #PCP@�            @w@                          �=@���[6@N            �^@������������������������       �:�R@1            �U@������������������������       �.���ʸ
@            �B@
                           �?�ҩ�m@�            v@                           �?�j�@�!@            �K@������������������������       �(���	@             7@������������������������       �ˣS��N@             @@                           �?"tVͅ�@�            �r@������������������������       �v9�)@R            �a@������������������������       �Nh��r@f            �c@                           @��	�O@C           Z�@                          �4@]��I�@�           �@                            �?ʊ�-@T           (�@������������������������       �8��C�@�             s@������������������������       �Y��I�@�            �n@                           �?^k��o@Z           ��@������������������������       �#�M�@�             m@������������������������       �'A���	@�           X�@                          �4@�����@�           А@                           @i,� ��@E           ؀@������������������������       ���S�	@�            �p@������������������������       �Rksv@�             q@                            �?e�\@P           Ȁ@������������������������       ����!��@U             a@������������������������       �I�4:Q@�            y@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �a@     �Y@     �v@     �K@     `}@       @     �h@     �@@     �|@     �[@     @Q@      G@     @Q@     @k@      Q@      u@     �t@     @{@     �U@     �\@     �B@      ?@      [@      "@      h@       @      T@      $@     �d@      A@      .@      @      8@     �T@      @     @]@     �W@     @b@      @@     �Q@      8@      6@     @U@      @     �c@             �E@      �?     �`@      9@      &@      @      *@     �O@      @     �T@     @S@     @\@      3@      O@      3@      2@      T@      @      b@             �C@      �?     @^@      1@      @              $@      K@             �Q@     �O@     @[@      *@      <@      *@      $@      @@              U@              5@             @T@      @      @              @      ?@              6@      C@     �R@      $@      A@      @       @      H@      @     �N@              2@      �?      D@      $@      @              @      7@              H@      9@     �A@      @       @      @      @      @              *@              @              *@       @      @      @      @      "@      @      *@      ,@      @      @       @      �?              @              @              @              @       @      @      @      �?      @       @      "@      *@      @      @              @      @      �?              @                              @              �?      �?       @      @      �?      @      �?      �?             �F@      *@      "@      7@      @      A@       @     �B@      "@      >@      "@      @              &@      4@      @      A@      2@     �@@      *@       @      @      �?      @              @       @      &@      @       @       @                              �?                      @      @              �?       @      �?       @               @       @      @                       @                              �?                       @       @              @      @              @               @              @      @       @                                                               @      @             �B@       @       @      1@      @      >@              :@      @      <@      @      @              &@      3@      @      A@      ,@      ;@      *@      1@      @      @       @      @      (@              .@      @      ,@       @       @              �?      &@              *@      @      ,@      &@      4@      @      @      "@      �?      2@              &@       @      ,@      @       @              $@       @      @      5@      "@      *@       @      i@     �Y@     �Q@     �o@      G@     `q@      @     �]@      7@     @r@     @S@      K@     �C@     �F@     �`@     �N@     `k@     �m@      r@      K@     @]@     �Q@     �M@     @c@     �B@     @^@      @     �R@      *@     �b@     �H@     �B@      4@     �A@     @T@     �D@     �a@      a@     �b@     �D@      D@      1@      .@     @P@      ,@     �H@      �?      0@      �?      F@      5@      $@      @      @      <@      0@     �K@     �E@     �R@      ;@      .@      @      &@      I@              =@              "@      �?      8@       @      @      @      @      ,@      $@      4@      :@     �F@      5@      9@      &@      @      .@      ,@      4@      �?      @              4@      *@      @              @      ,@      @     �A@      1@      >@      @     @S@     �J@      F@     @V@      7@      R@       @     �M@      (@     �Z@      <@      ;@      .@      <@     �J@      9@     @U@     @W@     �R@      ,@      &@      (@      3@      1@              7@       @       @      @      ?@      @      @               @      *@      $@      3@      :@      3@      �?     �P@     �D@      9@      R@      7@     �H@             �I@      "@      S@      6@      6@      .@      4@      D@      .@     �P@     �P@     �K@      *@     �T@     �@@      (@     @Y@      "@     �c@      @      F@      $@     �a@      <@      1@      3@      $@      K@      4@     �S@     �Y@     �a@      *@      >@      "@      @      F@              W@              2@      @      T@       @      $@      "@              6@      "@     �D@     �L@     @W@      $@      (@       @      �?      ;@             �B@              @             �M@              @      @              *@       @      5@      7@      H@      @      2@      @      @      1@             �K@              *@      @      5@       @      @       @              "@      @      4@      A@     �F@      @     �J@      8@       @     �L@      "@     @P@      @      :@      @     �N@      4@      @      $@      $@      @@      &@      C@     �F@      H@      @      &@       @      @      ;@              6@              @              *@      @              �?      @      @      @      @      .@      (@              E@      0@      @      >@      "@     �E@      @      7@      @      H@      ,@      @      "@      @      =@       @      A@      >@      B@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ{�/hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�S�@�	           ��@       	                    �?�n�I��@           *�@                          �4@a��XP @%           P�@                           �?u��~��@|            �@������������������������       ���ɉ�-@�             o@������������������������       �h"\!��@�            pv@                           �?ICͶ{@�            �p@������������������������       ��_�6O@7             X@������������������������       ��cO@r            @e@
                           @���F.�@�           ��@                          �1@��u�=@{           ȏ@������������������������       ���#!c�
@�            �s@������������������������       �5.�Ę@�           ��@                           @`Ꮏ@g           ��@������������������������       �He����@#           0|@������������������������       ��`���
@D            �[@                            @��
"�@�           Ж@                           @nP߈��@b           �@                           �?e֕�H@�           `�@������������������������       ������@�            �q@������������������������       ��H�-.@            }@                          �;@�.݊�@�            �n@������������������������       ��}�u@s             f@������������������������       ��}��@)             Q@                           @bLʕ��@'           0}@                           �?K��n@           �y@������������������������       �%��^Ai@�             r@������������������������       ������%@I             ^@                           �?��G���@%            �M@������������������������       ���x[
@             7@������������������������       ��HSvݤ@             B@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �v@     @_@     @U@      t@      D@     �}@      @     �m@      =@      z@     �Z@     �Q@      =@      L@     @n@      R@     w@      s@     @~@     �T@     �i@     �P@     �F@     �i@      ;@     �v@             �`@      &@     �q@      N@     �D@      $@      @@      b@      >@     �m@      h@     @t@     �G@     @V@      =@      9@     @R@      2@     @Y@              I@      "@     �R@      7@      4@              :@     �J@      .@     �R@      Q@     �Y@      6@     �P@      *@      .@     �G@      0@     @Q@              :@      @      F@      4@      *@              *@     �F@      (@     �J@     �H@     �T@      1@      >@      @      @      ,@      @      =@              @       @      2@       @      @              @      "@      "@      7@      5@     �D@      *@      B@      @       @     �@@      *@      D@              4@      @      :@      (@       @              "@      B@      @      >@      <@      E@      @      7@      0@      $@      :@       @      @@              8@       @      ?@      @      @              *@       @      @      6@      3@      4@      @      $@      @       @      &@       @      ,@              2@              @      �?      �?              &@                       @       @       @      �?      *@      *@       @      .@              2@              @       @      ;@       @      @               @       @      @      ,@      1@      (@      @     @]@      C@      4@     ``@      "@     @p@             �T@       @     �i@     �B@      5@      $@      @     �V@      .@     `d@     @_@     �k@      9@     �S@      7@      0@     @W@      @      c@             �K@             �c@      <@      @      @      �?      N@      @      X@     �Q@     �a@      3@      (@      @      @      7@      @      N@              7@             �K@       @      �?              �?      0@      �?      :@      7@     �K@      @     �P@      3@      *@     �Q@       @     @W@              @@             �Y@      :@      @      @              F@       @     �Q@      H@      V@      *@      C@      .@      @      C@      @     �Z@              <@       @      H@      "@      ,@      @      @      ?@      (@     �P@      K@     �S@      @      @@      .@      @      B@       @      U@              6@       @     �A@      @      &@      �?      @      5@      "@      K@      C@     �P@      @      @                       @      �?      7@              @              *@       @      @       @              $@      @      *@      0@      &@             �c@      M@      D@     �]@      *@     @\@      @      Z@      2@      a@     �G@      =@      3@      8@     �X@      E@     ``@     @\@      d@     �A@     �[@      E@      4@     @U@      &@     @V@      @      P@      @     �X@      <@      1@      ,@      $@      S@      @@      W@     �M@     �]@      1@     @Q@     �A@      *@     �P@      &@      P@      @     �M@      @      T@      7@      ,@      &@      @     �L@      =@      Q@     �F@      S@      0@      B@      @      @      2@      @      >@      �?      <@      @      :@       @      �?      @       @      9@      @      :@      6@      8@      @     �@@      @@      @      H@      @      A@       @      ?@              K@      .@      *@      @      @      @@      7@      E@      7@      J@      "@     �D@      @      @      3@              9@       @      @              3@      @      @      @      @      3@      @      8@      ,@     �E@      �?      @@      @      �?      1@              3@              @              &@      @      @       @      @      3@      @      1@      *@      6@      �?      "@       @      @       @              @       @                       @       @              �?      �?                      @      �?      5@              G@      0@      4@     �@@       @      8@      �?      D@      ,@     �B@      3@      (@      @      ,@      6@      $@     �C@      K@     �D@      2@     �B@      $@      1@      ?@              8@      �?     �C@      &@      A@      1@      $@      @      &@      .@      @     �A@      I@      C@      2@      7@      @      0@      5@              5@      �?      <@      &@      ,@       @      @      @       @      ,@      @      :@     �A@      ?@      (@      ,@      @      �?      $@              @              &@              4@      "@      @      �?      @      �?      �?      "@      .@      @      @      "@      @      @       @       @                      �?      @      @       @       @      �?      @      @      @      @      @      @              @       @      �?      �?                                      @      @       @                      �?       @      @                      �?              @      @       @      �?       @                      �?                               @      �?       @      @      �?      @      @       @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ4�-hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�D)N:�@�	           ��@       	                    @AfL�@�           ��@                           �? ��Z�y@�           `�@                          �4@Tѝވ @c           ��@������������������������       �/��&N@           Py@������������������������       �Ǘ���@[            @a@                          �3@��rI�@K           ȍ@������������������������       �."4@1           �}@������������������������       �*��)�)@            ~@
                          �5@\{����@K           8�@                           �?�t8 F�@           ��@������������������������       ����r�{
@           `{@������������������������       �����N@�            �w@                           �?FE��
@6            �T@������������������������       �f��i	@             J@������������������������       ���R�@             ?@                           @�m��إ@�           ��@                          �@@btvR@|           8�@                           @�m�t@\           ؎@������������������������       �ӹ��J�@�           ��@������������������������       �[�d��*@�            �r@                           �?��*_@             �I@������������������������       � ���$�@
             7@������������������������       ��W.��@             <@                           �?Vz�1�q@(           �}@                           @Κ��R�
@_            `b@������������������������       ����-�7@             B@������������������������       �ޖ4*�	@L            �[@                          �:@���?�@�            �t@������������������������       ����z��@�            �k@������������������������       �	C�u�@>            �Z@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       0u@      a@     @V@     �u@      C@     �}@       @     �m@      7@     �{@     �Z@      M@     �E@     �O@     �k@     �M@     �w@     �t@     �z@     �V@      g@     @Q@     �F@      l@      .@     Pv@      @     �a@       @     pq@     �I@     �D@      *@      =@     ``@      >@     @m@     @h@     pr@     �J@     �\@      H@     �@@     �b@      ,@     �f@      @     @U@      @     `e@      A@      ;@      @      ;@     @U@      <@     �c@     �`@      c@      F@     �G@      4@      (@      H@      @      U@       @      <@             @Q@      @      "@      �?      @      A@      �?     �M@      H@      J@      ,@      =@      *@       @      D@       @     �Q@              .@              O@      @      @      �?       @      ;@      �?      B@     �B@     �C@      (@      2@      @      @       @      �?      *@       @      *@              @       @       @              @      @              7@      &@      *@       @      Q@      <@      5@      Y@      &@      X@      �?     �L@      @     �Y@      =@      2@      @      4@     �I@      ;@     �X@     @U@      Y@      >@      ;@      .@      *@     �J@      @     �F@      �?      =@       @     �G@      3@      @      �?      @      2@      ,@     �L@      C@      Q@      $@     �D@      *@       @     �G@      @     �I@              <@      @     �K@      $@      &@      @      .@     �@@      *@      E@     �G@      @@      4@     �Q@      5@      (@     @S@      �?      f@             �L@       @      [@      1@      ,@       @       @      G@       @      S@     �N@     �a@      "@     @P@      0@       @     �P@      �?     �c@              J@      �?     @X@      *@      ,@       @       @     �E@       @     �Q@      N@     @a@       @      C@      "@      @      B@      �?     �V@              2@              I@      @      �?      @       @      9@              B@      8@     @V@      @      ;@      @      @      >@             @P@              A@      �?     �G@       @      *@      @              2@       @      A@      B@     �H@      @      @      @      @      &@              5@              @      �?      &@      @                              @              @      �?      @      �?      @      @      @      @              (@              @      �?      $@      @                              @              @                                       @      �?       @              "@               @              �?                                                      �?      �?      @      �?     @c@     �P@      F@     @^@      7@      ]@      @     �W@      .@      d@     �K@      1@      >@      A@     �V@      =@     �b@      a@     �`@      C@      V@      G@     �B@      T@      5@     @R@      @     �U@      *@     �Z@     �B@      0@      9@      ;@     @R@      6@     �W@     �U@      T@      7@     @T@     �A@     �A@     @S@      5@     @R@      @     @T@      *@      Z@      @@      ,@      4@      8@     �Q@      5@     �W@      U@      T@      7@      N@      5@      >@      M@      @     �L@      @      O@      $@      P@      >@      *@      .@      (@      H@      $@     �P@      O@      F@      .@      5@      ,@      @      3@      .@      0@              3@      @      D@       @      �?      @      (@      7@      &@      ;@      6@      B@       @      @      &@       @      @                              @               @      @       @      @      @       @      �?              @                      @      @               @                              @                      @               @               @      �?                                      @      @       @      �?                              �?               @               @      @      @                              @                     �P@      5@      @     �D@       @     �E@      �?       @       @     �K@      2@      �?      @      @      1@      @     �K@      I@     �K@      .@      3@      �?      @      (@      �?      0@               @              7@       @                              @              2@      4@      3@      @      @              �?      �?      �?      @               @              @                                      @                      *@                      *@      �?      @      &@              *@                              1@       @                              @              2@      @      3@      @     �G@      4@      @      =@      �?      ;@      �?      @       @      @@      0@      �?      @      @      $@      @     �B@      >@      B@      (@      ?@      1@       @      6@              3@              @      �?      :@      @              �?      @      @      @      7@      0@      <@      (@      0@      @      �?      @      �?       @      �?       @      �?      @      (@      �?      @      �?      @       @      ,@      ,@       @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�q8rhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@�`V)2�@�	           ��@       	                    @��
�@           d�@                            @b�����@�           T�@                           �?"���@�           8�@������������������������       �V:�);@|            �h@������������������������       �)Wr���
@           �@                           �?�I���@�            �r@������������������������       �M��D��@b            @e@������������������������       �Pہ�m�@U            �`@
                            @�gqx/@�            @t@                          �1@;�Ż_j@�            �n@������������������������       �.`�Rl�	@S            �`@������������������������       �$�z�
@E            �\@                          �2@f����@5            @S@������������������������       �Qr�":@&            �J@������������������������       �P:&У@             8@                           �?v�.�@+           `�@                          �9@`��<@�           ��@                            @.��R��@�           8�@������������������������       ��j*�@           p{@������������������������       �YA ���@�             s@                          �@@a��7@	           `y@������������������������       �
��[3@�            �v@������������������������       ����
@            �F@                          �9@�k�2�@R           ̔@                           �?g>dY��@m           @�@������������������������       ���b�e@�             x@������������������������       �Ex8��x@�           @�@                           @h&�R@�            �v@������������������������       ����c,@�             q@������������������������       ��,TE@<            �V@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       @u@      a@     �X@     @u@     @P@     �~@       @      k@     �@@      z@     @]@     �L@     �C@     @S@     �k@     @Q@     w@     0q@      }@     @S@     �Z@      >@      ?@     �`@      *@     �m@       @      S@      �?     �d@      <@      8@      @      (@      U@      3@      `@      W@      m@      *@     �R@      3@      4@     �Y@      *@     �f@       @     �P@      �?     �`@      9@      7@      @      $@     �N@      ,@     �W@      Q@     �g@      @     �H@      .@      "@     �R@      @     �a@              G@      �?     @Z@      &@      4@      @      @      D@      @     �Q@      E@      c@      @      .@      @      @      3@      @      :@               @      �?      8@      @      &@              @      *@              @      1@      @@      �?      A@      (@      @      L@             �\@              C@             @T@      @      "@      @      @      ;@      @      P@      9@      ^@      @      :@      @      &@      ;@      @     �C@       @      4@              =@      ,@      @              @      5@      @      7@      :@     �C@       @      $@       @      @      *@      @      .@       @      "@              *@       @      @              @      4@      �?      2@      *@      =@              0@       @      @      ,@              8@              &@              0@      @                              �?      @      @      *@      $@       @      ?@      &@      &@      >@             �L@              $@             �@@      @      �?               @      7@      @      A@      8@      E@      @      4@      @      @      6@             �F@               @              ;@      @      �?               @      2@      @      ?@      0@      C@      @      0@      @      �?      ,@              4@              @              3@              �?              �?      (@              @      &@      8@              @       @       @       @              9@              @               @      @                      �?      @      @      9@      @      ,@      @      &@      @       @       @              (@               @              @                                      @       @      @       @      @      @      "@      @      @      @              @              �?              @                                               @       @      @      @      @       @              @      @              @              �?                                                      @              �?      �?                     @m@     �Z@      Q@      j@      J@     �o@      @     �a@      @@      o@     @V@     �@@      A@     @P@     @a@      I@      n@     �f@      m@      P@     �Y@     �N@      H@     �W@     �B@     �R@      @      U@      1@     �X@      B@      3@      1@      G@     �L@      9@     �Z@     �R@     �\@      ?@     @R@      ?@      :@      M@     �@@      K@       @     �C@      &@     �T@      4@      $@      @      ;@      @@      &@     @S@      H@     �R@      ;@      G@      3@      (@     �C@      .@      4@       @      5@      @      H@      @      @               @      :@       @      H@      :@      O@      3@      ;@      (@      ,@      3@      2@      A@              2@      @     �A@      ,@      @      @      3@      @      @      =@      6@      *@       @      >@      >@      6@      B@      @      4@      @     �F@      @      0@      0@      "@      &@      3@      9@      ,@      >@      :@     �C@      @      >@      6@      ,@      @@      @      3@      @      C@      @      ,@      *@      "@      "@      ,@      8@      *@      ;@      :@     �C@      @               @       @      @              �?              @               @      @               @      @      �?      �?      @                             ``@      G@      4@     �\@      .@     `f@             �L@      .@     �b@     �J@      ,@      1@      3@     @T@      9@     �`@     @[@     �]@     �@@     �X@      C@      $@      V@      @      a@              F@      *@      ^@     �B@      &@      $@      $@     �N@      *@     @W@     @V@     �R@      3@      G@      *@      @      A@              L@              4@             �G@      1@       @               @      ?@              B@     �@@     �@@       @      J@      9@      @      K@      @     @T@              8@      *@     @R@      4@      "@      $@       @      >@      *@     �L@      L@     �D@      &@     �@@       @      $@      :@      (@      E@              *@       @      >@      0@      @      @      "@      4@      (@     �D@      4@     �F@      ,@      .@      @      @      .@      &@     �C@              @       @      8@      .@      @      @       @      3@      "@      ?@      $@     �A@      $@      2@      �?      @      &@      �?      @              @              @      �?                      �?      �?      @      $@      $@      $@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ<l\hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�L�|@�	           ��@       	                    �?�1`���@�            �@                            @{���U�@:           �@                          �6@���^@�             t@������������������������       �vCA�1@r             h@������������������������       �q4���_@R             `@                           �?��C]�@v             h@������������������������       ��q���
@!            �I@������������������������       �����g@U            �a@
                           @A��*�@�           �@                          �?@����@4           �~@������������������������       �U��g��@            �|@������������������������       � F�k�@            �@@                            �?2PE� a@�           ؂@������������������������       �~��$�@r            �e@������������������������       �_R��&@           �z@                          �3@]�0,@�           �@                            @�W�!@f           ��@                           @�Fb��
@�           ��@������������������������       ��nu�c�	@            �@������������������������       �����,�@l            �f@                           @s��4Ý@{            �g@������������������������       ���s9@N            @^@������������������������       ���2qZ�@-             Q@                           �?��^�@?           ��@                          �5@��K%4�@�           ��@������������������������       �z}J��@�            �i@������������������������       �.��U@           �z@                          �=@��[�@�           ��@������������������������       ��j.r�@�           �@������������������������       �{�Y�r�@!            �J@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     `b@     �U@     @w@      <@     p@       @      i@      A@     �{@      ]@     �L@      ;@     �S@     �k@      N@     0v@     t@     @}@     @R@     �Z@     @S@      P@      e@      7@      a@       @     @Z@      3@     �`@     �L@      ;@      *@      J@     @X@      ?@      a@      b@      f@      A@      8@      $@      6@      H@      @     �F@      �?     �E@      @      L@      ,@      @      @      .@     �B@      @      I@     �D@     @P@      .@      2@      $@      &@      ;@       @      @@              7@      �?      D@      @      @      @      @      6@      �?      @@      7@      G@      (@      .@      @      @      2@       @      4@              2@      �?      5@      @      �?              @      @              0@      1@      ?@      @      @      @      @      "@              (@              @              3@      @      @      @              .@      �?      0@      @      .@      @      @              &@      5@      �?      *@      �?      4@      @      0@      @      @              $@      .@      @      2@      2@      3@      @      @              �?      @      �?      @      �?      @              @      �?                              �?      �?      @      &@      @               @              $@      .@              "@              *@      @      $@      @      @              $@      ,@      @      .@      @      .@      @     �T@     �P@      E@      ^@      4@      W@      @      O@      (@      S@     �E@      4@      "@     �B@      N@      9@     �U@      Z@     �[@      3@      A@      ;@      :@     �M@      $@      D@      @      7@      "@     �@@      =@      &@      �?      3@      6@      &@      D@      C@      H@      @      A@      ,@      7@     �M@      "@      D@      @      5@      "@     �@@      <@      &@              0@      5@      &@      C@      A@      G@      @              *@      @              �?                       @                      �?              �?      @      �?               @      @       @             �H@      D@      0@     �N@      $@      J@             �C@      @     �E@      ,@      "@       @      2@      C@      ,@      G@     �P@     �O@      ,@      "@      0@      @      2@      @      6@              @              @              �?              $@      ,@      @      @      ,@      <@      @      D@      8@      &@     �E@      @      >@              @@      @     �C@      ,@       @       @       @      8@       @     �C@      J@     �A@      @     �i@     �Q@      6@     �i@      @     �v@             �W@      .@     �s@     �M@      >@      ,@      :@     @_@      =@     `k@      f@     @r@     �C@      N@      2@      @     �V@             `f@             �G@              e@      3@      @      �?      @     �M@      $@     �U@      Q@     @b@      $@      B@      .@      @     @R@             �b@              C@             �`@      (@      @      �?      @      G@      @     �R@     �L@      `@      @      1@       @      @      J@             @_@              A@             @\@      "@      @      �?      �?      A@      �?      O@      >@     �Z@      @      3@      @              5@              8@              @              5@      @                       @      (@      @      *@      ;@      7@      @      8@      @      �?      2@              >@              "@             �A@      @                       @      *@      @      &@      &@      1@      @      1@      @              &@              .@              �?              4@      @                              *@      @      &@      @      &@      �?      @              �?      @              .@               @              .@                               @                              @      @       @     `b@      J@      1@     @\@      @     `g@              H@      .@     �a@      D@      7@      *@      5@     �P@      3@     �`@      [@     @b@      =@     �R@      5@       @      L@      �?     �X@              8@      (@     @S@      ;@      "@      @       @      =@      "@      E@     �J@      P@      0@      *@      @              0@              8@              "@              5@      $@      @      @      @      @      �?      1@      6@     �C@      @     �N@      ,@       @      D@      �?     �R@              .@      (@      L@      1@      @      @       @      8@       @      9@      ?@      9@      $@     @R@      ?@      .@     �L@      @      V@              8@      @     �P@      *@      ,@      @      *@     �B@      $@     �V@     �K@     �T@      *@     �P@      >@       @     �J@      @     �U@              4@      @     �N@      $@      ,@      @      @      B@      $@      U@      J@     @S@      *@      @      �?      @      @              �?              @              @      @                      @      �?              @      @      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJF�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�M��.�@�	           ��@       	                    �?��"ѡ@:           `�@                          �9@�@]a@2@<           �@                           �?I�B��@�            px@������������������������       ��6~a)@`            �c@������������������������       �*�+L�@�            `m@                          �?@Z��+@K            �]@������������������������       �_��PW�@>            �W@������������������������       �����5E@             7@
                           @�X�h��@�           ؈@                           @ `맫k@�            `v@������������������������       �6���"�@�             i@������������������������       ��8�@V            �c@                            �?��i��
@           P{@������������������������       �w�;R��
@�             o@������������������������       ��E�4R
@�            �g@                           �?��&
�@r           b�@                          @A@�2�T@�           ��@                           �?+�%E/�@�           ��@������������������������       ��z8�@�            �s@������������������������       ��V	e��@�            �@                          �A@���Nf;@            �A@������������������������       ��HSvݤ@             2@������������������������       �"�]䁀�?             1@                          �4@e��q��@�           @�@                           @횉M'@�           8�@������������������������       ���`�@�           `�@������������������������       ��jx$��	@;            �V@                           @�٫L�y@�           H�@������������������������       �8K��s@           �{@������������������������       ��x�S@�            s@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �`@     �X@     @v@      B@     �~@      "@      k@      :@     �z@      ]@      O@      :@     �R@     �l@     �N@     �w@     �s@     |@     �S@      Y@      ;@      >@     �X@      "@     @i@       @     �V@      "@     �c@      ?@      ,@      @      3@     �Q@      "@     @a@      Z@      c@     �B@      B@      ,@      6@     �A@      @      I@       @      C@       @      C@      4@      &@      @      *@      ?@      @     �Q@     �E@      K@      $@      >@       @      .@      >@       @      G@              @@      @      B@      ,@      @      �?      &@      1@              M@      =@     �F@       @      $@               @      0@              4@              @      @      &@      $@      �?                      @              0@      0@      ;@      @      4@       @      @      ,@       @      :@              9@      @      9@      @       @      �?      &@      $@              E@      *@      2@      @      @      @      @      @       @      @       @      @       @       @      @       @      @       @      ,@      @      *@      ,@      "@       @       @      @      @      @       @      �?       @      @       @       @      @      @      @              ,@      @      &@      ,@      "@       @      @      @      @      �?              @                                              @               @              �?       @                              P@      *@       @     �O@      @      c@             �J@      �?     �]@      &@      @              @      D@      @     �P@     �N@     �X@      ;@      7@      @      @      ;@      @     �Q@              8@              I@      @      @              @      2@      �?      ?@      8@      C@      6@      0@      @              0@       @      >@              2@             �@@      @      �?                      @      �?      *@      ,@      ;@      ,@      @       @      @      &@      �?     �D@              @              1@      �?       @              @      &@              2@      $@      &@       @     �D@       @      �?      B@       @     @T@              =@      �?     @Q@      @                      �?      6@      @      B@     �B@      N@      @      6@      @      �?      7@       @      G@              5@      �?     �C@       @                      �?      @       @      7@      4@      A@              3@       @              *@             �A@               @              >@      @                              0@      �?      *@      1@      :@      @     �l@      [@      Q@      p@      ;@      r@      @     �_@      1@      q@     @U@      H@      6@     �K@     �c@      J@     �m@      j@     �r@      E@     @V@     �J@      F@     �[@      4@     �U@      @      M@      $@     @Y@      C@      7@      ,@      B@     �R@      <@      S@      Y@      _@      =@     @V@     �F@      C@     @[@      4@     �U@      @     �L@      $@     �X@      >@      6@      (@      B@     @R@      <@     �R@     �X@      _@      =@     �F@      @      (@      ?@      &@      :@              .@      @      :@      "@       @      @      @      (@      @      ;@      1@      F@       @      F@     �C@      :@     �S@      "@     �N@      @      E@      @     @R@      5@      4@      @      >@     �N@      5@      H@     @T@      T@      5@               @      @       @                              �?               @       @      �?       @               @              �?       @                              @      �?       @                                               @      �?      �?       @               @              �?      �?                              @      @                                      �?                      @                                                      �?                     �a@     �K@      8@     `b@      @      i@       @      Q@      @     �e@     �G@      9@       @      3@      U@      8@     @d@      [@     �e@      *@     �H@      6@      $@      T@      �?      [@             �B@             @X@       @      ,@      @             �E@      *@     �W@     �G@      [@      @     �C@      5@      $@     �S@             �V@              <@              W@      @      &@      @              D@      &@     @R@      E@     �X@      @      $@      �?               @      �?      2@              "@              @      �?      @                      @       @      5@      @      $@              W@     �@@      ,@     �P@      @     @W@       @      ?@      @      S@     �C@      &@      @      3@     �D@      &@      Q@     �N@     @P@      @      L@      6@      @      E@      @     �N@              ;@      @      D@      8@      @      @      @      ;@      $@     �D@      ?@      7@      @      B@      &@      "@      9@       @      @@       @      @              B@      .@      @              *@      ,@      �?      ;@      >@      E@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�v�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�]�Em�@�	           ��@       	                    �?/L+�@           �@                          �6@W ��D@j           8�@                           @���]V{@�            �t@������������������������       �Y�-?@�             o@������������������������       �.M�eZ�
@>            �U@                           @��C"�@�             o@������������������������       �x<g�O@N            ``@������������������������       ����v*1@E            @]@
                          �;@����@�           Ԑ@                           @�9~Rk@<           �@������������������������       �#�����@           X�@������������������������       �<E8��@9            �U@                           @��U�m�@k            �f@������������������������       ����
4@M            ``@������������������������       �8�>>�Y@            �H@                           �?�v1��d@�           ��@                           �?JXS�7@�           ��@                          �9@~��͌@           p{@������������������������       ��+�;�@�            Pw@������������������������       �	��5)@*            �P@                           @h~x�@�            �u@������������������������       �.�R�S
@�            q@������������������������       �}o,�]F
@0            @R@                           @zd���@�           �@                            �?�s�ٍ@$           l�@������������������������       ������@�            �x@������������������������       �qq4�@-           ��@                           @�H��7q@j             d@������������������������       ��$�lz@Q             ^@������������������������       ���1�h�	@            �D@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �a@     @T@     �v@      C@     0|@      *@     �m@      <@     @|@      U@      L@      J@     �M@     @o@     @R@     �v@     pt@      {@      W@     @a@     �Q@     �K@      b@      :@     @a@      "@     �`@      6@     �b@     �J@      @@      =@     �D@     @X@      C@     �`@     �b@     �d@      B@      G@       @      8@      A@      $@     �P@      @      H@      @      M@      3@      @      $@      "@      B@      .@      L@      I@     @P@      (@      A@      @      @      1@      @      J@              ;@              A@      .@      @      @      @      3@      @     �@@      :@      E@       @      .@       @       @      @      @      D@              1@              =@      (@      @      @      @      .@      @      @@      1@      A@      @      3@      �?       @      $@              (@              $@              @      @      �?                      @      �?      �?      "@       @      �?      (@      @      4@      1@      @      .@      @      5@      @      8@      @       @      @      @      1@      $@      7@      8@      7@      @      @      @       @      @       @      ,@      @      1@      @      "@      �?       @      @      @      @      @      "@      .@      $@      @       @              (@      &@      @      �?              @              .@      @               @       @      (@      @      ,@      "@      *@      �?      W@     �O@      ?@     �[@      0@     �Q@      @      U@      3@      W@      A@      9@      3@      @@     �N@      7@      S@     @Y@      Y@      8@     �T@      B@      9@     �W@      0@      P@      @      Q@      3@     �T@      <@      2@      $@      ;@      J@      5@     �P@     �Q@      V@      8@     �S@     �A@      8@     �U@      0@      J@      @      N@      3@     @S@      <@      .@      $@      5@     �F@      (@      N@     �N@      U@      8@      @      �?      �?       @              (@               @              @              @              @      @      "@      @      "@      @              "@      ;@      @      0@              @              0@              "@      @      @      "@      @      "@       @      "@      ?@      (@               @      6@      @      *@              @              &@              @      @      @      @      @      "@       @       @      .@      @              �?      @      �?      @              �?              @              @              �?       @      �?                      �?      0@       @             �f@     @Q@      :@     `k@      (@     �s@      @      Z@      @     �r@      ?@      8@      7@      2@      c@     �A@     `m@      f@     �p@      L@     �O@      &@      $@     �P@      @      _@             �D@              Z@      "@      @              @     @Q@      @     �R@      N@     @Z@      :@      E@      @       @      ?@      @     �O@              <@             @P@      @      @               @      E@       @      ;@      @@      L@      3@     �C@      @      @      :@      @     �M@              9@              I@      @                       @     �C@              6@      :@      J@      .@      @              @      @      @      @              @              .@      �?      @                      @       @      @      @      @      @      5@      @       @     �A@             �N@              *@             �C@      @                      @      ;@      @      H@      <@     �H@      @      ,@      @      �?      ?@              N@               @              <@       @                      �?      4@      @      D@      3@      A@      @      @              �?      @              �?              @              &@      �?                       @      @       @       @      "@      .@             @]@      M@      0@      c@      @     �g@      @     �O@      @     �h@      6@      5@      7@      *@      U@      <@      d@      ]@     @d@      >@     �Y@      F@      ,@     �a@      @     @e@      @      M@      @      f@      1@      3@      1@      *@     @P@      7@     `b@     �Y@      c@      >@      =@      .@      "@     �F@             �N@              $@              F@       @      @      "@      @      ,@      @      H@      1@     �M@      @     @R@      =@      @     �X@      @     @[@      @      H@      @     �`@      "@      *@       @      @     �I@      1@     �X@     @U@     @W@      8@      .@      ,@       @      $@      �?      3@              @              5@      @       @      @              3@      @      *@      ,@      $@              (@      ,@       @      @              1@              @              &@      @       @                      0@      @      (@       @      @              @                      @      �?       @              �?              $@                      @              @      �?      �?      @      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�d/hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@OG��@�	           ��@       	                    �?�c���d@D           ޠ@                            @�YOX�@x           ��@                           �?=��7{%@�           �@������������������������       ��"�Eз@3             W@������������������������       �L�ݴP�@�           8�@                          �1@��P�@�            �q@������������������������       ��?�'�@:            �W@������������������������       ��/��@�            �g@
                           �?_$�C۾@�           ��@                            @eI��̡@           P{@������������������������       �|0)�w@�             r@������������������������       �F⹿��@`            �b@                          �3@r�8��v@�           ؅@������������������������       �t��m_�@           �{@������������������������       ��J����@�             p@                           �?�?���@d           h�@                           �?}�V}�[@<            �@                           @'��c@�            �p@������������������������       ������r@x            �g@������������������������       �j����?@4             T@                           �?A�l�W]@�           ��@������������������������       �\����@�            �k@������������������������       ����/h@           �{@                          �;@0V���@(           ��@                           @��i�W@�           ��@������������������������       �d8���-@�           ȁ@������������������������       �F�Ƅ�@,            �P@                           @,�wfe�@u            @g@������������������������       �+# S�@9            �X@������������������������       ���6��@<             V@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       `s@     �`@     �T@     �t@      D@     �|@       @     `k@     �B@     0~@     �V@     �P@     �A@     @S@     �m@     �P@     0w@     �s@     `}@     @T@     �c@     �H@      A@     �g@      1@     �r@             �^@      (@     @r@     �A@      E@      .@      7@     @Z@      ?@     `k@     @f@     �r@     �B@     @S@      5@      (@     �S@      @      c@              K@             @`@      2@      2@      $@       @      F@      $@      Z@     @V@      e@      7@     �@@      .@      @      G@      @     @]@             �B@             �Y@      $@      .@       @      @     �A@      @     �S@     �O@     @a@      2@      "@              �?      "@       @      $@              �?              @       @       @              @       @              @      ,@      2@      @      8@      .@      @     �B@      �?     �Z@              B@             @X@       @      *@       @      @     �@@      @     @R@     �H@      ^@      &@      F@      @      @      @@      @     �A@              1@              ;@       @      @       @      �?      "@      @      :@      :@      >@      @      0@      @      @      *@      �?      *@              @              @      @                      �?      �?       @      &@      @      @       @      <@              @      3@      @      6@              ,@              5@       @      @       @               @      �?      .@      4@      9@      @     �S@      <@      6@      \@      $@     �b@             @Q@      (@     @d@      1@      8@      @      .@     �N@      5@     �\@     @V@     ``@      ,@     �G@      "@      *@      J@       @      C@              <@      "@     �F@       @      .@      �?      "@      8@       @      =@     �D@     �H@      $@      @@      @       @     �H@              7@              "@       @      @@               @              @      0@      @      0@      7@      A@      "@      .@       @      @      @       @      .@              3@      �?      *@       @      @      �?       @       @      �?      *@      2@      .@      �?      @@      3@      "@      N@       @      \@             �D@      @     @]@      .@      "@      @      @     �B@      *@     �U@      H@     �T@      @      6@      "@      @     �C@             �P@              :@      �?      V@      .@      @      �?      @      6@      "@      H@      7@     �L@              $@      $@      @      5@       @     �F@              .@       @      =@              @      @              .@      @      C@      9@      9@      @     @c@     �T@     �H@     �a@      7@     `c@       @      X@      9@     �g@     �K@      9@      4@      K@     ``@     �A@      c@     �a@     `e@      F@      M@      J@     �@@      R@      4@     �P@       @     �Q@      4@      T@      @@      5@      1@      C@     �M@      0@     �Q@      V@     @U@      :@      2@      0@      0@      5@      �?      B@       @      ,@      @      4@      @      @       @      $@      :@      @      0@      .@      ?@      @      1@      $@      *@      .@              <@       @      (@      @      &@      @      @      �?      @      (@       @      $@      $@      3@      @      �?      @      @      @      �?       @               @              "@                      �?      @      ,@      @      @      @      (@              D@      B@      1@     �I@      3@      ?@      @      L@      .@      N@      :@      .@      .@      <@     �@@      &@      K@     @R@      K@      7@      @      (@      @      &@      @      1@              1@      @      ;@      (@       @       @       @      *@      @      1@     �C@      &@      (@     �B@      8@      *@      D@      .@      ,@      @     �C@       @     �@@      ,@      *@      *@      4@      4@       @     �B@      A@     �E@      &@      X@      ?@      0@     �Q@      @      V@              :@      @     �[@      7@      @      @      0@      R@      3@     �T@     �J@     �U@      2@      R@      8@       @     �N@      �?     �Q@              8@       @     �U@      *@      @      �?      $@     �M@      *@     �Q@      D@     �M@      2@     �N@      6@       @     �L@      �?      P@              5@       @     �T@      $@      @              $@     �H@      "@      Q@      @@     �I@      2@      &@       @              @              @              @              @      @              �?              $@      @       @       @       @              8@      @       @      "@       @      2@               @      @      8@      $@               @      @      *@      @      (@      *@      ;@              ,@      @       @      @      �?       @              �?              5@      @                      @      @      @      @      @      &@              $@      @      @       @      �?      $@              �?      @      @      @               @       @      @              "@      "@      0@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�ehG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@
@�2�@�	           ��@       	                     @�uS���@n            �@                           @��;!�)@�           ��@                          �0@'��*��@�            �v@������������������������       �w�PC,�@*             L@������������������������       �'�˵�@�            s@                            �?�Q�
@�           P�@������������������������       ���i$�
@           �{@������������������������       �W�3d��@q            �e@
                          �2@ً�4W@�            Pw@                           @���]@�            �p@������������������������       � ^�7�p@�            �i@������������������������       ����1@&            �O@                           �?���s�
@?            �Y@������������������������       ���Q�4	@             J@������������������������       ���Lu�	@             �I@                          �<@-��%t@>           �@                           @iEc�C@x           ��@                           �?3���&@`           J�@������������������������       �iJ��@c           ��@������������������������       �׏	jm�@�           <�@                           �?/6��g�	@             B@������������������������       ��	�o�� @             $@������������������������       ���n#�@             :@                           @�\v�Vq@�            �s@                           �?�c��h@g            �c@������������������������       �0#dA�@7             U@������������������������       ��ݧ=@0             R@                           @��d�a@_            �c@������������������������       �E�x�m@N            �_@������������������������       �K2��0@             =@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@      _@     �T@     �v@      E@      }@       @     �i@     �A@     �{@      ^@      N@      E@     �M@      o@      S@     �v@     `s@     �|@     �U@     �S@      :@     �@@      ^@      @     �i@       @     �T@      @     �g@      ?@      .@      @      "@     �Q@      5@     @_@     @Y@     @j@      1@     �F@      5@      6@      V@       @     �a@             �I@      @      c@      .@      $@      @      @     �M@      ,@      U@     @R@     @f@      (@      2@      "@      ,@      D@       @      >@              2@      @      F@      $@      @      @      @      6@      @      :@      <@     �Q@      "@       @                      &@              @              "@              @                              @      @               @      "@       @              0@      "@      ,@      =@       @      8@              "@      @     �D@      $@      @      @      @      3@      @      8@      3@      O@      "@      ;@      (@       @      H@             �[@             �@@              [@      @      @      �?             �B@      "@      M@     �F@      [@      @      3@      &@      @      A@             @P@              9@              V@      @       @      �?              >@      "@      H@      ;@      R@       @       @      �?       @      ,@             �F@               @              4@      �?      @                      @              $@      2@      B@      �?      A@      @      &@      @@      @     �P@       @      @@              C@      0@      @              @      &@      @     �D@      <@      @@      @      6@      @      @      <@      @     �E@       @      :@              >@       @      @                      $@      @      @@      3@      3@      @      *@      �?       @      6@      @     �@@       @      7@              7@      @      �?                      "@      @      <@      0@      0@      @      "@      @      @      @              $@              @              @      �?      @                      �?      @      @      @      @       @      (@              @      @              7@              @               @       @                      @      �?      �?      "@      "@      *@              @               @       @              ,@              @              @      @                              �?      �?      @      �?      @              @              @       @              "@               @              �?      @                      @                      @       @       @             �m@     �X@     �H@     @n@     �A@     @p@      @     �^@      @@     p@     @V@     �F@      C@      I@     `f@     �K@      n@      j@     �n@     @Q@      j@     �R@      C@     �j@      =@      o@      @     �[@      @@     �l@      S@      E@      9@      E@      d@     �G@      l@      e@     �j@      O@      j@     �Q@      C@     �j@      8@     �n@      @      [@      @@     @l@      S@      E@      4@      E@     @c@      F@     �k@     �d@     �j@      O@     �V@      @@      6@     �V@      0@     @Q@      @      L@      9@     �X@      C@      >@      &@      >@     �O@      7@     �X@     �M@     �V@      A@     �]@      C@      0@     @_@       @     @f@              J@      @     �_@      C@      (@      "@      (@     �V@      5@     @^@      [@     �^@      <@              @                      @      �?               @              @                      @              @      @      @      �?      �?                                                      �?                               @                                      @               @              �?                      @                      @                       @              �?                      @               @      @       @      �?                      >@      7@      &@      ;@      @      (@      �?      (@              <@      *@      @      *@       @      3@       @      1@     �D@     �@@      @      1@      0@      @      @      @       @      �?      @              4@      @      @       @      @      *@      @       @      .@      @              @      @      @      �?      @      @               @              "@      @      @      @      @      @       @       @      .@      @              (@      $@      �?      @       @       @      �?      @              &@       @              �?       @       @      @      @              �?              *@      @      @      4@      �?      @              @               @      @              @      @      @       @      "@      :@      :@      @      &@      @      @      4@              @              @              @      @              @       @      @       @      @      3@      1@      @       @                              �?                                      �?       @                      �?                      @      @      "@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ2ڪshG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@˝_ʿ�@�	           ��@       	                     @��ӭ@@x           ��@                          �0@��k*��@<           ��@                           @$8bMT5@^             c@������������������������       �x
�o�@F             \@������������������������       ��gA��@            �D@                           �?*���u@�           D�@������������������������       �-DP�a�@Q           0�@������������������������       �~��Ff�@�           X�@
                           �?�鳱@<           �@                           �?I�z��@�            �n@������������������������       �����!@O            �`@������������������������       ��U��/�	@F             \@                           @��6x��@�            �p@������������������������       ��H�tШ@~            �h@������������������������       �jz��
@)            �Q@                            @�WLѾi@O           ��@                           �?vP���@�           �@                           �?�Oz��@D           �@������������������������       �SP�o@�@�             o@������������������������       ��/>�C@�            0p@                          �9@���r� @z           P�@������������������������       ���dB�[@�           (�@������������������������       ��趸^w@�            Pv@                           @����@�           ��@                           @>�ŕ/@b           x�@������������������������       ��l])�@[            �@������������������������       ��QUL>. @             .@                           @��Ω��	@/            @R@������������������������       �y"|GT@            �C@������������������������       �Ij�Q��@             A@�t�b��     h�h5h8K ��h:��R�(KKKK��h��B`       s@     `a@     �V@     `v@     �F@     ~@      @     @k@      5@     `@     �\@      K@     �D@     �U@     Pp@      M@     pt@     �p@     �|@     �U@     �\@     �C@      E@     �c@      0@     0p@              V@       @      p@     �D@      6@      @      4@      [@      :@      b@     @]@     �p@     �@@      R@      A@      7@     �\@      @     �h@              L@      @      g@      1@      1@      @      &@     �U@      ,@     @X@     @U@      j@      9@       @       @              *@             �A@              @              0@               @              �?      &@       @      *@      $@      D@               @                      @              ;@              @              .@              �?              �?       @       @      (@      @      ?@                       @              $@               @              �?              �?              �?                      @              �?      @      "@             �Q@      @@      7@     @Y@      @      d@              I@      @      e@      1@      .@      @      $@     �R@      (@      U@     �R@      e@      9@      ;@      ,@      "@     �D@       @      T@              :@             �V@       @       @      @      �?     �C@      @      @@     �D@     @U@      *@     �E@      2@      ,@      N@      @     @T@              8@      @     �S@      "@      *@      �?      "@      B@      "@      J@      A@      U@      (@      E@      @      3@      F@      $@     �O@              @@       @     @R@      8@      @       @      "@      6@      (@      H@      @@      O@       @      ;@      �?      @      ?@      @      =@              .@              =@      (@      �?              @      @      @      6@      &@     �C@      @      0@      �?      @      .@       @      ,@               @               @      (@      �?              @      @      �?      0@       @      1@      �?      &@               @      0@      �?      .@              @              5@                                       @      @      @      @      6@      @      .@      @      *@      *@      @      A@              1@       @      F@      (@      @       @      @      .@       @      :@      5@      7@      @      @      @      &@      &@      @      =@               @       @      ;@      (@       @       @      �?      ,@      @      1@      .@      4@      @      "@               @       @              @              "@              1@               @              @      �?      �?      "@      @      @             �g@      Y@      H@      i@      =@     �k@      @     @`@      *@     �n@     @R@      @@      A@     �P@      c@      @@     �f@     `b@     `g@     �J@      a@     @Q@     �@@     ``@      *@     @g@      �?     �R@      @     �f@      E@      3@      8@      G@     �Y@      6@      _@     �V@      a@     �B@     �B@      5@      2@      D@       @     @T@              =@             @P@      ,@      @      @      &@      7@      @     �E@     �B@     �K@      2@      7@      $@      @      3@              G@               @              B@      @      �?      �?      @      $@       @      4@      0@      9@      ,@      ,@      &@      (@      5@       @     �A@              5@              =@      @      @      @      @      *@      �?      7@      5@      >@      @      Y@      H@      .@     �V@      &@     @Z@      �?      G@      @     @]@      <@      *@      4@     �A@     �S@      3@     @T@      K@     @T@      3@      R@      9@      @     �P@       @     @Q@      �?      .@       @      T@      3@      "@      "@      6@      N@      "@      M@     �@@      B@      *@      <@      7@       @      9@      @      B@              ?@      @     �B@      "@      @      &@      *@      3@      $@      7@      5@     �F@      @      K@      ?@      .@     @Q@      0@      B@      @     �K@      @      O@      ?@      *@      $@      4@     �I@      $@      M@      L@     �I@      0@     �H@      9@      .@     �M@      0@      @@      @     �K@      @      I@      <@      *@      $@      4@     �B@      $@     �K@     �J@     �D@      *@     �H@      9@      .@     �M@      *@      @@      @     �K@      @      I@      <@      *@      $@      4@      ?@      $@     �I@      J@      D@      *@                                      @                                                                              @              @      �?      �?              @      @              $@              @                              (@      @                              ,@              @      @      $@      @       @      @              @               @                              @      @                              @              �?               @      �?      @                      @               @                               @                                      @               @      @       @       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�b�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��TP�@�	           ��@       	                    �?`���BF@           :�@                            @!K�00�@~           X�@                           �?s$>�6@~           ��@������������������������       ������@�             m@������������������������       ��\r,`�@�            @w@                          �5@o�A�@            �x@������������������������       �G;�mA@o             f@������������������������       ��gP��n@�            �k@
                          �5@�t^��@�           Ȗ@                          �3@�h�Q~w@d           ��@������������������������       �����
@�           ��@������������������������       ���"$�@�            �q@                           @oM��&�@.           �}@������������������������       ���Gڭ@�            �v@������������������������       �_|�=\5
@J            �\@                          �3@%d� 9@�           ��@                          �2@��c�@           `{@                           @��U��@�            Pu@������������������������       �C,�Cv@y            �g@������������������������       ��j���@Y             c@                            �?�q�V�!@?            @X@������������������������       �m�XY�l@             9@������������������������       ��-���@0             R@                          �;@s�8o�@�           ��@                           @����<y@           P�@������������������������       ��" �8�@�            �r@������������������������       ��U���@N           �@                           �?6N�V@}            �i@������������������������       ���/C�>@J             ^@������������������������       �'�.X�@3             U@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �r@     `b@      V@     �v@      ?@     P|@      &@      j@     �A@     P|@     @Y@      I@      H@      O@      o@     @R@     �w@     �r@     @}@     �V@      g@     @S@      I@     �k@      2@     �s@      $@     @a@      ,@     Pt@     @P@      :@      :@      C@     @b@      ?@     �n@     �f@     �q@     �O@     �P@      C@     �@@      U@      *@      W@      $@     @R@      @     �X@      =@      ,@      3@     �@@     �L@      3@     �Y@     @W@     @W@      >@      C@      8@      ,@      M@      @     �J@       @     �E@      @      R@      ,@      $@      $@       @      B@      &@     @P@      I@      O@      5@      $@      @      "@      &@      @      8@      @      0@             �A@      @      @       @      �?      ,@      @      5@      ;@      :@      @      <@      2@      @     �G@              =@      �?      ;@      @     �B@       @      @       @      @      6@       @      F@      7@      B@      .@      <@      ,@      3@      :@      "@     �C@       @      >@      @      :@      .@      @      "@      9@      5@       @     �B@     �E@      ?@      "@      4@      �?      @      $@      @      7@      �?      0@              "@      @      �?      �?      @      "@      @      6@      6@      3@               @      *@      ,@      0@      @      0@      �?      ,@      @      1@      $@      @       @      5@      (@      @      .@      5@      (@      "@     �]@     �C@      1@     @a@      @     `l@             @P@      @     `l@      B@      (@      @      @     @V@      (@     �a@     �U@      h@     �@@      K@      5@      &@     @Y@              e@             �H@       @     `d@      1@       @      @       @     �D@      @     @Z@     �P@     �a@      3@      B@      (@       @     @S@             �^@             �@@       @     �`@      *@      @               @      9@      @     �Q@     �@@     �[@      &@      2@      "@      @      8@              G@              0@              >@      @      @      @              0@      @      A@     �@@     �@@       @      P@      2@      @     �B@      @     �M@              0@      @      P@      3@      @       @      @      H@      @     �B@      5@     �H@      ,@      L@      "@      @      >@      @     �J@              0@      @     �F@      .@      @       @      @     �@@      @      9@      0@      8@      *@       @      "@      @      @              @                              3@      @      �?                      .@              (@      @      9@      �?     @]@     �Q@      C@      b@      *@     �`@      �?     �Q@      5@      `@      B@      8@      6@      8@     �Y@      E@     �`@     �^@     �f@      ;@      F@      ,@      (@     �C@              M@              2@              @@      (@      @               @      C@      (@      8@      D@     @S@      "@      C@      &@      "@      ?@              E@              0@              >@       @      @               @      :@      "@      &@      ?@     �P@      @      7@       @      @      6@              ,@              @              0@      @      @               @      ,@      @      @      8@     �A@      @      .@      "@       @      "@              <@              $@              ,@      @      �?                      (@      @       @      @      ?@              @      @      @       @              0@               @               @      @                              (@      @      *@      "@      &@      @      �?      �?                              @              �?                      �?                                              @       @      @      @      @       @      @       @              (@              �?               @      @                              (@      @      $@      @      @             @R@      L@      :@     �Z@      *@      S@      �?      J@      5@      X@      8@      1@      6@      6@      P@      >@      [@     �T@     �Z@      2@      M@     �E@      0@     �U@      &@      Q@              @@      5@     @S@      2@      ,@      2@      2@     �M@      8@      X@     �N@     �S@      (@      *@      ,@      @      G@       @      5@              *@      (@      4@      @      "@      (@       @      1@       @      ;@      8@      =@      @     �F@      =@      &@      D@      @     �G@              3@      "@     �L@      &@      @      @      $@      E@      0@     @Q@     �B@     �H@      @      .@      *@      $@      4@       @       @      �?      4@              3@      @      @      @      @      @      @      (@      6@      <@      @       @      *@      @      .@       @      �?              ,@               @      �?      @      @       @      @      @      @      ,@      (@       @      @              @      @              @      �?      @              &@      @                       @       @       @      @       @      0@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�!PehG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���ㆱ@�	           ��@       	                   �4@�ގ@           ��@                            �?�Ѷ�$$@v           �@                          �3@���4��@�            0r@������������������������       �)�e�B@�            �j@������������������������       ��C��%*@3            @S@                          �3@�Y(���@�            �s@������������������������       �I3�p!�@�            �l@������������������������       �tT3/ƪ@+            �T@
                           �?<V�0J@�           ,�@                          �:@��-���@�            v@������������������������       �0��0E�@�            pp@������������������������       �T
��v@<            �V@                            �?n��H�@�           P�@������������������������       �dÓ�@�            `g@������������������������       �u�\K�@4           �~@                           �?_���8@�           ¡@                          �3@"텆�/@�           \�@                            �?�S$�p`
@?           �@������������������������       ��M���
@�            pt@������������������������       �����	@t            `g@                           �?��8G��@�           ��@������������������������       ��ϭ���@�            �o@������������������������       � ��-:@�            �u@                          �6@�W(�F�@�           (�@                          �2@F����@�           �@������������������������       ���#[�@�            �u@������������������������       �3�~��@           �{@                          �7@�}���@�            �v@������������������������       �զ��}@6            @U@������������������������       �^�%�d@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        s@     �a@     @X@     0u@      E@     }@      @     �k@      B@     �{@     @X@      M@      :@     �R@     @o@      S@     pw@     �u@     �{@     @Q@      a@     �Q@     �K@     �`@      ;@     @`@      @      ^@      7@     @d@      L@     �B@      0@      M@     @[@     �@@     �b@     �a@      a@      C@      Q@      "@      8@     �G@      $@     �K@       @      <@      @     �L@      8@      .@      @       @     �H@      @      I@     �L@     �O@      7@      <@      @      *@      =@              =@              *@      @     �C@      @      $@              @      .@      @      .@      :@     �D@      &@      2@       @      (@      :@              6@              @      @      7@      @      $@              @      "@       @       @      4@      C@      @      $@      @      �?      @              @              @              0@      �?                      �?      @       @      @      @      @      @      D@      @      &@      2@      $@      :@       @      .@      �?      2@      4@      @      @      @      A@       @     �A@      ?@      6@      (@      9@      @      &@      (@      @      9@       @      ,@              (@      (@      @       @      �?      :@      �?      ?@      ;@      .@      @      .@                      @      @      �?              �?      �?      @       @       @      @       @       @      �?      @      @      @      @     @Q@     �N@      ?@      V@      1@     �R@      @      W@      2@     @Z@      @@      6@      &@      I@      N@      ;@     �X@     @U@     �R@      .@      9@      "@      *@      8@       @      5@       @      @@      @      =@      *@       @      @      7@      ?@      @      B@      >@      @@      @      6@      @      @      6@      @      3@      �?      2@       @      8@      @       @              2@      2@       @      >@      =@      6@      @      @      @      @       @      @       @      �?      ,@      @      @      @              @      @      *@       @      @      �?      $@              F@      J@      2@      P@      "@      K@       @      N@      (@      S@      3@      ,@       @      ;@      =@      7@     �O@     �K@      E@      &@      "@      ,@       @      6@      @      ,@      �?      1@      "@      2@      @      @       @      @      @      @      .@      2@      *@      @     �A@      C@      0@      E@      @      D@      �?     �E@      @      M@      0@      &@      @      5@      7@      3@      H@     �B@      =@      @     �d@     �Q@      E@     �i@      .@     �t@             �Y@      *@     �q@     �D@      5@      $@      0@     �a@     �E@     @l@     �i@      s@      ?@     �U@      @@      .@     �W@      $@     @f@              J@      (@     @`@      8@      $@      @      @     �Q@      *@      W@      ]@     �a@      9@      >@      @             �F@       @     �W@              <@             @R@      �?      @       @              =@       @     �I@     �I@     �U@       @      2@      @              @@       @     �L@              2@              N@              �?       @              4@              =@      ?@      G@      @      (@       @              *@              C@              $@              *@      �?      @                      "@       @      6@      4@      D@      �?     �L@      :@      .@      I@       @     �T@              8@      (@     �L@      7@      @       @      @      E@      &@     �D@     @P@      L@      1@      6@      @      &@      ,@      @     �A@              0@              <@      &@       @               @      8@      @      1@      :@      8@      "@     �A@      5@      @      B@      @      H@               @      (@      =@      (@      @       @      �?      2@       @      8@     �C@      @@       @      T@     �C@      ;@     @[@      @     �c@             �I@      �?     @c@      1@      &@      @      *@     �Q@      >@     �`@     �V@     @d@      @      F@      5@      2@     �R@      @     @^@              F@      �?     �Y@      @      &@       @       @     �H@      2@     �X@      N@     @[@      @      9@      $@      @      >@              P@              3@             �I@      @       @       @      @      *@      (@     �C@      9@      G@              3@      &@      ,@     �F@      @     �L@              9@      �?      J@      @      "@               @      B@      @      N@     �A@     �O@      @      B@      2@      "@      A@       @      B@              @             �I@      $@              @      @      5@      (@     �A@      >@     �J@       @      1@      @      @      @              @              �?              &@      @                      �?      �?       @      *@      "@      @       @      3@      .@      @      <@       @      @@              @              D@      @              @      @      4@      @      6@      5@      I@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�;�+hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?D��:�@�	           ��@       	                     @{XG5��@            �@                          �5@��� �@u           ��@                           @a��,@           pz@������������������������       ��P{K�@�            �q@������������������������       ��G�023@Y            �a@                          �6@Z� $6 @j           X�@������������������������       ���O��@4             V@������������������������       �mX���@6           0@
                           @��C��@�           P�@                           �?�����@�            s@������������������������       ��6R���@1             S@������������������������       �e}3ZxX@�            �l@                          �<@� %ݵ@�            �u@������������������������       ���W>p@�            �r@������������������������       ��ٺ?Q@#            �H@                           @H4��y\@�           ��@                           @g���W@N           ؚ@                          �5@-))8&@�           H�@������������������������       �;Tʄ�@�           ��@������������������������       ���%�@f           ؁@                          �9@�Z웖<@h            �d@������������������������       �f��آ@W            �`@������������������������       �X"�P��@             >@                          �5@�/$ƞ�@Z           ��@                           �?3S_�(@�            �r@������������������������       �����@P            �_@������������������������       �����3@p            �e@                          �8@p���@�            �m@������������������������       �b L�� @G            �]@������������������������       �^��)5@S            �]@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �a@     @V@     `v@     �@@      |@      @      k@      7@     �|@     �X@      L@     �@@     @R@     �p@     �Q@     `y@     �r@     {@     �U@     �^@      S@      N@     �c@      7@      a@      @     @Y@      0@     �b@     �L@      =@      3@     �I@      Y@      @@     �f@     �a@     @d@      C@     �S@      H@     �@@      \@      "@     @U@      @     �K@      $@     @Y@      =@      4@      (@      9@      N@      8@     @Y@     �P@     @[@      :@     �E@      ,@      (@     �K@             �A@              0@      "@     �H@      &@      "@      �?       @      5@      @     �B@     �B@      I@      &@      9@      @       @      H@              4@              "@      @     �C@      @      @      �?      @      (@      �?      <@      ;@      A@      @      2@      @      $@      @              .@              @       @      $@      @      @              @      "@      @      "@      $@      0@      @      B@      A@      5@     �L@      "@      I@      @     �C@      �?      J@      2@      &@      &@      1@     �C@      3@      P@      =@     �M@      .@      @              @      @       @      1@       @      "@      �?       @              �?      �?       @      �?      @      @      �?      .@      @      @@      A@      0@     �I@      @     �@@      @      >@              F@      2@      $@      $@      .@      C@      .@      M@      <@      F@      (@     �E@      <@      ;@      G@      ,@      J@      �?      G@      @      I@      <@      "@      @      :@      D@       @     �S@     �R@     �J@      (@      *@      ,@      *@      7@      @      8@              @@       @      5@      (@      @              *@      7@      @      @@     �E@      6@      @      @      @       @      @      �?      @               @      �?       @      @      �?              �?       @      @      @      ,@       @      �?      @      &@      &@      2@       @      5@              8@      �?      *@      @      @              (@      .@       @      =@      =@      4@      @      >@      ,@      ,@      7@      &@      <@      �?      ,@      @      =@      0@      @      @      *@      1@      @     �G@      @@      ?@      @      7@      @      *@      2@      $@      <@      �?      ,@      @      ;@      ,@      @      @      "@      0@      @      G@      7@      :@      @      @      @      �?      @      �?                                       @       @              @      @      �?              �?      "@      @      �?     @h@     �P@      =@      i@      $@     �s@             �\@      @     s@     �D@      ;@      ,@      6@      e@      C@     @l@     �c@     �p@      H@     �a@     �D@      5@     �c@      "@     �o@             �W@      @     �j@      ?@      8@      @      .@      `@      @@      e@     �^@     �j@     �E@      `@      A@      1@     @c@      "@     @m@             �U@      @     @i@      7@      4@      @      .@     @\@      7@     �b@     @Y@     �g@     �E@     �L@      4@      (@     �Y@      �?     �c@             �G@             ``@      (@      0@      @      @      S@      $@     �Y@     �M@     �b@      4@      R@      ,@      @     �I@       @     @S@             �C@      @     �Q@      &@      @      �?      $@     �B@      *@     �G@      E@      D@      7@      (@      @      @      @              2@               @              (@       @      @       @              .@      "@      2@      5@      6@               @      @      �?      @              0@               @              &@      @      @       @              .@       @      0@      3@      &@              @      �?      @                       @                              �?      @                                      �?       @       @      &@             �J@      9@       @      E@      �?     �N@              5@      �?     �V@      $@      @       @      @     �D@      @      M@      B@      M@      @      <@      (@       @      3@             �F@              1@      �?     �D@      @       @      @      �?      =@       @     �@@      6@     �A@       @      &@       @      �?      (@              4@              &@      �?      &@       @                      �?      .@       @      2@       @      $@      �?      1@      $@      �?      @              9@              @              >@      �?       @      @              ,@              .@      ,@      9@      �?      9@      *@      @      7@      �?      0@              @              I@      @      �?      @      @      (@      @      9@      ,@      7@      @      @       @      @      5@      �?      @               @              @@      @                      @      @       @      &@      $@      @       @      4@      @      @       @              (@               @              2@      @      �?      @       @      @       @      ,@      @      2@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJUhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?F7K��m@�	           ��@       	                    �?�ݯ��@�           d�@                           @pӸx�]@W           x�@                          �:@z-+@�            �v@������������������������       ���8C��@�            Pr@������������������������       �\�LU3�@)            �Q@                           @�2e�x�@w            �h@������������������������       �Q�؟�@^            �c@������������������������       �_�8r7@             C@
                          �:@��[���@�           ��@                          �1@�U)(�@           ��@������������������������       ���e@<            �X@������������������������       ���թ��@�           ��@                           �?��n�ae@�             o@������������������������       ��Gv@@'            @P@������������������������       ��Lkv�*@s            �f@                            �?x�܍�+@�           �@                           �?�j���@�           ��@                          �1@>\<�3S@t            �e@������������������������       �ɈsBz�@             C@������������������������       �Y��!�2@[            �`@                           @A�V�@           {@������������������������       ���Ƿ��@�            �s@������������������������       �r�Z
/�@G            �]@                          �3@�O�!@0           H�@                           �?� �O��@�           ��@������������������������       �|���
@�            @t@������������������������       �)�h�U�@�            w@                          �>@MA���@r           �@������������������������       �+�*f�r@T           8�@������������������������       ��qc�&	@             K@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       `u@     �_@      W@      w@      B@      @      .@     �j@     �B@     �}@     �W@      L@      @@      H@     `n@     �O@     �u@     �s@     �{@     @P@      a@     �Q@      O@     �d@      5@     �c@      *@     �X@      8@     �c@      A@      C@      1@      A@     @\@      <@     �b@      `@     �b@      =@     �L@      (@      6@      E@       @      O@      @     �@@      @     �O@      0@      *@      @      &@      F@      @     �D@     �E@      L@      (@      =@      @      &@      3@      @      K@      @      ;@      @      F@      ,@      (@       @      @      5@      @      <@      ;@     �B@      @      ;@      @      @      ,@      @     �I@      @      2@      �?      D@      @      (@              @      0@      @      :@      5@      @@      @       @      �?      @      @              @      @      "@      @      @       @               @      @      @      �?       @      @      @              <@      @      &@      7@      @       @              @      �?      3@       @      �?      @      @      7@              *@      0@      3@      @      *@      @      $@      4@      @      @              @              $@      �?      �?      @      @      6@              (@      ,@      3@      @      .@              �?      @      �?      @                      �?      "@      �?                              �?              �?       @                      T@     �M@      D@     �^@      *@     �W@      @     @P@      2@     �W@      2@      9@      (@      7@     @Q@      5@     �Z@     �U@     �W@      1@      O@     �B@      =@     @V@      &@      U@      @      G@      2@      T@      2@      0@       @      3@      L@      $@      V@      J@     �R@      0@      $@               @      (@              "@      @       @              $@              @                      *@              @      @      ,@              J@     �B@      ;@     @S@      &@     �R@      �?      C@      2@     �Q@      2@      &@       @      3@     �E@      $@      U@     �F@      N@      0@      2@      6@      &@     �@@       @      &@       @      3@              ,@              "@      @      @      *@      &@      3@      A@      5@      �?      @      @              @              @       @      @              @              @                      �?              $@      @      "@              &@      .@      &@      ;@       @      @              ,@              "@              @      @      @      (@      &@      "@      <@      (@      �?     �i@      L@      >@     �i@      .@     Pu@       @     �\@      *@      t@      N@      2@      .@      ,@     @`@     �A@      i@     `g@     0r@      B@      M@      3@      1@     �L@             �W@              6@       @     �R@      1@      @       @      @      C@      @      J@      H@     @S@      "@      1@              @      7@              =@              (@       @      4@      �?                              1@      �?      0@      ,@      (@      @      �?                      @               @                               @                                      @      �?       @      �?      @       @      0@              @      2@              5@              (@       @      (@      �?                              &@              ,@      *@       @       @     �D@      3@      (@      A@             @P@              $@              K@      0@      @       @      @      5@      @      B@      A@     @P@      @      6@      ,@      "@      ?@              D@               @             �E@      (@      @       @      @      2@      @      6@      ?@      D@      @      3@      @      @      @              9@               @              &@      @                      �?      @              ,@      @      9@             `b@     �B@      *@     `b@      .@     �n@       @     @W@      &@     �n@     �E@      .@      @      $@      W@      <@     �b@     `a@     �j@      ;@      @@      $@      @      Q@      @     �Y@             �D@             �_@      $@      @       @      @     �D@      2@      N@     �L@      Z@      @      .@      @       @      ?@      @     �N@              .@             �G@      @      �?               @      1@      �?      >@     �@@      L@       @      1@      @      @     �B@             �D@              :@             �S@      @      @       @      �?      8@      1@      >@      8@      H@      �?     �\@      ;@      @     �S@      &@      b@       @      J@      &@      ^@     �@@      "@      @      @     �I@      $@     @V@     �T@     �[@      8@      [@      :@      @     �S@       @     �a@              J@      &@     �[@     �@@      "@      @      @      I@      "@      S@     �T@     �Y@      7@      @      �?      �?              @      @       @                      $@                               @      �?      �?      *@              @      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �:@}r��n�@�	           ��@       	                   �3@�܁��@/           0�@                           @���!��@[           ��@                          �1@���|!d@P           ��@������������������������       ��w�>�O@           �{@������������������������       ��wĄ��@=           �@                            �?[��լ�@            {@������������������������       ���'L�@�            �p@������������������������       ����@p            �d@
                           �?H�cq �@�           ��@                            @{9�β�@!           ��@������������������������       ��9��M�@A           �@������������������������       �S]�� @�            �u@                           @�1����@�           x�@������������������������       �W�CwK@0           @@������������������������       �����@�           P�@                           @��sƛH@`           ��@                          �<@��t@�             s@                           �?�օ@\            @a@������������������������       ��5TL�@7             U@������������������������       ���Z�f�@%             K@                            @<�Z��@k            �d@������������������������       �Կ����@D             Y@������������������������       ������@'            �P@                           �?�����@�            p@                            �?r�z��g@Z            �b@������������������������       �v����
@             I@������������������������       ������@<            �X@                           @Z��0�@?             [@������������������������       ��F����@             F@������������������������       �%����@%             P@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@     �a@     �T@     Pv@      G@     �@      @     �k@      ;@     �|@     @\@     �K@      E@     �R@     �j@      N@     �u@     @r@     �{@     �T@     �r@     �\@     �M@     �r@      D@     �}@      @      f@      2@     �y@      U@     �G@      7@      M@     �f@     �D@     �s@      n@     �x@     �Q@     @Y@      B@      6@     @`@      &@     �k@      �?     @S@       @      h@     �A@      3@      @      ,@      S@      *@      ]@      X@     `i@      *@     @R@      3@      (@     �T@      &@      b@      �?      J@       @     �b@      3@      .@      @      @     �K@      @     �R@     �L@     �c@      $@      <@       @       @      ?@      $@     @T@      �?      7@      �?      Q@      $@      @      �?      @      <@      @      <@     �@@     �Q@      @     �F@      1@      @      J@      �?     �O@              =@      �?     �T@      "@      $@      @      �?      ;@      �?     �G@      8@     �U@      @      <@      1@      $@     �G@             �S@              9@             �D@      0@      @              "@      5@      @     �D@     �C@      G@      @      ,@      &@      @     �@@             �D@              ,@              ;@      @       @              "@      &@      @      6@      >@      A@       @      ,@      @      @      ,@              C@              &@              ,@      &@       @                      $@       @      3@      "@      (@      �?     �h@     �S@     �B@      e@      =@     �o@       @     �X@      0@     �k@     �H@      <@      3@      F@     �Z@      <@     �h@      b@     @h@     �L@      T@      A@      <@     �L@      5@     @V@       @      E@      *@      U@      8@      1@      @      ?@     �H@      0@      W@     �P@     �R@      6@      K@      8@      ,@      D@      "@      L@       @      2@      @     �J@      $@      "@              *@      ?@       @      J@      @@      N@      *@      :@      $@      ,@      1@      (@     �@@              8@      @      ?@      ,@       @      @      2@      2@       @      D@     �A@      .@      "@     @]@      F@      "@      \@       @     `d@             �L@      @     @a@      9@      &@      (@      *@     �L@      (@     �Z@     @S@     �]@     �A@      G@      1@       @      L@       @     @P@              @@             �R@      (@              @      �?      ;@      @      G@      4@     @Q@      4@     �Q@      ;@      @      L@      @     �X@              9@      @     �O@      *@      &@      @      (@      >@      @      N@     �L@      I@      .@      G@      ;@      7@      M@      @      >@      @      F@      "@      E@      =@       @      3@      1@     �@@      3@      B@      J@      G@      *@      ?@      4@      0@      6@      @      &@      @      6@      @      .@      .@      @      ,@      @      6@      *@      4@      @@      1@      @      &@       @      �?      2@       @      @      @      .@      @       @       @      @      @       @      @      @      $@      4@      (@       @      @      �?      �?      *@       @              @      (@      @      �?      @      @      @      �?      @      @      @      0@      @       @       @      �?              @              @              @       @      �?      @      �?              �?      @              @      @       @              4@      2@      .@      @      @      @      �?      @              *@      @       @      &@      @      .@      "@      $@      (@      @      @      *@      ,@      @       @              @      �?      @              $@      @              &@      @      $@      @      @      @      �?              @      @      "@       @      @                      @              @       @       @              �?      @      @      @      @      @      @      .@      @      @      B@      �?      3@              6@      @      ;@      ,@       @      @      &@      &@      @      0@      4@      =@      @      @      @      @      <@              @              0@              ,@      @       @       @      @       @      @      @      &@      6@       @              �?      @       @              �?              @                       @               @      @               @       @      "@       @      �?      @      @      �?      4@              @              &@              ,@      @       @               @       @      �?      @       @      ,@      �?      "@               @       @      �?      ,@              @      @      *@      "@              @      @      @      @      $@      "@      @      @      �?                                      ,@                      @      @      @              @      �?      �?      �?       @      @      @               @               @       @      �?                      @               @      @                      @       @       @       @      @       @      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJW>=khG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@b9PG��@�	           ��@       	                     �?I�n���@v           ؕ@                           �?����r?@�           p�@                          �2@���@�            �r@������������������������       ��z!��
@�            @l@������������������������       �/�E ��@0            �R@                           @�TQ�d@9           ~@������������������������       ��tǩH@�            �p@������������������������       �7���v�
@�            `j@
                           @s5�T�@~           @�@                           @m�o��U@           �z@������������������������       �t��ԉ@�            Pr@������������������������       �_�Q��
@U             a@                           @޿�0�J	@h            `g@������������������������       ��MZk��@J            �_@������������������������       ������@             N@                           �?}�(l.�@I           ��@                           @Q��(@@�           $�@                           �?j��t�,@           @�@������������������������       ��ȬR@�            �o@������������������������       ��M��d4@`           P�@                           @)S�o��@�            v@������������������������       �R��@            �A@������������������������       �!�jG��@�            �s@                           @o�x5�@X           (�@                          �5@Ϟ<Qp:@           P�@������������������������       �:ݟ#�@�            �r@������������������������       ��3?��@H            �@                           @W-��@U            �@������������������������       �m�8�@_            @c@������������������������       � jͭC@�            `x@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �`@     �\@     �w@     �D@     0~@      @      n@      A@     `z@     @[@     �Q@      A@     �O@     �l@     �F@      v@     �q@     �{@     �X@     �W@      =@      <@     �b@      @      k@             @S@      @      f@      =@      8@      @      @     �S@      @     �_@     �Z@      j@      9@      G@      6@      $@     �Y@              Z@             �D@      @     �[@      0@      &@      @      @      A@       @     @P@      M@      `@      1@      :@      @      @      E@             �G@              5@       @      I@      "@       @               @      ,@              *@      .@     �G@       @      1@       @      @      =@              @@              4@      �?     �C@      @                       @      @              *@      ,@     �B@       @      "@      �?              *@              .@              �?      �?      &@      @       @                       @                      �?      $@              4@      3@      @     �N@             �L@              4@      @     �N@      @      "@      @       @      4@       @      J@     �E@     �T@      .@      "@       @      @      G@              7@              $@      @      <@      @      @      �?       @      1@      �?      A@      9@      E@      &@      &@      1@      �?      .@              A@              $@             �@@      �?       @      @              @      �?      2@      2@      D@      @      H@      @      2@      H@      @     @\@              B@             �P@      *@      *@      @       @      F@       @      O@      H@     �S@       @      D@      @      *@      B@      @     �Q@              ;@             �B@      *@      (@      @      �?      7@       @      F@     �C@      I@      @      <@      @      *@      0@      @     �C@              1@              8@       @      "@      �?      �?      3@              B@      <@      B@      @      (@                      4@      �?      ?@              $@              *@      @      @       @              @       @       @      &@      ,@               @              @      (@             �E@              "@              =@              �?              �?      5@              2@      "@      =@       @      @              @       @              >@              "@              9@              �?              �?       @              ,@      "@      1@       @      @                      @              *@                              @                                      3@              @              (@             `m@     �Z@     �U@      l@     �A@     �p@      @     `d@      =@     �n@      T@     �G@      ;@     �L@      c@     �D@      l@     @f@     �m@     @R@      Z@     �N@     �I@     �W@      8@     @V@      @     �V@      4@     �Y@      C@      9@      .@      C@      M@      ;@      Z@     �Q@     �Y@      E@     @S@      B@     �B@     �R@      ,@     �Q@      @      M@      ,@     @P@     �A@      1@       @      5@      ?@      3@     �R@      L@     �O@      ?@      =@       @      &@      .@       @      7@       @      2@      @      7@      $@      �?      @      @      &@       @      ;@      1@      ?@      @      H@      <@      :@      N@      @      H@      @      D@      $@      E@      9@      0@      @      0@      4@      1@      H@     �C@      @@      :@      ;@      9@      ,@      3@      $@      2@              @@      @      C@      @       @      @      1@      ;@       @      =@      .@     �C@      &@               @              �?                               @                                              @       @      �?      @       @      @      @      ;@      7@      ,@      2@      $@      2@              8@      @      C@      @       @      @      *@      9@      @      :@      *@      A@      @     ``@     �F@     �A@     ``@      &@      f@       @     @R@      "@     �a@      E@      6@      (@      3@     �W@      ,@     @^@     �Z@     �`@      ?@     �R@      ;@      ,@     �R@      @      ^@             �I@              X@      6@      @      @      @      N@      @     �S@      M@     �U@      4@      *@      .@      @      >@             �I@              2@              7@      @      @      @      �?      3@       @      B@      :@      C@      $@      O@      (@      "@     �F@      @     @Q@             �@@             @R@      2@      �?       @      @     �D@      �?     �E@      @@     �H@      $@      L@      2@      5@      L@      @     �L@       @      6@      "@      G@      4@      1@      @      *@     �A@      &@      E@     �H@      H@      &@      *@       @      @      3@      @      .@              $@      �?      (@      &@      @       @              *@      "@      .@      $@      @      @     �E@      0@      0@     �B@      �?      E@       @      (@       @      A@      "@      &@      @      *@      6@       @      ;@     �C@     �E@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJbhhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�k;�y�@�	           ��@       	                     @[��#��@�           ��@                          �3@�5�@8           H�@                           �?VUwRk@r           ��@������������������������       �>���_
@�            �x@������������������������       ����֦�@�           8�@                           �?�=���@�           ��@������������������������       �F��@�            Pq@������������������������       ����>	3@$           �|@
                           @·I�,C@�           ��@                           �?�+P��@�            �r@������������������������       ���]il@d            `c@������������������������       ��I�ϣ�
@`            �b@                          �4@��!�B@�             t@������������������������       ��b��?v@�             m@������������������������       �WC[��
@8            @V@                           @��2~r�@�           �@                           �?�?S3
@�           ��@                            @%߂�^@
           �z@������������������������       �Bi �/@�            �r@������������������������       ��Ξ���@M            ``@                            @��$ؙ@�           ��@������������������������       � ?�@F@.           �}@������������������������       �&G1��D@�             l@                           @X)-=�@           �y@                          �;@Bk6y@�            �w@������������������������       �zV�'G@�            �p@������������������������       �nEhB��@K            @\@                          �9@�����	@             @@������������������������       �m�u5x@             4@������������������������       �B8iY�o @             (@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �c@     @X@     �v@     �D@     �}@      "@     �m@      =@     0z@     �`@      N@      <@      P@      k@     �L@     x@     Ps@     @z@      U@     `d@     �P@      I@     �n@      2@     Pv@      �?     �a@      &@     Pq@      P@     �D@      "@      2@     @[@      8@     �o@     �h@     @q@     �F@     �]@     �G@      >@      i@      @      q@             @U@      $@     �j@      A@      >@       @      $@     @T@      4@     �g@     @a@     �k@      A@     �N@      6@      2@      _@      @     �c@              I@             �b@      (@      3@      @      @      E@      @     �X@     �S@     �a@      1@      7@      @      @     �K@             �P@              8@             �S@      �?      @              �?      3@      �?     �@@      6@     �I@       @      C@      1@      (@     @Q@      @      W@              :@              R@      &@      0@      @      @      7@      @     �P@      L@     �V@      "@     �L@      9@      (@      S@      @     �\@             �A@      $@      P@      6@      &@      @      @     �C@      ,@     �V@      N@     �S@      1@      7@      &@      @      7@             �F@              &@              ,@       @      �?              @      .@              E@      >@      B@      "@      A@      ,@      @     �J@      @     @Q@              8@      $@      I@      ,@      $@      @       @      8@      ,@      H@      >@      E@       @     �F@      3@      4@     �G@      (@     @U@      �?     �L@      �?     �O@      >@      &@      �?       @      <@      @     @P@     �N@      L@      &@      ;@      @      &@      0@      @      H@             �E@      �?      6@      @       @              @      &@      �?      =@      =@      A@      @      (@      @      $@              @      1@              8@      �?      (@       @       @              @      @      �?      0@      2@      4@              .@      @      �?      0@              ?@              3@              $@      @                              @              *@      &@      ,@      @      2@      *@      "@      ?@      "@     �B@      �?      ,@             �D@      8@      "@      �?      �?      1@      @      B@      @@      6@      @      (@       @      @      ;@      "@      7@      �?      "@              9@      .@      @      �?      �?      .@      @      8@      8@      6@      @      @      @       @      @              ,@              @              0@      "@      @                       @              (@       @                     �d@      W@     �G@     @\@      7@      ^@       @     @X@      2@     �a@      Q@      3@      3@      G@      [@     �@@     ``@     �[@      b@     �C@      Z@     @Q@     �A@     �V@      &@      Y@       @     @P@      0@      Z@      M@      3@      .@      <@     @T@      1@     �X@     �T@     @W@      B@     �@@      *@      1@      9@      �?      C@       @      8@      @      G@      7@      @      @       @      D@      $@      F@      E@      ?@      0@      :@      @      (@      1@      �?     �B@              *@              ?@      (@      @      @              >@      @      ?@      ?@      7@      $@      @      @      @       @              �?       @      &@      @      .@      &@       @               @      $@      @      *@      &@       @      @     �Q@      L@      2@     �P@      $@      O@      @     �D@      "@      M@     �A@      *@       @      :@     �D@      @      K@      D@      O@      4@     �G@     �F@      "@      H@      @     �H@      @      ;@      @     �I@      8@       @      @      ,@      <@      @      @@      5@     �E@      (@      8@      &@      "@      2@      @      *@       @      ,@      @      @      &@      @      @      (@      *@      �?      6@      3@      3@       @     �N@      7@      (@      6@      (@      4@              @@       @      C@      $@              @      2@      ;@      0@     �@@      <@     �I@      @      N@      4@      (@      5@       @      4@              @@       @     �A@      @              @      2@      :@      .@      <@      7@      G@      @     �J@      *@      $@      *@      @      1@              *@       @      6@      @                      *@      5@      (@      2@      "@     �C@              @      @       @       @      �?      @              3@              *@       @              @      @      @      @      $@      ,@      @      @      �?      @              �?      @                                      @      @                              �?      �?      @      @      @              �?      @                      @                                      @                                      �?      �?      @      @                                              �?                                                      @                                               @      �?      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�ªhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�3Jk��@�	           ��@       	                    @��UX@U           ��@                            �?T��6�@           `�@                           �?�nc�H@           |@������������������������       �~�;]u@k            �e@������������������������       �:�*o�@�            @q@                           �?"�dd�(@�            �v@������������������������       �����}(@�            �p@������������������������       ��=���@>             W@
                           @�sH�
�@G           ��@                           @<jv�lH@w            �f@������������������������       �c�}K�`
@R            �_@������������������������       �5�_��@%             K@                           �?BUn*@�           ��@������������������������       ��@e��C
@�            @r@������������������������       �겘�@           �{@                            @�@����@b           �@                           @_�҅��@�           ܗ@                            �?��We"P@2           (�@������������������������       �1��Ē@�            �u@������������������������       ��]鹌�@_           H�@                           @h|�J�@�           ��@������������������������       �?i�R֝@            z@������������������������       ��n��o@�             j@                          �;@�ޕ:�=@�           ��@                          �:@���	@K           Ȁ@������������������������       �]b�O�@&           �}@������������������������       ����s.i
@%            �O@                           @-��d0a@T            �^@������������������������       ��rF@L            @[@������������������������       �[�����?             ,@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       pt@     �a@     �S@     0u@      I@     ~@       @     �n@      @@     @}@     �Z@     �P@     �B@     �O@     �k@     @P@     0w@     �r@     �z@     �T@     �_@      D@      9@     �b@      0@     �p@       @     �W@      "@     �k@      C@      >@      (@      ,@      W@      :@     �d@     �a@     �m@      4@      M@      2@      2@     �V@      ,@      Z@       @      F@      @     �S@      =@      *@      @      &@      D@      4@     �S@     �S@     @V@      *@      ;@       @      @     �O@              P@              5@      @     �G@      (@      &@      �?      @      5@      &@     �E@     �@@     �N@      &@      $@      @      �?      .@              A@              *@              4@      @       @      �?               @      �?      3@      (@      :@      @      1@      @      @      H@              >@               @      @      ;@      "@      "@              @      *@      $@      8@      5@     �A@       @      ?@      $@      (@      <@      ,@      D@       @      7@      @      ?@      1@       @      @      @      3@      "@     �A@      G@      <@       @      :@      @      &@      1@      *@      =@       @      2@      @      4@      &@       @      @      @      ,@       @      8@     �A@      9@      �?      @      @      �?      &@      �?      &@              @              &@      @                              @      @      &@      &@      @      �?      Q@      6@      @      M@       @     �d@             �I@       @     �a@      "@      1@      @      @      J@      @     �U@     �O@     �b@      @      @      @              0@              9@              @             �@@      @       @                      $@       @      0@       @     �@@      @      @      @              &@              8@               @              9@      �?      @                      "@      �?      0@      @      ,@      @      @       @              @              �?              @               @      @      @                      �?      �?              @      3@             �N@      0@      @      E@       @     �a@              G@       @     @[@      @      "@      @      @      E@      @     �Q@     �K@     �\@              =@              @      ,@       @     �M@              :@      �?      B@      @                      @      1@      �?      8@      9@      H@              @@      0@      @      <@             @T@              4@      �?     @R@       @      "@      @              9@      @      G@      >@     �P@              i@     �Y@     �J@     �g@      A@     �j@      @     �b@      7@      o@      Q@      B@      9@     �H@     @`@     �C@     �i@     �c@      h@     �O@     �a@     @Q@      =@     �a@      3@     �d@      @      V@      "@      h@      F@      0@      1@      9@     �X@      ?@     @b@     @[@      b@     �B@     �W@      B@      6@     �P@      @     @]@      �?     �K@      @      ^@     �@@      &@      $@      $@     �I@      "@      V@      L@     �T@      =@     �C@      1@      .@      @@       @     �C@      �?      =@      @      E@      0@       @      @      @      3@       @      6@      .@     �A@      "@      L@      3@      @     �A@      @     �S@              :@      �?     �S@      1@      "@      @      @      @@      @     �P@     �D@     �G@      4@      H@     �@@      @     �R@      ,@      H@      @     �@@      @      R@      &@      @      @      .@     �G@      6@      M@     �J@     �O@       @      4@      =@      @      H@      @      :@              ;@      @     �L@       @      @      @      @      B@      2@      D@      ;@      F@       @      <@      @       @      :@      "@      6@      @      @       @      .@      @                      $@      &@      @      2@      :@      3@              M@     �@@      8@     �H@      .@     �G@       @     �N@      ,@      L@      8@      4@       @      8@      @@       @     �N@      I@      H@      :@      F@      2@      4@      B@       @      G@       @      L@      (@     �G@      4@      3@      @      2@      6@      @     �L@     �E@      B@      7@     �D@      2@      3@      <@       @      C@              F@      &@      G@      2@      &@      @      2@      4@      @      L@      D@      9@      7@      @              �?       @               @       @      (@      �?      �?       @       @                       @              �?      @      &@              ,@      .@      @      *@      @      �?              @       @      "@      @      �?      @      @      $@      @      @      @      (@      @      ,@      .@      @      &@      @      �?              @       @      "@      @      �?      @      @       @      @      @      @      $@      @                               @                                                      �?                               @              �?               @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJl8�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��k6G�@�	           ��@       	                   �:@�\�ɔ�@           ,�@                            �?h^pD`�@1           ��@                           �?-����Y@�           ��@������������������������       �7���.�@�            �r@������������������������       ��"n���@�            pw@                            @$�n9+@�           H�@������������������������       ���}"�@B            �Z@������������������������       �
��]m@M           ��@
                           �?BW:%v@�            0v@                          �=@�і��Q@7            �T@������������������������       �S�j��@$             I@������������������������       ����@            �@@                            �?Ke�P�V@�             q@������������������������       �j �iخ@1            @R@������������������������       �	=h�@~            �h@                           �?�X]@�           |�@                           @���4C�@�           ��@                            �?�s��s@�           �@������������������������       ����@G�
@~            @h@������������������������       �|�^�d @I           �@                            �?{0�=�m@�            x@������������������������       ������@�             l@������������������������       �TlM{�@i             d@                           @8����@�            �@                           @�B4'@�           ��@������������������������       ������@T           ��@������������������������       �����/�@j            �c@                          �4@>�c�@+            }@������������������������       �yk\��L@�            @n@������������������������       �P*�zB@�            �k@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       Ps@     `b@     �Y@     �v@      >@     �|@      @      k@      @@     �~@     �[@     �P@      =@     �P@     �k@      R@     v@     `s@     �{@     �T@     �`@     @S@     �S@     @c@      4@     @a@      @      Y@      8@     �e@      J@      B@      1@     �E@     �Y@      <@      a@     �a@     `e@     �D@     @[@      J@      L@     @^@      .@     �`@      @      P@      6@     @b@      E@      =@      @     �B@     @U@      0@      \@     @Z@     @`@     �B@     �F@      :@      ?@     �S@      @     @P@      @      >@      (@     @S@      .@      8@      @      0@     �G@      &@      L@     �A@     �R@      ,@      8@      (@      4@      ?@              A@       @      $@       @      >@      &@      @      @      @      1@      "@      6@      (@     �C@      @      5@      ,@      &@      H@      @      ?@      �?      4@      $@     �G@      @      4@              "@      >@       @      A@      7@      B@      @      P@      :@      9@      E@       @     �P@              A@      $@     @Q@      ;@      @      @      5@      C@      @      L@     �Q@     �K@      7@      $@      @              "@       @      ,@              @              4@       @                      �?      @              @      &@      ,@      @      K@      5@      9@     �@@      @     �J@              ?@      $@     �H@      9@      @      @      4@      A@      @     �I@     �M@     �D@      0@      8@      9@      7@     �@@      @      @       @      B@       @      <@      $@      @      $@      @      2@      (@      9@      C@     �D@      @      @      �?      @      @              @      �?       @              &@      �?      �?      @      �?       @      �?      &@      @      ,@       @       @      �?      @                       @      �?      @              @      �?      �?      @              �?              @      @      &@       @       @                      @               @               @              @                              �?      �?      �?      @       @      @              4@      8@      2@      ;@      @       @      �?      <@       @      1@      "@      @      @      @      0@      &@      ,@      ?@      ;@       @      �?      @       @      "@      �?      �?              $@              @      �?              @      @      @       @      @      @      $@       @      3@      5@      0@      2@      @      �?      �?      2@       @      $@       @      @       @       @      &@      "@      $@      8@      1@              f@     �Q@      8@      j@      $@     0t@             @]@       @     t@     �M@      >@      (@      7@     @]@      F@      k@     �d@     �p@      E@     �T@      ;@      $@     @Z@       @      c@             �N@      @      f@      8@      (@      @      @     �E@      2@      X@     �S@     �b@      ;@     �H@      1@      @      K@      @      Y@             �I@      @      a@      0@       @      @      @      8@      @     �N@     �A@      [@      4@      *@      @              .@      �?      @@              .@              F@              �?      @              @      �?      9@      @      0@      @      B@      $@      @     �C@      @      Q@              B@      @      W@      0@      �?      @      @      1@      @      B@      <@      W@      *@     �@@      $@      @     �I@      @      J@              $@      �?      D@       @      $@      �?       @      3@      ,@     �A@     �E@      D@      @      8@      @      @      @@       @      7@              @              6@       @              �?      �?      .@       @      6@      >@      5@      @      "@      @      @      3@      �?      =@              @      �?      2@              $@              �?      @      @      *@      *@      3@      @     �W@     �E@      ,@      Z@       @     `e@              L@      @      b@     �A@      2@      @      0@     �R@      :@      ^@     @V@     �^@      .@      H@      7@      "@      S@       @     �[@              @@      �?      V@      6@      $@      @      @      E@      7@     �R@      L@     �M@      @      D@      3@      "@     �N@       @     �S@              *@             @R@      ,@      @       @      @      B@      2@     �N@      C@     �I@      @       @      @              .@              @@              3@      �?      .@       @      @      �?              @      @      *@      2@       @              G@      4@      @      <@              N@              8@       @     �L@      *@       @       @      (@      @@      @      G@     �@@     �O@      $@      2@      @      @      *@             �F@              1@       @     �C@      @      @      �?              ,@       @      6@      ,@      =@       @      <@      *@       @      .@              .@              @              2@      $@      @      �?      (@      2@      �?      8@      3@      A@       @�t�bub��     hhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ|��OhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@oҫ�u�@�	           ��@       	                    �?o~9��@+           \�@                          �2@#17y��@a           �@                          �1@���g�@R           ��@������������������������       �+R��ƺ@�            �t@������������������������       �j!�Ñ�
@|            @i@                          �3@��x��@           �z@������������������������       ��ˎj�	@_            �b@������������������������       �h�k
J?@�            `q@
                            @}��@�           ��@                           @�{�&�@           ��@������������������������       �����@           `y@������������������������       ��Zd��E@            |@                          �2@Ђ8��@�            `q@������������������������       ��S/��@W            @a@������������������������       �ڞ�ۋO@Z            �a@                           �?�:��@�           l�@                            �?�i{w@�            �s@                            �?��U��@r            @i@������������������������       ��vV���@5            �V@������������������������       �u1f�	@=             \@                            @ȮcM�@F            @\@������������������������       ��G �]@             :@������������������������       ��{Ab3@5            �U@                           �?�.��@�           ��@                          �9@.3�|$�@?           �~@������������������������       ��D\�0@�            �r@������������������������       ����K�@~             h@                           @$�@��@�           ��@������������������������       �8g����@�           Ђ@������������������������       ��>�@           �y@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@      `@     �U@     �v@     �F@     P@      $@      n@      >@     �{@     �W@      J@      D@     �O@     �m@     �Q@     @v@     �r@     �{@     �S@      d@     �K@      6@     @k@      ,@     Pt@      @     ``@      @     `p@      A@      8@      &@      .@     �^@      >@     `h@     �d@     �p@     �@@     �T@      3@      @     @T@      @     �e@             @Q@             `a@      &@      "@       @      @      I@      @      S@      R@     �`@      1@      C@      ,@      @      J@      @      T@              H@              W@      @      �?       @      @      ;@       @     �A@     �E@     �R@      $@      7@      @      @      8@      @     �I@             �A@              L@      @      �?               @      .@       @      6@      >@     �G@      @      .@       @              <@              =@              *@              B@                       @      �?      (@              *@      *@      ;@      @      F@      @      @      =@             �W@              5@             �G@      @       @      @      �?      7@      @     �D@      =@      M@      @      *@       @      �?      "@              C@              @              3@      @       @                      "@      �?      ,@      @      <@       @      ?@      @      @      4@              L@              2@              <@      @      @      @      �?      ,@      @      ;@      8@      >@      @     �S@      B@      .@      a@       @     �b@      @      O@      @     �^@      7@      .@      @      &@      R@      8@     �]@      W@      a@      0@     �O@      8@      &@      ]@       @     �[@              E@      @      X@      2@      $@      @      @      L@      ,@      W@     �N@     @\@      ,@      =@      @      @      M@       @     �L@              3@      @      I@      �?      @       @             �@@      @      H@      8@     �I@      @      A@      1@      @      M@             �J@              7@       @      G@      1@      @      �?      @      7@       @      F@     �B@      O@      $@      0@      (@      @      5@      @     �D@      @      4@       @      ;@      @      @              @      0@      $@      ;@      ?@      7@       @       @       @       @      "@              3@      @      "@              4@               @              �?      &@       @       @      3@      $@      �?       @      @       @      (@      @      6@              &@       @      @      @      @              @      @       @      3@      (@      *@      �?     �d@     @R@      P@     `b@      ?@      f@      @     @[@      7@      g@      N@      <@      =@      H@     @]@      D@      d@     �`@     �e@     �F@      4@      ,@      4@      B@      �?      B@      @      7@      @      6@      @      "@      @      @      <@      "@      1@      3@      A@      @      *@      &@      *@      9@              6@               @              *@      @      @      @       @      4@       @      "@      .@      9@      @      @      @      @      $@              $@              @              @       @               @       @      @      @      @       @      .@       @      "@      @       @      .@              (@              �?              "@       @      @      @              *@      @      @      @      $@      @      @      @      @      &@      �?      ,@      @      .@      @      "@      �?      @              �?       @      �?       @      @      "@      �?      @                                      @              @              @               @                                               @      @              @      @      @      &@      �?      "@      @       @      @      @      �?      @              �?       @      �?       @       @      @      �?     `b@     �M@      F@     �[@      >@     �a@      @     �U@      2@     `d@     �K@      3@      8@     �F@     @V@      ?@      b@     �\@     �a@     �C@      :@      0@      0@     �@@       @      L@              @@      @      O@      0@      @      @      *@      C@      "@      H@      E@      G@      5@      3@      "@      "@      4@              C@              7@              G@      &@              �?      $@      <@      �?      :@      ;@      6@      @      @      @      @      *@       @      2@              "@      @      0@      @      @       @      @      $@       @      6@      .@      8@      ,@     @^@     �E@      <@     �S@      <@      U@      @      K@      ,@     @Y@     �C@      (@      5@      @@     �I@      6@      X@     @R@     �W@      2@     �Q@      8@      5@      H@      ,@      M@      @      =@      $@      G@      A@       @      ,@      7@      >@      "@     �L@      E@      L@      @     �I@      3@      @      >@      ,@      :@              9@      @     �K@      @      @      @      "@      5@      *@     �C@      ?@     �C@      *@�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�^�YhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��K��@�	           ��@       	                   �:@='ΫH�@           x�@                           �?5by���@3           �@                           @r���Ѣ@0           @@������������������������       �܈���@�            �n@������������������������       �jg]2@�            �o@                            @�E�!��@           p�@������������������������       ����ǵ@/           �~@������������������������       ��>§�@�            `v@
                          �;@��uο�@�            �u@                            �?Gª�Δ@3            �T@������������������������       ��Ȓ��@            �A@������������������������       ���@-�g@             H@                           �?cZ!�F�@�            �p@������������������������       ���'�s@)            @Q@������������������������       �?���|@�            �h@                          �6@�����@t           V�@                           @C���@�           ��@                           �?Uȍ-@�           ��@������������������������       �;�¢��
@�            �k@������������������������       �+����@�            py@                           �?�=.��f@5           H�@������������������������       ������@�            @t@������������������������       �����x@i           (�@                           �?g����@�           `�@                           �?�c��u�@�             k@������������������������       �g����@S            �^@������������������������       � � �2
@A            �W@                           �?c,	7#7@)           0}@������������������������       ��N湬=@�            �j@������������������������       �H��]
�@�            �o@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �`@     �U@     �t@     �C@     �@       @     �n@     �C@     p{@     @Y@      R@      G@     �R@     `m@     @T@     �v@     �p@     �z@     @T@     �a@     @Q@      J@     @b@      8@      e@       @     �]@      :@     �b@      H@     �H@      6@      F@     �Y@      A@     @c@      ^@      f@     �E@     �[@     �D@      C@     @\@      7@     �b@      @     @U@      9@     @`@      C@      C@      "@      B@     �U@      4@     @`@     @W@      a@     �C@      K@      (@      0@      E@      @     �I@       @     �@@      �?      G@      (@      ,@      @      @     �D@      @      F@     �B@     �O@       @      6@      @      @      2@              9@       @      9@              9@      @       @      @      @      0@      @      5@      1@      C@      @      @@       @      *@      8@      @      :@               @      �?      5@       @      @               @      9@      �?      7@      4@      9@      @      L@      =@      6@     �Q@      0@      Y@      �?      J@      8@      U@      :@      8@      @      =@      G@      .@     �U@      L@     �R@      ?@     �A@      0@      0@      H@       @     �K@      �?      3@      1@      K@      ,@      ,@      �?      ,@      <@      .@      C@      6@      L@      1@      5@      *@      @      7@       @     �F@             �@@      @      >@      (@      $@      @      .@      2@              H@      A@      2@      ,@      >@      <@      ,@     �@@      �?      1@      @      A@      �?      3@      $@      &@      *@       @      .@      ,@      8@      ;@      D@      @      �?               @      *@              @      @      $@               @              @      �?              @      @      @      *@      ,@      �?                              @              @              @                                      �?                       @       @      @       @      �?      �?               @       @              �?      @      @               @              @                      @      @      �?      @      @              =@      <@      (@      4@      �?      (@      �?      8@      �?      1@      $@      @      (@       @      (@      "@      5@      ,@      :@      @      $@      @       @      @              $@              @      �?      @               @       @       @      @              @      �?      $@              3@      5@      $@      1@      �?       @      �?      4@              (@      $@      @      $@      @      "@      "@      ,@      *@      0@      @      h@     �P@      A@     `g@      .@      u@             @_@      *@      r@     �J@      7@      8@      >@     �`@     �G@      j@     �b@     �o@      C@     �Y@      A@      9@     �a@      @     Pq@             @X@      @     �h@      ;@      .@      ,@      *@     �U@      A@     �a@      Y@     �h@      2@     �D@      0@      (@     @Q@      �?     �W@              A@             �V@      ,@      @      @      @     �C@      ;@      R@     �C@      M@      @      ,@      @       @      6@              F@              *@              @@       @                       @      0@      �?      ;@      ,@      9@      @      ;@      *@      $@     �G@      �?     �I@              5@              M@      (@      @      @      @      7@      :@     �F@      9@     �@@      �?      O@      2@      *@     �R@      @     �f@             �O@      @     �Z@      *@      (@       @      @      H@      @     �Q@     �N@     `a@      &@      <@      @      @     �@@      @     �Q@              <@      �?      6@      @                      @      5@       @      (@      9@     �L@      �?      A@      (@      "@     �D@             �[@             �A@      @      U@      "@      (@       @      @      ;@      @      M@      B@     �T@      $@     @V@      @@      "@      F@       @     �M@              <@      @     �W@      :@       @      $@      1@      G@      *@     �P@     �I@     �L@      4@      ;@       @      @      "@       @      3@              &@              B@      @      @              �?      2@       @      <@      4@      3@       @      (@              @      "@       @      @              "@              7@      @       @              �?      "@      �?      (@      &@      $@       @      .@       @      �?                      (@               @              *@      @       @                      "@      �?      0@      "@      "@              O@      >@      @     �A@      @      D@              1@      @      M@      3@      @      $@      0@      <@      &@      C@      ?@      C@      (@      >@      *@              1@      @      8@               @      @      >@      "@       @      �?      �?      *@      @      "@      0@      ,@      @      @@      1@      @      2@              0@              "@              <@      $@       @      "@      .@      .@      @      =@      .@      8@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJߦjxhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�Ju.�@�	           ��@       	                     @P^n�z@�           �@                          �2@:JD�@X           �@                           �?��o��@�           ��@������������������������       �w���@j            �f@������������������������       �r��,�@           ��@                            �?�d���n@o           ��@������������������������       ��Ҿ�@�           ��@������������������������       �qXVKB�
@�            @p@
                           �?�yL�rZ@�           ��@                           @��Al�@�            `s@������������������������       �	�z0H�@\            ``@������������������������       ���c�H�@d            `f@                           @α~�!�@�            �t@������������������������       ���G��@�            Pr@������������������������       �oXi<}�@             B@                           �?V��:�@�           �@                           �?6V��@k           P�@                           �?�#�ׅ@�            �l@������������������������       �t��^�	@'             K@������������������������       ����7@u            �e@                          �7@܆u��@�            Pt@������������������������       �	�R�@(            @P@������������������������       �R�"�3@�            @p@                            @Q�a���@B           Ȍ@                           �?Pb�-�Q@r           ��@������������������������       ��7�g��@�            �r@������������������������       ���ƀK@�            r@                           @��2@�            �t@������������������������       ���1��@�             r@������������������������       ���0j@            �C@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        u@     �`@     �V@     �u@      C@     }@       @     @n@      :@     0@     @Z@      L@      B@     �P@      k@     �P@      v@     @s@      {@     @V@     @h@      N@      H@     �k@      1@     �v@      �?     �a@      $@     �u@     �M@      =@      &@     �@@      `@      =@     `l@      f@     �q@     �J@     ``@     �D@      >@     `f@      @     �p@             �Y@      @     �p@      @@      8@       @      0@     @Y@      3@     �d@     �_@     �l@      F@     �G@      (@       @      R@      @      \@              N@      �?     @a@      &@      @      @      $@     �@@      @     �J@     �N@     `a@      @      *@       @      @      7@       @      .@              &@      �?      8@       @      �?      @      @      $@      �?      @      .@      E@      �?      A@      $@      @     �H@      �?     @X@             �H@             �\@      "@      @      �?      @      7@      @     �H@      G@     @X@      @      U@      =@      6@     �Z@       @     �c@              E@      @     �`@      5@      2@      @      @      Q@      (@      \@     @P@     �V@     �B@     �Q@      ;@      5@      T@       @     �Y@              A@      @      X@      3@      ,@      @      @     �I@      (@     �P@      I@      R@      :@      ,@       @      �?      ;@             �J@               @      @     �B@       @      @               @      1@             �F@      .@      3@      &@     �O@      3@      2@     �E@      (@     �X@      �?      C@      @     @S@      ;@      @      @      1@      <@      $@      O@      I@      L@      "@      E@       @      &@      6@      @     �F@              .@             �C@      .@               @      @      *@      @      ;@      9@      A@      @      *@      �?      @      (@      @      9@              "@              @      "@               @      @      @              ,@      @      2@       @      =@      �?       @      $@      @      4@              @              @@      @                               @      @      *@      4@      0@      @      5@      1@      @      5@      @     �J@      �?      7@      @      C@      (@      @      �?      ,@      .@      @     �A@      9@      6@      @      4@      1@      @      1@      @      H@      �?      3@      @      ;@      (@      @      �?      $@      &@      @      A@      9@      4@      @      �?                      @              @              @              &@                              @      @              �?               @             �a@     �R@     �E@      `@      5@     �X@      �?     �Y@      0@     �b@      G@      ;@      9@     �@@      V@      C@     @_@     �`@     @b@      B@     �P@      &@      ,@     �G@      $@     �B@              C@      &@     @R@      0@      @      @      @     �D@      @     �I@     �E@     �L@      ,@      0@       @      *@      (@      @      "@              2@      @      <@      @      �?      @      @      0@       @      >@      3@      ?@      @       @              @       @              �?              @              &@      �?                              @              @       @      (@      �?      ,@       @      "@      $@      @       @              .@      @      1@      @      �?      @      @      &@       @      :@      &@      3@      @     �I@      "@      �?     �A@      @      <@              4@      @     �F@      "@      @       @      @      9@      @      5@      8@      :@      "@      0@                      ,@              @                       @      @       @                              @               @      *@      @             �A@      "@      �?      5@      @      8@              4@      @     �C@      @      @       @      @      6@      @      3@      &@      7@      "@     �R@      P@      =@     �T@      &@      O@      �?      P@      @     �S@      >@      7@      2@      ;@     �G@      ?@     �R@     @V@     @V@      6@     �I@      I@      .@     �J@      @      A@      �?      ?@              N@      2@      *@      $@      0@      ?@      6@      J@     �J@     �P@      $@      3@      =@       @      @@      @      &@      �?      5@              >@       @      "@      @      &@      $@      &@      ;@      9@      @@      @      @@      5@      @      5@              7@              $@              >@      $@      @      @      @      5@      &@      9@      <@      A@      @      8@      ,@      ,@      =@      @      <@             �@@      @      2@      (@      $@       @      &@      0@      "@      6@      B@      7@      (@      4@      $@      ,@      8@      @      <@             �@@      @      (@      @      $@      @      $@      *@       @      6@     �A@      3@      $@      @      @              @                                              @      @              @      �?      @      �?              �?      @       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJʡm`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�ک�@�	           ��@       	                    �?C��u�T@t            �@                            �?6-á�+@�           p�@                           @����=@�             x@������������������������       ��! ��
@�            `t@������������������������       �s�k9<�	@&             N@                           @��ښU�@�            �p@������������������������       ����@O            �\@������������������������       ��sm��	@f            @c@
                            @��2���@�           ȑ@                           @C9?�e(@           �@������������������������       �_�Z�@p            @f@������������������������       ���P�}�@�           ��@                           @P��7UU@�             s@������������������������       �н���@}            `g@������������������������       � g�.m@D            @]@                          �:@ˆ7 AN@8           ��@                           @��g���@�           ��@                          �7@06���-@6           ��@������������������������       ��@~{F�@G            �@������������������������       �bn #��@�            �w@                            �?~p��@�           �@������������������������       ��lH�d@z            �f@������������������������       ���M�@           �|@                          �@@�H�!@m           X�@                           �?�\
��	@D           8�@������������������������       �=�:��@            `i@������������������������       ��ׄ`�T@�            �s@                           @%��pe�@)             Q@������������������������       �,sZ��@             2@������������������������       �k�F�R	@             I@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@     `a@     @Y@     �t@      B@     �~@      @      i@      ?@      }@     �Y@      L@      <@     �Q@     @k@      Q@     `w@     �t@     �z@     @T@      b@     �A@      @@     �d@      ,@     0p@             @U@      "@      m@     �E@      :@       @      .@     �V@      8@     �d@     @d@     �m@     �C@      J@      @       @      K@      @      X@              E@       @     �X@      .@      @              @     �D@      @      K@      I@     �Y@      .@      ;@      @      @      F@      �?      J@              >@      �?     �Q@      @       @                      8@       @      :@      <@     �L@      "@      8@      @      �?      D@      �?      G@              6@      �?      K@      @       @                      3@              9@      8@     �I@      "@      @               @      @              @               @              0@      @                              @       @      �?      @      @              9@      @      @      $@      @      F@              (@      �?      <@       @       @              @      1@      �?      <@      6@      G@      @      1@      @      @      @      @      "@              $@      �?      &@       @                              &@      �?      ,@      &@      "@       @       @              �?      @      �?     �A@               @              1@      @       @              @      @              ,@      &@     �B@      @     @W@      =@      8@     @\@      "@     `d@             �E@      @     �`@      <@      6@       @      "@      I@      5@     @\@      \@      a@      8@      L@      8@      .@     �U@       @     �_@              @@      @     �Z@      4@      0@       @      @     �C@      *@     @T@     @R@     �\@      .@      .@              @      1@              ;@              @       @      5@       @       @      @      �?      @      "@      8@      *@      3@      @     �D@      8@      (@     @Q@       @     �X@              :@       @     �U@      2@       @      @       @     �A@      @     �L@      N@     �W@      &@     �B@      @      "@      ;@      @     �B@              &@      @      ;@       @      @              @      &@       @      @@     �C@      6@      "@      5@      �?      @      4@      @      6@              @              ,@       @      @              @      @      @      6@      7@      1@      @      0@      @      @      @              .@              @      @      *@               @              �?      @      @      $@      0@      @      @     @i@      Z@     @Q@     �d@      6@     �m@      @      ]@      6@      m@      N@      >@      4@      L@     �_@      F@     �i@      e@     �g@      E@     �b@     �Q@     �F@      ]@      $@     �h@             @T@      .@      g@     �D@      5@       @     �D@     @X@      >@     `d@      ]@      ^@      <@      U@     �A@      ?@     �M@      @      `@              L@      @     �]@      >@      "@      @      ;@      I@      @      U@     �N@      T@      5@      N@      2@      ,@     �B@      �?     �U@              ?@      @      H@      ,@      @      @      0@      9@      @      O@      =@      D@      (@      8@      1@      1@      6@      @     �D@              9@      �?     �Q@      0@      @              &@      9@      �?      6@      @@      D@      "@     �P@     �A@      ,@     �L@      @     @Q@              9@      $@     �P@      &@      (@      @      ,@     �G@      7@     �S@     �K@      D@      @      ,@      9@       @      (@      @      .@              �?       @      .@      @      @              @      ,@      "@      ,@      4@      1@       @     �J@      $@      (@     �F@              K@              8@       @     �I@      @      @      @      $@     �@@      ,@     @P@     �A@      7@      @     �I@      A@      8@     �I@      (@     �C@      @     �A@      @      H@      3@      "@      (@      .@      >@      ,@      F@      J@     �Q@      ,@     �D@      :@      .@     �I@      (@      C@      @      <@      @     �G@      .@      @      &@      ,@      ;@      *@     �D@     �D@     �P@      ,@      2@       @      "@      ,@      @      &@      @      *@      @      5@      @      @      "@      "@      &@      @      2@      $@      2@      @      7@      8@      @     �B@      @      ;@      @      .@              :@       @      �?       @      @      0@      @      7@      ?@     �H@       @      $@       @      "@                      �?              @              �?      @      @      �?      �?      @      �?      @      &@      @               @              @                      �?               @              �?      �?       @              �?      �?      �?                                       @       @      @                                      @                      @       @      �?               @              @      &@      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��  hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @#H1Y�@�	           ��@       	                   �6@k��h��@�           ��@                           @<sK@R           �@                            �?�0���@l           ��@������������������������       �xyK�@           �}@������������������������       ����Jl0@N           Ȁ@                          �1@,�H��@�           8�@������������������������       �)C�l�z	@�            �p@������������������������       �ɦ���Q@D           �@
                            �?�Aفa�@z            �@                          �<@6e���@�            px@������������������������       �ӈ����@�            �r@������������������������       �=!|l��@3            �V@                           �?Y�P�Q�@{           Ȃ@������������������������       �b1cvS�@�            �o@������������������������       ��'�Bƅ@�            �u@                           �?h ���n@�           ��@                           @"
֛
�@           �}@                           @E��nI@�            �z@������������������������       ��2���@�            �v@������������������������       �E�z]#@%             M@                           �?��- !@            �H@������������������������       ��P��r
@             ;@������������������������       �m�*���@             6@                           @ԆL�@�           ��@                           @~a(s �@/           }@������������������������       �Z�
���@�            0w@������������������������       �B�"�[�
@@            �W@                           @f�6'@q            `h@������������������������       ��TE�`�@G            �^@������������������������       �"jU!��@*             R@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@     �`@      V@     �t@     �E@     �|@      @     �o@      A@     @~@     �V@     �O@      ;@     �O@      k@     �O@     �w@     `r@     �|@     �U@     �m@     �T@     �H@     �p@      0@     �u@       @     �c@      8@     Pw@     �M@      D@      1@     �B@     �c@      C@     �o@      i@     Pv@      Q@     �`@     �B@      ;@     @g@      @      p@             �Z@      4@     `o@      5@      :@      $@      1@     @U@      3@     @e@      ]@     �o@      G@     �S@      8@      4@      \@      @     �\@             �G@      *@     `c@      *@      1@      @      ,@     �I@      .@      X@     �L@     @a@      B@      ?@      &@      (@     �L@              G@              :@      @     �Q@      @      ,@      @      @      @@       @     �@@      8@      R@      7@     �G@      *@       @     �K@      @     @Q@              5@      @     @U@      @      @       @      "@      3@      *@     �O@     �@@     �P@      *@     �L@      *@      @     �R@      �?     �a@             �M@      @      X@       @      "@      @      @      A@      @     �R@     �M@     �\@      $@      "@       @              6@              E@              6@              I@              @                      .@      @      5@      6@      J@       @      H@      &@      @      J@      �?     �X@             �B@      @      G@       @      @      @      @      3@             �J@     �B@     �O@       @     @Y@      G@      6@      T@      $@     �V@       @     �I@      @     �^@      C@      ,@      @      4@      R@      3@     �T@     @U@      Z@      6@      >@      <@      (@      >@      @     �A@       @      :@      @      C@      *@       @      @      1@      :@       @      ?@      @@      A@      ,@      :@      4@      �?      >@      @      ;@       @      2@              =@      &@       @      �?      &@      5@      @      :@      5@      =@      ,@      @       @      &@                       @               @      @      "@       @               @      @      @      @      @      &@      @             �Q@      2@      $@      I@      @     �K@              9@      �?      U@      9@      (@      @      @      G@      &@      J@     �J@     �Q@       @      7@       @      @      ?@              .@              ,@             �D@      ,@       @      �?              2@       @      5@      *@     �A@      �?      H@      $@      @      3@      @      D@              &@      �?     �E@      &@      @      @      @      <@      "@      ?@      D@     �A@      @     �[@     �H@     �C@     �P@      ;@      \@      �?      X@      $@     �[@      ?@      7@      $@      :@      N@      9@      _@     @W@      Y@      3@      I@      .@      1@      A@      $@      G@              H@      @     �M@      $@       @      @      @      4@      $@      B@      <@      N@      @     �F@      ,@      *@      >@      "@     �D@             �F@      �?     �H@      "@      @      @      @      3@      "@     �@@      :@      N@      @      C@      ,@      *@      3@      "@     �A@              B@      �?      G@       @      @      @      @      2@      "@      @@      :@      F@      @      @                      &@              @              "@              @      �?      �?                      �?              �?              0@       @      @      �?      @      @      �?      @              @      @      $@      �?      @              �?      �?      �?      @       @                      @              @      @      �?      �?              @      @       @      �?                      �?              �?              �?                              �?              �?              @                               @              @                      �?              @      �?                     �N@      A@      6@     �@@      1@     �P@      �?      H@      @      J@      5@      .@      @      3@      D@      .@      V@     @P@      D@      (@     �B@      2@      .@      >@      *@      J@      �?      C@      @     �@@      0@      "@      @      .@      8@      &@      N@      K@      3@      (@      6@      (@      .@      5@      *@     �D@      �?      @@      @      7@      (@      "@      @      .@      1@      &@     �H@      E@      1@      &@      .@      @              "@              &@              @              $@      @                              @              &@      (@       @      �?      8@      0@      @      @      @      ,@              $@              3@      @      @      @      @      0@      @      <@      &@      5@              5@      "@      @       @              $@              $@              *@      @      @      �?      �?      @      �?      *@      "@      0@              @      @       @      �?      @      @                              @      �?       @       @      @      (@      @      .@       @      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�	hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �3@)'n���@�	           ��@       	                    �?�����@�           ,�@                           @n�6�l�
@K           8�@                            @q�Y'/@�            0t@������������������������       �R�����	@�            �k@������������������������       �&w�Κ�@F             Y@                           @W}��@n            �h@������������������������       ���u�M@>            �\@������������������������       �o4��@0            �T@
                           @m��P\�@8            �@                           �?�|v��@�           �@������������������������       ��S�)�j@�            �j@������������������������       ��((��@�            �x@                           �?T���=@�            r@������������������������       ����N}k	@M            @^@������������������������       ���6@"@i             e@                           @XK��@7           |�@                            @���f*�@           �@                           @V���%@G           К@������������������������       ����<YP@8           ��@������������������������       �ޣO-J�@           p{@                           @��׋@�           ��@������������������������       �R@R�`@^           x�@������������������������       �Q��˟E@t             i@                           �?�j�r�	@            �I@������������������������       ��o���@             1@                          �6@�w}7j7@             A@������������������������       ���#@             1@������������������������       �����@
             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B         s@     @a@     @W@     �v@     �B@     0|@      @     �j@     �D@     �{@      \@     @P@     �@@     �S@     �l@     �N@     �w@     0r@     P}@     �Y@     �U@      9@      :@     �d@      @     �i@       @      S@      @     �e@     �@@      2@      @      ,@      U@      1@      `@     @Z@     �k@      :@      A@       @      @     �L@             @U@              =@      �?     �R@      &@       @      �?      @      E@      @      ;@      ?@     @Y@       @      @@       @      @      A@             �F@              &@              I@      &@       @      �?      @      ?@       @      5@      2@     �K@       @      .@       @      �?      ;@              A@              @              E@      @       @              @      7@              .@       @      E@       @      1@               @      @              &@              @               @       @              �?               @       @      @      $@      *@               @               @      7@              D@              2@      �?      9@                               @      &@      �?      @      *@      G@      @       @               @      &@              ;@               @              &@                                      @              @      @     �@@      @                              (@              *@              $@      �?      ,@                               @      @      �?              @      *@      @     �J@      7@      5@      [@      @     @^@       @     �G@      @     @X@      6@      0@      @      "@      E@      ,@     @Y@     �R@     @^@      2@      @@      .@      "@     @R@      @     �Q@       @      ?@      @     �S@      3@      0@      @      @      >@       @     �Q@     �D@     �U@      (@      *@      @      @      :@      @      *@       @      @      @      3@      (@       @              @      ,@       @      2@      3@      :@      $@      3@       @      @     �G@              M@              :@             �M@      @       @      @              0@      @     �J@      6@      N@       @      5@       @      (@     �A@              I@              0@              3@      @                      @      (@      @      >@     �@@     �A@      @      $@       @      �?      4@              8@              @              @      �?                              @              $@      7@      (@       @      &@      @      &@      .@              :@              $@              ,@       @                      @      @      @      4@      $@      7@      @      k@     @\@     �P@     @i@      A@     �n@      @      a@     �A@      q@     �S@     �G@      =@     @P@      b@      F@     @o@     @g@     �n@      S@     �j@     @\@     �P@     @i@      <@     �n@      @     �`@     �A@     `p@     @S@     �G@      ;@     @P@     `a@     �E@     �n@     `f@      n@      S@     �b@      T@      C@     �b@      "@     @h@      @     �S@      5@      h@     �H@      ?@      6@      D@     �Y@      B@     �f@     �[@      f@     �H@     �\@      P@      8@     @]@      @     �b@      @     �Q@      *@      b@      B@      :@      3@      =@     �S@      A@     @_@      S@      [@      C@     �B@      0@      ,@     �@@      @      F@               @       @      H@      *@      @      @      &@      7@       @     �L@      A@     @Q@      &@     �O@     �@@      =@      J@      3@     �I@              L@      ,@     @Q@      <@      0@      @      9@     �B@      @      P@     @Q@     �O@      ;@     �F@      6@      6@     �D@      ,@      A@             �D@      (@      A@      :@      &@      @      7@      9@      @      H@      J@     �F@      8@      2@      &@      @      &@      @      1@              .@       @     �A@       @      @               @      (@      @      0@      1@      2@      @      @                              @                      @              $@       @               @              @      �?      @      @      @                                                                       @              �?       @                              @              @      �?      @              @                              @                      �?              "@                       @              �?      �?      �?      @      @              @                              @                                      @                       @                      �?                       @                                              @                      �?              @                                      �?              �?      @       @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ/��@hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�W����@�	           ��@       	                    @&��B*�@�           ��@                          �3@�?��S�@�           ��@                           @�S��ʡ@�           (�@������������������������       ��Ϲ�kx@%           |@������������������������       �ƐE�a.@c            �d@                           �?��Jg�@g            �@������������������������       �r���@�            `k@������������������������       �9�WgD�@�            �v@
                          �0@��9��@�           ��@                           �?�'��	@P            �`@������������������������       ���i�t�@,             R@������������������������       ���=�@$            �O@                           �?���8�@�           ��@������������������������       ���~k	�@           �y@������������������������       �¦�0��@�           X�@                           �?	�L���@�           ؗ@                           @��'�@           0x@                           �?���L�@�            �p@������������������������       ������@I            @\@������������������������       ��f�\{o@n            �c@                           �?�ф��2
@K             ]@������������������������       �͔�~�	@/             Q@������������������������       ���/�@�@             H@                            @0���r�@�           ̑@                           @�m��@�           ��@������������������������       ���)z��@�           ��@������������������������       ���v�%@N             `@                          @@@X�ѵ�C@�            �u@������������������������       �z�GH'@�             t@������������������������       �쒚L�@             <@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       @t@     �a@     @T@     0u@      F@     �|@      $@     @k@      A@     �|@     @Y@     �N@      E@     �S@     �p@     �O@     �w@     �r@     �z@     @V@      f@     �Q@      E@      k@      3@     �u@       @     �a@      2@     �q@      G@     �G@      0@      @@      c@      6@     @o@     @f@     �q@     �D@      Y@      A@      <@     @`@      0@     �b@       @     �P@      ,@     �_@      ?@      2@      @      8@     �U@      1@      `@     @U@      [@      7@     �D@      ,@      .@     �U@      @     @S@      �?     �@@      @     �K@      0@      $@              @      G@      @      M@      J@      S@      $@      7@      @      @      K@      @     �O@      �?      8@      @     �H@      .@      $@              @      C@      @      E@      A@      M@      @      2@      @       @      @@              ,@              "@              @      �?                       @       @      @      0@      2@      2@      @     �M@      4@      *@      F@      (@      R@      �?      A@      "@      R@      .@       @      @      1@     �D@      $@     �Q@     �@@      @@      *@      A@      @      @      &@              :@      �?      2@              :@      @      �?       @      @      (@      @      6@      7@      4@      �?      9@      0@      $@     �@@      (@      G@              0@      "@      G@      $@      @       @      (@      =@      @     �H@      $@      (@      (@      S@      B@      ,@     �U@      @      i@              S@      @     �c@      .@      =@      (@       @     �P@      @     @^@     @W@     �e@      2@      @      @      @      @              :@              "@              ,@                               @      &@       @      &@      @      C@              @              �?      @              &@               @              $@                                      @              @              6@              �?      @      @                      .@              �?              @                               @      @       @      @      @      0@              R@     �@@      "@     �T@      @     �e@             �P@      @     �a@      .@      =@      (@      @     �K@      @     �[@     �U@      a@      2@      B@      @      �?     �A@      �?     �R@              :@      �?      F@      @       @              @      =@       @      ;@      >@      Q@       @      B@      :@       @     �G@       @     �X@             �D@      @     �X@       @      5@      (@      @      :@      �?     �T@     �L@     @Q@      $@     �b@     �Q@     �C@     �^@      9@     �[@       @     �R@      0@     �e@     �K@      ,@      :@      G@     �]@     �D@     �_@     �^@     �a@      H@     �C@      @      *@      9@       @      A@      �?      9@      @      H@      ;@      @      $@       @     �@@       @      >@      ;@      ?@      3@      2@      @      &@      3@       @      6@      �?      3@      @      =@      9@      @      $@       @      2@       @      0@      3@      7@      0@      "@       @      @      @       @       @      �?      $@       @      &@      (@      �?      @              @      @      @      &@       @      @      "@      @      @      (@              ,@              "@      �?      2@      *@       @      @       @      &@      @      &@       @      .@      (@      5@               @      @              (@              @              3@       @                              .@              ,@       @       @      @      ,@               @      �?              "@              @              "@      �?                              "@              @      @      @      @      @                      @              @                              $@      �?                              @              &@      �?      @             @[@      P@      :@     �X@      7@     @S@      @      I@      *@      _@      <@      &@      0@      F@     @U@     �@@     @X@     �W@     �[@      =@     �U@      K@      (@     �R@      (@      O@      @     �@@      @     @V@      ,@       @      @      6@     �P@      <@     @R@     �J@     @R@      1@     �P@      F@      &@     @R@       @     �H@      @      :@      @     @S@      *@       @      @      5@      L@      6@      J@     �D@     �P@      1@      5@      $@      �?      �?      @      *@              @              (@      �?               @      �?      &@      @      5@      (@      @              6@      $@      ,@      8@      &@      .@      @      1@      $@     �A@      ,@      @      &@      6@      2@      @      8@      E@     �B@      (@      6@      @      ,@      4@      @      .@      @      .@      $@     �@@       @      @      &@      6@      2@      @      7@     �C@     �A@      (@              @              @      @                       @               @      @                                              �?      @       @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��wphG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�����@�	           ��@       	                    @xe���@�           �@                            �?��4��v@Q           <�@                           �?�H�~��@`           �@������������������������       ���D�� @�           �@������������������������       �i�M&�@�           (�@                           �?�1'�@�            �x@������������������������       ���$�#;@n            @e@������������������������       �>�_pX�
@�            `l@
                           �?�o�b�@�           ��@                           �?��G*� @           �y@������������������������       ��M���|@             G@������������������������       �� �=]@�            �v@                           @�<��@�           x�@������������������������       �T��n@-           @~@������������������������       ���h�@d            `e@                           @OǷ@�           H�@                           �?����hl@�           Ȉ@                           �?H�-~�@)           �}@������������������������       �,)�q�@G            �\@������������������������       �wpɭ?�@�            �v@                           @t����@�            �s@������������������������       ��L�6��@�            `n@������������������������       �d�M�Q@1            �R@                           @��� #c@�            �s@                           �?]��v�@�            �h@������������������������       �f.�Q�@/            �P@������������������������       ��G�@W            ``@                          �5@cu,��@D            �\@������������������������       �}Q<���@             G@������������������������       ��X��rS@*            @Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       pu@     �a@      U@     @u@     �E@     �}@      @     �m@      @@     �{@     @_@     �H@      @@     �Q@     �m@      N@     �x@     Ps@     �y@     �S@      l@     �Y@      E@      n@      ;@     0v@      @     �d@      .@     �u@     �S@      =@      :@      C@     `f@      A@     Pr@     �k@     0u@      I@      c@     �L@      <@     �a@      &@     �o@      @     �X@      @     �n@      E@      ,@      2@      7@     �Z@      .@     �g@     �\@     �h@      ;@     @`@      I@      4@     �]@       @     �e@      @     �R@      @     �f@     �B@      $@      .@      5@      T@      ,@     �a@     �U@     �c@      6@     �M@      8@      ,@     �J@      @      V@      @      F@      �?      [@      $@      @      $@      @     �C@       @     �R@     �C@     @S@      "@     �Q@      :@      @     �P@       @     �U@      �?      >@      @      R@      ;@      @      @      1@     �D@      (@      Q@     �G@     �S@      *@      7@      @       @      7@      @     �S@              9@      �?     �P@      @      @      @       @      :@      �?      G@      =@      E@      @      $@                      "@      @      ?@              *@      �?      8@      @      �?               @      $@      �?      (@      *@      @@      @      *@      @       @      ,@             �G@              (@              E@              @      @              0@              A@      0@      $@       @     �Q@     �F@      ,@     �X@      0@     �Y@             @P@      $@     @Y@      B@      .@       @      .@     @R@      3@     @Z@     �Z@     �a@      7@      ?@      1@      @     �C@      ,@     �F@              &@      @      @@      *@       @      @       @     �D@      @      A@      G@     �K@      &@       @              �?      �?              @                              @                                      @               @      @      0@              7@      1@      @      C@      ,@      E@              &@      @      =@      *@       @      @       @     �A@      @      @@      D@     �C@      &@      D@      <@      $@     �M@       @      M@              K@      @     @Q@      7@      *@      @      *@      @@      .@     �Q@      N@     �U@      (@      <@      9@      @      I@       @      C@             �I@      @      L@      1@       @       @      @      8@      ,@      D@     �E@     �M@       @      (@      @      @      "@              4@              @              *@      @      @       @      @       @      �?      ?@      1@      ;@      @     �]@      D@      E@      Y@      0@     �]@       @     �R@      1@     @W@     �G@      4@      @     �@@     �L@      :@     �Y@      V@      S@      <@     �U@      7@      ;@     �R@      $@     @W@       @     �H@      .@     �I@      D@       @       @      <@      A@      6@     �S@     �Q@     �L@      5@      K@      2@      8@     �J@      @     �B@       @      =@      *@      5@      :@      @      �?      6@      ,@      *@      J@     �F@      :@      *@      0@      @      @      2@       @      &@      �?      @      �?      @      @      �?              �?      @      @      &@      @      @      @      C@      (@      1@     �A@      @      :@      �?      6@      (@      0@      5@      @      �?      5@      &@      $@     �D@     �C@      5@       @     �@@      @      @      6@      @      L@              4@       @      >@      ,@       @      �?      @      4@      "@      :@      :@      ?@       @      <@      @      @      ,@      @     �G@              0@       @      ;@      $@       @                      $@      "@      8@      2@      4@      @      @       @               @              "@              @              @      @              �?      @      $@               @       @      &@       @      @@      1@      .@      9@      @      9@              :@       @      E@      @      (@      @      @      7@      @      9@      1@      3@      @      9@      "@      (@      *@       @      *@              6@       @      >@      @      @      @      @      $@      �?      *@      (@      (@      @      (@      �?      @      @              @              "@              @      �?      @      �?      �?              �?      @      @      @      �?      *@       @      @      @       @      "@              *@       @      7@      @      @       @       @      $@              "@       @      @      @      @       @      @      (@      @      (@              @              (@       @      @      �?       @      *@      @      (@      @      @       @       @      @               @              @               @              @      �?       @              �?      @       @      (@      �?      @       @      @      @      @      $@      @      @               @              "@      �?      @      �?      �?      $@      �?              @      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJz̲6hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @eHL��@�	           ��@       	                   �6@}FN1X@�           ,�@                           �?Q���+@_           ��@                          �3@� ts�@�           x�@������������������������       ��j�Ơ
@           �|@������������������������       �)mx4@�             p@                          �0@�����@�           t�@������������������������       ���R��L@;            �W@������������������������       ����@e           ��@
                           �?�@3�@�           ��@                           �?]�^^*@*           �|@������������������������       �ĕ�X7@j            `e@������������������������       �G���3�@�            r@                            �?�e1��?@k           ��@������������������������       �tׇ�K@�             y@������������������������       �ſ<�+�@n            �i@                           @F�2B��@�           ̐@                          �;@0�4�@�           ��@                           �?�-�^3@�           �@������������������������       �c�	D��@           �y@������������������������       �VV=�ɽ@�            @r@                           �?�##fm@6             V@������������������������       ���6N�@+            �Q@������������������������       ��V���@             2@                           �?�	�S�@�            �q@                           @}҈=�@G             [@������������������������       �hGr:g@.            �P@������������������������       ����\yu
@            �D@                          �8@���p��@t            @f@������������������������       �ĶQD)	@M             ^@������������������������       �?/��4@'             M@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �b@      V@     0u@      F@     �~@      @     �o@     �A@     }@     �Z@      Q@      C@     �R@      m@     �R@     Pv@     �r@     �y@     �O@     `k@     @Y@     �I@      p@      6@      x@      @     �d@      9@     Pv@     @P@      K@      =@     �A@     `e@     �L@     �p@      j@     0t@      F@     �]@     �F@      7@     �c@      @     �r@             @Y@      .@     �n@      B@     �D@      *@      $@      X@      <@     `d@      `@     �k@      ;@      H@      .@       @     �N@       @     �a@              D@      @     �Z@      @      *@       @      @      A@      �?     �P@     �K@     �Y@      "@      5@      @      �?      D@      �?      W@              ?@      @     �T@      �?      "@       @       @      7@      �?      E@      A@     �P@      @      ;@      &@      @      5@      �?     �H@              "@              7@       @      @              @      &@              9@      5@     �A@      @     �Q@      >@      .@     �W@      @     �c@             �N@      "@     �a@     �@@      <@      &@      @      O@      ;@      X@     @R@     @^@      2@      @      �?               @              4@              (@              @              �?                      @               @       @      6@             �P@      =@      .@     �U@      @      a@             �H@      "@      a@     �@@      ;@      &@      @     �K@      ;@      V@     @P@     �X@      2@     @Y@      L@      <@      Y@      1@     @V@      @     �O@      $@     �[@      =@      *@      0@      9@     �R@      =@     �Y@     @T@      Y@      1@      6@      B@      2@      =@      &@      >@      @      A@      �?      G@      ,@      $@      &@      ,@      C@      *@     �I@     �@@      B@       @      &@      @      ,@      @      @      $@      @      0@      �?      5@       @       @      @      �?      3@      @      4@      &@      &@       @      &@      @@      @      6@      @      4@       @      2@              9@      (@       @      @      *@      3@       @      ?@      6@      9@      @     �S@      4@      $@     �Q@      @     �M@              =@      "@      P@      .@      @      @      &@     �B@      0@     �I@      H@      P@      "@     �L@      0@      @      C@      @      @@              8@      @      D@      ,@      @      @      &@      9@       @     �@@      ?@     �H@      @      6@      @      @     �@@       @      ;@              @      @      8@      �?               @              (@       @      2@      1@      .@      @     @X@     �H@     �B@     �T@      6@     �Z@       @      V@      $@      [@     �D@      ,@      "@      D@     �N@      1@      W@      W@     �U@      3@     �P@      =@      ;@      O@      1@     �U@       @      P@      @     �Q@     �B@       @      @      B@     �F@      (@      N@     �R@      Q@      (@      K@      4@      6@     �H@      .@     �U@       @     �N@      @     �P@     �B@       @      @      >@      C@       @      K@     �P@      P@      "@      B@       @      5@      6@      ,@      F@       @      @@      @      A@      9@      @      @      9@      8@      @      <@      @@      B@      @      2@      (@      �?      ;@      �?     �E@              =@             �@@      (@      �?              @      ,@       @      :@      A@      <@      @      (@      "@      @      *@       @                      @       @      @                              @      @      @      @      "@      @      @      $@      @      @      "@                              @       @                                      @      @      @      @      "@      @               @       @              @       @                                      @                                       @                                      @      ?@      4@      $@      5@      @      4@              8@      @      C@      @      @      @      @      0@      @      @@      1@      3@      @      1@      @      @      ,@       @      @              "@       @      0@      @      @       @              �?              @      "@      $@              $@      @       @      @              @              @               @              @       @                              @      @      "@              @      �?      �?      @       @                      @       @       @      @                              �?               @       @      �?              ,@      *@      @      @      @      0@              .@       @      6@      �?      @      �?      @      .@      @      :@       @      "@      @      $@      &@      @      @      �?      &@              *@       @      1@      �?       @              �?      @      @      4@      @              @      @       @      @      @       @      @               @              @              �?      �?      @       @              @       @      "@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�4ghG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?6�H6F�@�	           ��@       	                     @m�#��r@�           d�@                           @�4��У@�           h�@                          �4@^�rG�,@Q           ��@������������������������       �����K@�            `l@������������������������       �_̋��@�            �s@                           @b\�Լ-
@l           ؁@������������������������       �D`E���	@�            �w@������������������������       �_�,��	@}            @h@
                           �?Ý����@�            �w@                           �?_��;�@�             j@������������������������       �����|6@j            �d@������������������������       ��^X�*@             F@                           �?�ւ<�@g            �e@������������������������       �����~B@:            @W@������������������������       �!�NF)�@-            �T@                           �?(D���@           �@                          �5@e�x��@�           ��@                           @�s����@           P|@������������������������       �#��(2n@�            @q@������������������������       �L�!S�v@d             f@                           @��_@�           ȁ@������������������������       �wѬ��@5           �|@������������������������       �L���"@K            @[@                           @�nu�"�@y           ȕ@                           @�Hl�s�@a           $�@������������������������       �@��J{_@�           �@������������������������       ��+��/�@i           `�@                           �?���u	@            �D@������������������������       ���ܤ�@
             .@������������������������       �jޱnu:@             :@�t�b��     h�h5h8K ��h:��R�(KKKK��h��B`        v@      \@      U@     �t@     �B@     P�@      "@     �j@      <@     p|@     �Z@      P@      B@      Q@      l@      N@      x@     �s@      z@     @X@     �\@     �A@     �B@      [@      &@     �o@      �?      V@      @     �e@     �G@      0@      @      3@     �U@       @     �b@     @^@      f@      G@      T@      7@      6@     �V@      @     �i@      �?     �M@             �`@      ?@      (@      @      @      K@      @      ]@     �U@      b@     �@@     �C@      1@      &@     �C@      @      U@      �?      C@             �Q@      8@      "@      @      @      :@      @      H@      E@      G@      >@      3@      @      @      3@      �?      >@              1@             �D@      @      @                      $@              .@      9@      5@      "@      4@      *@      @      4@      @      K@      �?      5@              =@      4@      @      @      @      0@      @     �@@      1@      9@      5@     �D@      @      &@     �I@             �^@              5@             �O@      @      @               @      <@      �?      Q@     �F@     �X@      @      3@       @      @      E@             �W@              .@             �D@      @       @              �?      5@      �?     �F@     �@@     �H@       @      6@      @      @      "@              <@              @              6@      @      �?              �?      @              7@      (@     �H@      �?      A@      (@      .@      2@      @      G@              =@      @      D@      0@      @              (@     �@@      @      @@      A@     �@@      *@      0@       @      *@      (@      �?      1@              7@      @      3@      @      @              $@      &@      @      5@      4@      2@      @      $@      @      $@      "@              *@              6@      @      3@      @       @              @      $@      @      4@       @      1@       @      @      @      @      @      �?      @              �?      �?                       @              @      �?              �?      (@      �?      �?      2@      @       @      @      @      =@              @              5@      &@                       @      6@              &@      ,@      .@      $@      @               @      @       @      1@              @              @      @                              0@              @      @      &@      "@      &@      @               @       @      (@               @              ,@       @                       @      @              @       @      @      �?     �m@     @S@     �G@     �k@      :@     �p@       @     �_@      8@     �q@     �M@      H@      @@     �H@      a@      J@     �m@      h@      n@     �I@     �X@      9@     �B@     �X@      5@     �R@       @     �L@      0@     @[@      5@      :@      ,@      ?@      K@      7@     �V@     �S@     �[@      =@      H@      @      5@      C@      $@     �D@              1@      @      D@      &@      .@      �?      @      5@       @      E@     �J@     �J@      1@      9@      �?      @      :@      $@      <@              @      @      8@       @      $@      �?      @      (@      @     �@@      :@     �A@      *@      7@      @      2@      (@              *@              &@      �?      0@      @      @              �?      "@      @      "@      ;@      2@      @     �I@      4@      0@     �N@      &@      A@       @      D@      &@     @Q@      $@      &@      *@      8@     �@@      .@      H@      9@     �L@      (@      C@      ,@      0@      K@      @      ;@       @     �B@      "@     �N@      "@       @      &@      5@      8@      @      B@      4@     �F@      $@      *@      @              @      @      @              @       @       @      �?      @       @      @      "@      "@      (@      @      (@       @     `a@      J@      $@     �^@      @     @h@             @Q@       @     �e@      C@      6@      2@      2@     �T@      =@     @b@     �\@     ``@      6@     �`@      J@      $@     �^@      @      h@             �P@       @      e@      C@      6@      ,@      2@     @T@      ;@     �a@     @Y@      `@      6@     �Q@      A@      @     �R@      @     �Y@              F@       @     �[@      ;@      1@      "@      "@     �G@      7@     @Q@     �P@      O@      (@      P@      2@      @      H@      �?     @V@              7@              M@      &@      @      @      "@      A@      @     @R@     �A@     �P@      $@      @                                       @               @              @                      @               @       @      @      *@      @               @                                                       @              @                                       @               @      @      �?               @                                       @                               @                      @                       @       @      $@       @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJc,� hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?i��0l�@�	           ��@       	                   �:@�I��x�@           ��@                            �?�6mUKd@7           x�@                          �2@�W��z�@�            y@������������������������       ����/
@7             U@������������������������       ��W\�P3@�            �s@                           �?���ecR@@           h�@������������������������       �P��T�@�            �v@������������������������       ��P�$*@j           �@
                          �?@�f�A!@�             u@                           �?�xBO@�             o@������������������������       ��W�ˀ@7            �S@������������������������       �����m@o            @e@                           �?#|�}��@:            @V@������������������������       ����JF�@             9@������������������������       �~����+@)             P@                          �4@$쑾�@�           ��@                           @%�b@�           ؒ@                          �3@��TZ�@6           @@������������������������       ��Q���@�            �v@������������������������       �0��t�@Q            �`@                           �?>�o�-�@�           �@������������������������       ����O�?
@�            �w@������������������������       ��>��@�            0t@                            @����g@�           ��@                           �?�~ϐ�1@&           Ȋ@������������������������       �xX6|�@�            �o@������������������������       �T4c��@�           Ђ@                           @�&���@�            @i@������������������������       �Wx�н@[             a@������������������������       �����.9
@%            �P@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       `u@     �_@     �Z@     @u@     �G@     p~@      @     `m@      >@     `z@     �^@     �K@      A@     �J@      n@      R@     @w@     �r@     �z@      W@     �c@     �K@     @Q@     �a@      @@      b@      @     �`@      8@     @a@      I@      9@      2@     �@@     �X@      D@      b@     `a@     `c@     �F@      a@     �C@      G@     �[@      =@     �`@      �?     @V@      5@     �\@     �C@      2@       @      7@     �S@      :@     �^@     �Z@     @`@     �B@      ?@      (@      $@      H@      &@     �E@      �?      <@      "@      ?@      @      @      �?      @      :@      "@      :@      B@     �I@      ,@      "@              @      (@      @      "@              @              @                      �?      �?      @              �?       @      4@              6@      (@      @      B@       @      A@      �?      8@      "@      :@      @      @              @      4@      "@      9@      <@      ?@      ,@     �Z@      ;@      B@      O@      2@      W@             �N@      (@      U@      B@      (@      @      2@      J@      1@     @X@     �Q@     �S@      7@      A@      ,@      6@      6@       @     �E@              <@      @      <@      0@      �?      @      "@      7@      @      D@      =@      =@      (@      R@      *@      ,@      D@      0@     �H@             �@@       @      L@      4@      &@      @      "@      =@      ,@     �L@     �D@      I@      &@      4@      0@      7@     �@@      @      "@      @     �E@      @      7@      &@      @      $@      $@      4@      ,@      6@     �@@      9@       @      .@      @      ,@      :@      @      @      @      C@      @      4@       @      @      @      @      3@      "@      1@      6@      8@      @      @      �?      "@      @      @      �?      @      $@      @      @      @               @      @      @      �?      @       @       @              $@      @      @      4@               @      �?      <@              ,@      �?      @       @       @      0@       @      (@      4@      0@      @      @      &@      "@      @              @              @              @      @       @      @      @      �?      @      @      &@      �?      @              �?      @      �?                              @                      @              @      @              @                      �?              @      $@      @      @              @              �?              @               @      @       @      �?              @      &@              @      g@      R@     �B@     �h@      .@     pu@             �Y@      @     �q@     @R@      >@      0@      4@     �a@      @@     `l@     �c@     @q@     �G@      R@      >@      0@     �_@       @     �f@              P@      �?      e@      7@      &@      @      @     �Q@      2@     �_@     �T@     �f@      3@      2@      &@      @     �P@             �O@              3@             �S@      (@      @      @      @      =@      0@     �M@      @@     �O@      ,@      2@      @      @     �H@              I@              *@              M@      &@      �?              @      ;@      "@      I@      4@      C@      $@              @      @      1@              *@              @              5@      �?       @      @               @      @      "@      (@      9@      @      K@      3@      "@      N@       @     �]@             �F@      �?     @V@      &@       @      @      �?      E@       @     �P@      I@      ^@      @      ;@      @      @     �C@       @     �P@              1@             �H@      @      @                      3@             �D@      2@     �T@       @      ;@      (@      @      5@              J@              <@      �?      D@      @      @      @      �?      7@       @      :@      @@      C@      @     @\@      E@      5@     �Q@      *@     @d@             �C@      @      ]@      I@      3@      "@      ,@      R@      ,@     @Y@     @S@     @W@      <@     �U@      A@      1@      L@      "@      b@              @@      @     @U@      D@      0@      @      (@      F@      (@     �U@     @P@     �U@      6@      8@      @      &@      ,@       @      H@              1@              @@      @                              *@              <@      3@      <@      "@     �O@      <@      @      E@      @      X@              .@      @     �J@      B@      0@      @      (@      ?@      (@      M@      G@      M@      *@      :@       @      @      .@      @      2@              @              ?@      $@      @      @       @      <@       @      .@      (@      @      @      1@      @      @       @      @      1@              @              7@      $@      �?       @      �?      (@       @      (@      @      @      @      "@      @              @              �?                               @               @       @      �?      0@              @      @      @       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJU��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@��Iٿ@�	           ��@       	                    �?�6=�mw@           d�@                            �?-��h@           �{@                           @����C�@�            `j@������������������������       ��w\�~}@o             e@������������������������       �(^���@            �E@                          �2@���K4�@�            �l@������������������������       ���î�@g            @d@������������������������       ����>�@%            �P@
                           �?�o�v@h           �@                           @u��<�
@:           }@������������������������       ��b^ް
@�            0q@������������������������       �Ʃx�f
@{            �g@                           �?�}T��@.            }@������������������������       �5�Y�
@e            `c@������������������������       �j�G��Y@�            Ps@                          �7@j�+k}�@C           �@                           �?�2,��@1           d�@                          �4@�m���@'           }@������������������������       ����s@^            �b@������������������������       ��n�(�@�            �s@                           �?�æex@
           @�@������������������������       ��RD\ܟ@�            �t@������������������������       ����4�@@           �@                           �?\�>VG�@           \�@                            �?�L�h~@�            �u@������������������������       ����MhB@x            @h@������������������������       �u� #d�@h            @c@                          �8@h.k F�@2           ؋@������������������������       �zVHۑ@�            `k@������������������������       �"��]@�            �@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �`@     �X@     �u@     �D@     �|@      @     �l@      =@     �{@     @X@     �P@     �F@     @Q@     `m@     �Q@     �w@     �r@      }@      S@     �W@      7@      ;@     @b@      @     `j@             @R@      @      f@      5@      1@      @      (@     �S@      2@     �`@     �Z@     �i@      .@      C@      "@      4@     �A@      @      L@              0@       @      A@      $@      @      @      @      =@      @      =@     �J@     �S@      @      0@      @      "@      9@              ;@              @       @      1@      @      @       @       @      &@      �?      @      8@     �H@      @      (@      @      @      7@              3@              �?       @      1@      @      @       @       @      "@      �?      @      6@      ?@      @      @      �?      @       @               @               @                                                       @              �?       @      2@              6@      @      &@      $@      @      =@              *@              1@      @              �?      @      2@      @      6@      =@      >@      @      *@      @      @      $@      @      .@              (@              ,@      @              �?      �?      0@      @      ,@      7@      0@      @      "@              @                      ,@              �?              @      @                      @       @               @      @      ,@              L@      ,@      @     �[@       @     `c@             �L@      �?     �a@      &@      (@              @      I@      (@     @Z@      K@     �_@       @      >@       @      @     �L@       @     �R@             �A@             �P@              �?              �?      9@      @     �H@      @@     @Q@      @      (@      @      @     �B@      �?      F@              (@             �B@              �?              �?      0@      @      >@      1@      I@      @      2@       @       @      4@      �?      ?@              7@              >@                                      "@              3@      .@      3@      �?      :@      @      �?      K@              T@              6@      �?     �R@      &@      &@              @      9@       @      L@      6@     �L@      @      *@                      3@              A@              @      �?      3@      @      @               @       @       @      "@       @      7@       @      *@      @      �?     �A@              G@              .@              L@      @      @              @      1@      @     �G@      ,@      A@       @     �m@     @[@     �Q@     �i@      B@     �n@      @     �c@      :@     �p@      S@     �H@      E@     �L@     �c@      J@     @n@     �g@     Pp@     �N@      `@      I@      8@      ^@      *@     @c@      @      N@      2@      a@      ?@     �@@      $@      3@      R@      <@     �b@     �W@      `@      B@     �H@      *@      ,@      A@       @      N@      @      7@      @     �B@      ,@      @              @      B@      �?     �L@      A@     �L@      1@      (@      �?      @      $@       @      0@              @      @      ,@       @      �?                      @      �?      $@      5@      7@      "@     �B@      (@       @      8@              F@      @      0@              7@      @      @              @      =@             �G@      *@      A@       @     �S@     �B@      $@     �U@      &@     �W@             �B@      .@     �X@      1@      =@      $@      (@      B@      ;@     �V@      N@     �Q@      3@      D@      @      @     �C@      @      C@              ,@      @     �@@      $@      $@      @      @      3@      @      8@      9@      A@      @     �C@      @@      @     �G@      @      L@              7@       @     �P@      @      3@      @      "@      1@      4@     �P@     �A@     �B@      ,@     �[@     �M@     �G@      U@      7@     �V@      @     �X@       @      `@     �F@      0@      @@      C@      U@      8@     �W@      X@     �`@      9@      1@      "@      3@      &@      @      >@      �?     �A@       @     �J@      0@       @      .@      @      3@      @      =@      :@     �B@      "@      @      @      0@      @      @      3@              2@              C@      @      �?      ,@      @      (@      �?      2@      @      4@      �?      $@      @      @      @              &@      �?      1@       @      .@      "@      @      �?      �?      @      @      &@      4@      1@       @     @W@      I@      <@     @R@      4@     �N@       @     �O@      @      S@      =@       @      1@      A@     @P@      3@     @P@     �Q@      X@      0@      1@      1@      @      3@      @       @               @      @      :@      @      �?      @      0@      .@      @      7@      5@      &@      "@      S@     �@@      7@      K@      .@     �J@       @     �K@       @      I@      8@      @      ,@      2@      I@      *@      E@     �H@     @U@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��4thG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��RC!�@�	           ��@       	                   �3@#C{?W�@/           ��@                            @�`5�;@a           P�@                            �?b;�u_
@
           �x@������������������������       ����t�@^             b@������������������������       �Q5T�@�             o@                           �?�͸B�4@W            @`@������������������������       �{��כx
@-            @Q@������������������������       �?�Ǣ¸
@*            �N@
                          �7@u����@�           (�@                            �?ދf<@@            `z@������������������������       ��{#+%�@�            �n@������������������������       �&����@n             f@                            @����d@�            �s@������������������������       �ã���@�            �l@������������������������       �kq-HYO@=            �V@                            �?��i�.�@�           ��@                           �?&�4Rn�@�           X�@                          �:@��[��@�            �s@������������������������       ��ښ��c@�            �p@������������������������       �����*�@             G@                           �?ܶ\�R@(           �|@������������������������       �ćB�5�@�            `l@������������������������       �.�7�x�@�            �m@                          �6@<�-���@�           <�@                          �5@S����@�           `�@������������������������       ����#�@M           ��@������������������������       �Z4��@a            �d@                           @)<�Y(�@�           ��@������������������������       �FKQE�@@           `~@������������������������       �X~yb
@�            q@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       `t@     �a@      W@     �v@     �@@      @      @      k@      9@      |@      [@     �M@      H@     �P@     �o@      R@      v@     �r@      {@      S@     @Y@      ;@      ?@     �[@      @     �g@             @T@      @     @b@      ?@      .@      .@      *@     �W@      &@     @]@     �S@     �c@      A@      B@      @       @      I@              Z@              >@      �?     �P@      @      @      �?       @      C@      @      C@      ?@      V@      @      9@      @      @     �D@             �S@              5@      �?     �I@       @      @                      :@       @      <@      ;@      R@      @      *@              @      2@              7@              &@              .@       @       @                      $@       @       @      ,@      3@      @      (@      @              7@              L@              $@      �?      B@              @                      0@              4@      *@     �J@              &@              @      "@              9@              "@              0@      @              �?       @      (@      @      $@      @      0@      @      @               @      @              1@              @              @      @              �?               @              "@       @      "@      @       @               @      @               @              @              *@      �?                       @      @      @      �?       @      @             @P@      6@      7@      N@      @     �U@             �I@       @     �S@      8@      $@      ,@      &@      L@      @     �S@      H@     �Q@      <@      E@      (@      ,@     �D@      @      M@              7@              G@      (@      �?               @      =@              L@      :@      >@      4@      ;@       @      @     �@@              B@              &@              6@      @                      @      *@             �A@      4@      5@      @      .@      @      "@       @      @      6@              (@              8@      @      �?              @      0@              5@      @      "@      .@      7@      $@      "@      3@      @      <@              <@       @     �@@      (@      "@      ,@      @      ;@      @      7@      6@      D@       @      1@      @      @      (@       @      6@              3@              ;@      @      @      ,@      �?      4@      @      2@      2@      9@      @      @      @      @      @      �?      @              "@       @      @      @      @               @      @       @      @      @      .@      @      l@     �\@     �N@     �o@      :@      s@      @     �`@      6@     �r@     @S@      F@     �@@     �J@      d@     �N@     `m@     �k@      q@      E@      G@     �K@      0@      O@      @     �S@      �?      @@      @     @Z@      3@      &@      .@      6@     �B@      2@     �N@     �L@     �\@      2@      4@      2@      (@      6@      @     �A@      �?      $@      �?      J@      @      @      &@      @      4@       @      <@      :@      ;@      @      4@      0@      @      6@      �?      @@      �?      "@              H@      @      @       @       @      4@              9@      6@      8@      @               @      @              @      @              �?      �?      @      �?              @      @               @      @      @      @              :@     �B@      @      D@       @     �E@              6@      @     �J@      ,@      @      @      1@      1@      $@     �@@      ?@     �U@      (@      $@      4@       @      "@       @      1@              *@      @      3@      @      @       @      (@      "@      @      0@      8@      D@      &@      0@      1@       @      ?@              :@              "@              A@       @       @       @      @       @      @      1@      @     �G@      �?     `f@     �M@     �F@     �g@      3@     �l@      @     �Y@      1@     �h@      M@     �@@      2@      ?@      _@     �E@     �e@     �d@      d@      8@     �W@      <@      .@      ]@      $@     @f@      �?     �N@      @     �_@     �@@      ;@       @      &@     @R@      =@     �X@     @W@     �W@      (@     �S@      8@       @     �Y@       @     @b@      �?     �H@      @     @[@      7@      5@       @      &@     �L@      8@     �T@     �V@     �V@      (@      0@      @      @      ,@       @      @@              (@       @      2@      $@      @                      0@      @      0@      @      @              U@      ?@      >@     �R@      "@      I@      @      E@      $@     �Q@      9@      @      0@      4@     �I@      ,@     �R@      R@     @P@      (@      F@      4@      >@      I@      @      >@       @     �A@      "@      D@      1@      @      $@      ,@      >@      @      F@      J@     �B@      @      D@      &@              8@       @      4@      �?      @      �?      >@       @       @      @      @      5@      "@      ?@      4@      <@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�\RF�f@�	           ��@       	                    �?8a�Ԙ@           ��@                          �8@DXO��@e           H�@                          �2@@^�v@           y@������������������������       ��˥��O@U            �`@������������������������       �@�oâ@�            �p@                           �?�)�w�@a             c@������������������������       �8e.��I@              F@������������������������       �9A��@A             [@
                            @Fi	��@�           �@                           �?sQ�hOV@i           ��@������������������������       �m�t|."@n            �h@������������������������       �H��о�@�            �y@                           �?�ԾX�@:           �~@������������������������       �[� 'Y@j            �d@������������������������       ���ǌA<@�            @t@                           �?$�ً5@�           ��@                          �9@	�An�;@           `�@                          �3@B����@�           ��@������������������������       �/��d�
@�            �x@������������������������       �kBG��d@�            �t@                          �<@�T=��@;            �U@������������������������       ��2�ec�@*             O@������������������������       ��ܩQ/|@             8@                            �?'ך��@�           ��@                           @/���"�@           �@������������������������       ��6��Ѫ@�           ��@������������������������       �kBT�
@<            @T@                            @ ��/B�@�           X�@������������������������       �ⷠ_|@�            �t@������������������������       �l1?J�\@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@      a@     �U@     �w@      B@     @@      @      i@      9@     0|@      \@      I@      >@      M@     �p@     �M@     �v@      s@     �z@      U@      b@     �O@     �I@     `d@      7@     �c@      @     �W@      6@     �c@     �K@     �A@      0@     �A@     @[@      :@      b@     �a@      d@      F@     �K@      4@      8@     �M@      @      L@      @      ;@      �?     �F@      3@       @      �?      @      C@      $@      J@     �H@     @P@      &@      E@      ,@      5@      I@      @      F@              (@      �?      <@      0@      @              @      5@      $@     �B@      >@     �J@       @      0@      �?      @      5@      �?      (@              @              $@      @      �?              �?      "@      @      @      .@      ;@              :@      *@      .@      =@      @      @@              "@      �?      2@      *@      @              @      (@      @      @@      .@      :@       @      *@      @      @      "@              (@      @      .@              1@      @      @      �?      �?      1@              .@      3@      (@      @      @      �?      �?       @              @       @      @               @      �?              �?      �?      @              @       @       @               @      @       @      @              "@      �?      (@              "@       @      @                      ,@              (@      &@      $@      @     @V@     �E@      ;@      Z@      3@     @Y@       @      Q@      5@      \@      B@      ;@      .@      =@     �Q@      0@      W@     �W@      X@     �@@      D@      A@      *@     �P@      &@     �N@      �?      =@       @     @R@      ,@      2@      @      *@      @@      "@     �I@      G@     �N@      4@      .@      @      @      ,@      @      8@      �?      ,@      �?      7@      @      "@      �?      �?      *@      @      8@      @      *@      $@      9@      ;@      @      J@      @     �B@              .@      @      I@      "@      "@      @      (@      3@      @      ;@     �C@      H@      $@     �H@      "@      ,@      C@       @      D@      �?     �C@      *@     �C@      6@      "@      &@      0@     �C@      @     �D@      H@     �A@      *@      2@      @      @      ,@      �?      1@              ,@      @      0@      $@              @      @      &@              *@      1@      ,@      @      ?@      @      "@      8@      @      7@      �?      9@       @      7@      (@      "@       @      *@      <@      @      <@      ?@      5@      $@     �g@     @R@     �A@     `k@      *@     pu@             @Z@      @     `r@     �L@      .@      ,@      7@     �c@     �@@     �k@      d@     �p@      D@     @P@      2@      (@     �O@      @     �a@              F@              ]@      2@      �?              "@     @P@      @     �Q@      L@     �Y@      5@      P@      2@      $@      L@       @      `@              D@             @X@      ,@                      @     �N@      �?      P@     �K@     �V@      1@      >@      �?      @      @@       @     @T@              9@              J@      @                      @     �@@      �?     �A@      6@     @P@      @      A@      1@      @      8@              H@              .@             �F@      $@                       @      <@              =@     �@@      :@      &@      �?               @      @      �?      (@              @              3@      @      �?               @      @      @      @      �?      &@      @      �?               @      @      �?      @              @              "@      @      �?              �?      @      @      @              $@      @                               @              @                              $@                              �?              @      �?      �?      �?             �^@     �K@      7@     �c@      $@     @i@             �N@      @     @f@     �C@      ,@      ,@      ,@     �W@      :@      c@     @Z@     �d@      3@     �S@      B@      0@     @T@      @     @Y@              >@      �?     �W@     �@@      $@      $@      &@      H@      &@     �V@     �Q@     @X@      (@     �Q@      @@      ,@      T@      @     @W@              2@      �?     @V@      <@      $@      @      &@      C@      &@     @T@     �O@     �V@      (@      @      @       @      �?               @              (@              @      @              @              $@              "@      @      @             �F@      3@      @     �R@      @     @Y@              ?@       @     �T@      @      @      @      @      G@      .@      O@     �A@      Q@      @      5@      @      @      D@      @     �P@              .@       @     �@@      @      @      @       @      =@      @     �B@      2@      C@      @      8@      *@       @     �A@      @     �A@              0@              I@      @              �?      �?      1@      "@      9@      1@      >@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�o�\hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@��&Hz�@�	           ��@       	                    �?�R5���@�           ��@                           @{���]@�           ��@                            �?*�j��*@           P�@������������������������       ��.
�@�            `n@������������������������       ���LZ\@z           ��@                           @+�(B:@�            �m@������������������������       �FOQWn�
@Y             d@������������������������       �/�7&�Z	@0            @S@
                            �?�(^/�@6           8�@                          �2@}w�ni�@�            @x@������������������������       �|m��ۊ	@j            `d@������������������������       ��$d��@�             l@                          �3@L5izz�@=           P�@������������������������       �U���R�@=            @������������������������       ��"���@            �y@                           @m̝⥫@�           �@                           �?]�? g�@�           ��@                            �?�%S�U�@           �z@������������������������       ���K��@�            �l@������������������������       �#D�
@s            @i@                            @��nR@�           ��@������������������������       �DPNQع@           @z@������������������������       �b��̅@�            �j@                          �;@��0"Sc@(           �}@                           �?1����@�            Pt@������������������������       ���6"@e            `c@������������������������       �>��WG�@b            @e@                           �?J���
@a             c@������������������������       �SM��@            �F@������������������������       ��R��;�@F            �Z@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �d@     �U@     �v@     �E@     �|@      @     �h@      <@     �z@     �U@     �P@     �C@     �M@     �m@     �Q@     `x@     u@     `{@      V@      f@     �R@      G@      l@      6@     pu@       @      ]@      2@     �q@      C@      E@      0@      0@     �_@      @@     p@      h@     `r@      K@     @U@      9@      2@     �T@      &@     @f@      �?     �G@             �`@      (@      4@      @      @      K@      @     @]@     �Y@      d@      6@      J@      0@      .@     �M@      &@     `b@      �?      B@             @]@      $@      ,@      @      @      G@      @     @S@     �P@      b@      1@      .@      @       @      0@             �A@      �?      (@             �G@      @       @      @              (@              8@       @      @@       @     �B@      $@      @     �E@      &@      \@              8@             �Q@      @      @              @      A@      @     �J@     �M@     @\@      "@     �@@      "@      @      7@              ?@              &@              0@       @      @                       @              D@     �A@      0@      @      2@      "@       @      5@              2@              @              &@       @       @                      @              =@      :@       @      @      .@              �?       @              *@              @              @              @                      @              &@      "@       @             �V@      I@      <@     �a@      &@     �d@      �?     @Q@      2@     �b@      :@      6@      $@      *@      R@      =@     �a@     �V@     �`@      @@      8@      *@      $@      L@              K@              2@       @      I@       @      @      @       @      3@      @      7@      6@     �K@      @      (@      @       @      @@              A@              @              1@      @      �?      @      �?      �?              $@       @      >@      �?      (@      "@       @      8@              4@              .@       @     �@@      @      @      @      �?      2@      @      *@      ,@      9@      @     �P@     �B@      2@     �U@      &@     �[@      �?     �I@      $@     @Y@      2@      .@      @      &@     �J@      7@     @]@      Q@     �S@      :@     �B@      0@      &@      E@      �?      Q@      �?      :@      @      J@      ,@      &@      �?      �?      B@      0@      L@      D@      L@      @      >@      5@      @     �F@      $@     �E@              9@      @     �H@      @      @       @      $@      1@      @     �N@      <@      6@      3@     `c@     @V@      D@      a@      5@     @\@      @     �T@      $@     �a@      H@      8@      7@     �E@      \@     �C@     �`@      b@      b@      A@      X@     �L@      B@     @W@      &@     �X@      @     �M@      "@     @W@      C@      4@      1@      <@     @S@      4@     @V@      Y@     �U@      =@     �C@      (@      $@      B@       @      J@      @     �@@      @      I@      2@      @      @      @      6@       @      ?@      I@      ?@      *@      6@      @      @      .@       @     �C@              (@      �?      D@      "@       @      @       @       @      �?      7@      3@      1@              1@      @      @      5@              *@      @      5@      @      $@      "@      @      @      �?      ,@      @       @      ?@      ,@      *@     �L@     �F@      :@     �L@      "@      G@       @      :@      @     �E@      4@      .@      &@      9@     �K@      (@      M@      I@      L@      0@     �E@      A@      *@     �A@       @     �B@              .@              A@       @      &@      @      $@     �B@      @     �E@      A@     �E@      @      ,@      &@      *@      6@      @      "@       @      &@      @      "@      (@      @      @      .@      2@      @      .@      0@      *@      "@     �M@      @@      @     �E@      $@      .@              8@      �?     �H@      $@      @      @      .@     �A@      3@      F@     �F@     �L@      @     �E@      9@      �?     �A@      @      &@              $@      �?      B@      @      @      @      $@      <@      ,@     �@@      9@      ?@      �?      ,@       @              3@      @      $@              @      �?      8@               @              @      &@      @      1@      $@      0@      �?      =@      1@      �?      0@              �?              @              (@      @      �?      @      @      1@      $@      0@      .@      .@              0@      @      @       @      @      @              ,@              *@      @      �?       @      @      @      @      &@      4@      :@      @       @      @                       @                      @              �?      �?               @      �?              @      @      @      @      �?       @      @      @       @      �?      @              $@              (@       @      �?              @      @              @      ,@      4@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�
hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @$e�邛@�	           ��@       	                    @H]oS@           �@                            �?��ZV�@:           p�@                          �4@,)����@�           X�@������������������������       �ČY��@�             s@������������������������       ����ע@#           �{@                            �?ij@jBx@V           ��@������������������������       �����$�@�           H�@������������������������       �J`��W@�            �r@
                          �2@�32��@�           ��@                            �?%�
���	@           �z@������������������������       �7
�
@�            `r@������������������������       ��7�~1@O            @`@                           @.�h�f�@�            �@������������������������       �@���@�            @t@������������������������       �n���m=@�            �w@                          �6@z��7�@�           �@                           @�J �z@�           P�@                           @���H�F@C           P@������������������������       �qvGM)�@�            Ps@������������������������       �¿W��b@{             h@                           �?�2��@B            @]@������������������������       ����7!�@$            �N@������������������������       �/a%��	@             L@                          �8@tg�E:@,           �}@                           @��� v@g            �e@������������������������       �;ʿ�X@\            @b@������������������������       ��~t�z @             ;@                           �?���� �@�            �r@������������������������       �\)�(�@@             Z@������������������������       �s�i��@�            �h@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@     @`@     @W@     �s@     �D@     �~@      @     �l@      8@     �|@     �Z@     �R@     �C@     �Q@      l@     �M@     �x@     �r@      {@     @S@     �l@     @W@     �M@      m@      7@     �w@       @     �c@      2@     `v@      O@     �K@      8@      E@     �c@      D@     r@      k@      u@      G@     @_@     �L@     �E@     �b@      3@     �e@       @      \@      @      k@      D@      D@      3@     �@@      Y@      @@     @e@      _@     @h@     �@@     �L@      9@      .@     �P@      &@     �R@       @     �M@      @     �W@      *@      *@      *@      7@     �G@      $@     �L@     �I@     �W@      1@      6@      @      "@     �B@      �?      F@              7@      �?     �E@      @      @      �?      @      .@       @      9@      0@      F@      "@     �A@      6@      @      >@      $@      ?@       @      B@       @      J@       @      $@      (@      4@      @@       @      @@     �A@      I@       @      Q@      @@      <@     �T@       @      Y@             �J@      @     �^@      ;@      ;@      @      $@     �J@      6@     @\@     @R@      Y@      0@     �G@      :@      6@     �K@       @     �M@              =@      @     @S@      6@      1@      @      @      C@      3@     �U@      F@      S@      (@      5@      @      @      <@      @     �D@              8@             �F@      @      $@              @      .@      @      :@      =@      8@      @     �Y@      B@      0@     �T@      @     �i@              G@      &@     �a@      6@      .@      @      "@     �L@       @     �]@      W@      b@      *@      2@      @      �?      9@       @     @Z@              8@              Q@      @      @       @              3@             �J@      9@      P@      @      1@      @              2@       @      K@              2@             �K@      @      @                      ,@              E@      1@     �D@       @      �?      �?      �?      @             �I@              @              *@                       @              @              &@       @      7@      �?     @U@      >@      .@     �L@       @      Y@              6@      &@     @R@      2@      $@      @      "@      C@       @     �P@     �P@      T@      $@      <@      "@      @      5@             �H@              .@      @      G@       @      @                      .@       @     �B@      <@     �H@      @     �L@      5@      "@      B@       @     �I@              @      @      ;@      $@      @      @      "@      7@      @      =@     �C@      ?@      @     �^@     �B@      A@      T@      2@     �\@       @     @R@      @     �X@     �F@      3@      .@      <@      Q@      3@     �Z@     @T@      X@      ?@      T@      5@      2@      E@      (@     @V@      �?     �A@             �O@      3@      $@      @      $@      C@      @      M@      E@      N@      *@      Q@      3@      1@     �@@      (@      R@      �?      9@             �H@      2@       @      @      @      9@      @      L@      A@      C@      (@     �H@      &@       @      2@      $@     �G@      �?      3@              ?@      "@       @       @      @      ,@      @      ;@      &@      @@       @      3@       @      "@      .@       @      9@              @              2@      "@      @      �?              &@      �?      =@      7@      @      @      (@       @      �?      "@              1@              $@              ,@      �?       @              @      *@               @       @      6@      �?      @       @              @              .@              @              @      �?                              @              �?      @      *@      �?      @              �?      @               @              @              &@               @              @      $@              �?      @      "@              E@      0@      0@      C@      @      9@      �?      C@      @      B@      :@      "@      (@      2@      >@      .@      H@     �C@      B@      2@      "@      @      @      $@      �?       @              ,@       @      5@      *@      @       @      @      $@       @      (@      8@      @      ,@      "@      @      @      @      �?       @              ,@       @      ,@      *@      @       @      @      $@       @      (@      ,@      @      $@                              @                                              @                               @                              $@      �?      @     �@@      &@      &@      <@      @      1@      �?      8@      @      .@      *@      @      $@      &@      4@      @      B@      .@      @@      @      0@      @       @      "@       @       @      �?      &@      �?      @      @              @      @      @      @      (@      @      "@      �?      1@      @      "@      3@      @      .@              *@      @       @      @      @      @      @      .@      @      8@      (@      7@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ\R#hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @5g˽4�@�	           ��@       	                    �?�3z:1@�           ��@                           �?�u����@]           ��@                           @(/��@�            `v@������������������������       �>Ǵ��@�            �t@������������������������       ����$�(@             8@                            �?Oު��@�           p�@������������������������       ���S�L@U           Ѐ@������������������������       �<���@2             U@
                            �?��w@�           ��@                          �3@�����@R           ̔@������������������������       ��5�@u           Ȃ@������������������������       ���nHZ'@�           І@                           @�;�}}?@B           @@������������������������       �n��)@           �z@������������������������       �M�p��	@2             S@                           �?�G(�@�           8�@                          �:@p)����@�           �@                           @XU�� {@W           ؀@������������������������       ���2�{@           y@������������������������       �'��)u@T            @a@                           �?�:ۈI@V             a@������������������������       �G����
@             4@������������������������       ��2��@H             ]@                           @>-���@           �z@                          �9@MR��M@�            q@������������������������       �ʝ˜�7@�             l@������������������������       ���ADr@             H@                           @Ϟ1�@\            @c@������������������������       �4�OAY@             ?@������������������������       ��[���j@J            �^@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �^@     @V@     0v@      >@     @~@      "@     �o@      =@     �}@     �[@     �S@     �@@     @P@     �m@     �M@     �v@     �q@      {@     �V@     `j@     @V@      N@     `o@      0@     `w@      @      d@      .@      w@     �S@      L@      5@      E@     �d@     �B@     �p@     �g@     �u@      N@     @R@      D@     �@@     @S@      $@     @T@      @     �S@      @     �Y@      ?@      ?@      @      9@      M@      .@     @U@     �T@     �Z@     �@@      =@      @      1@      0@      @     �C@      @     �A@              C@      @      @      @      $@      4@      @      >@      >@     �I@       @      2@      @      0@      0@       @      C@      @     �A@              @@      @      @      @      $@      4@      @      <@      =@      I@       @      &@              �?              �?      �?                              @                                                       @      �?      �?              F@     �@@      0@     �N@      @      E@      �?     �E@      @      P@      8@      8@      @      .@      C@      &@     �K@     �J@      L@      9@      B@      =@      0@      J@      @     �B@      �?      E@      @     �I@      8@      5@      @      *@      =@      &@      F@      G@      H@      6@       @      @              "@      �?      @              �?              *@              @               @      "@              &@      @       @      @     @a@     �H@      ;@     �e@      @     Pr@      �?     �T@       @     �p@     �G@      9@      .@      1@     @[@      6@     `f@      [@     �m@      ;@     @[@     �E@      3@     �^@      @     �g@              M@      @      j@      C@      1@      $@      .@     �Q@      3@     @^@     @T@     `f@      8@      =@      .@      @     �P@       @     �V@              >@      �?     �^@       @      @       @      @      :@       @     �L@      9@     �X@       @      T@      <@      ,@     �K@       @      Y@              <@       @     �U@      >@      ,@       @      (@      F@      &@      P@      L@      T@      0@      =@      @       @      J@       @     �Y@      �?      9@      @     �L@      "@       @      @       @     �C@      @      M@      ;@      M@      @      5@      @      @      I@       @     @U@              6@      @      H@      @      @      @             �C@      @      G@      5@     �H@      @       @              @       @              2@      �?      @              "@       @      �?               @                      (@      @      "@             �Y@      A@      =@      Z@      ,@     �[@      @      W@      ,@      [@      @@      6@      (@      7@     @Q@      6@      Y@     @W@      V@      ?@      O@      2@      :@      N@      (@     �N@      @     �L@      *@     �L@      8@      ,@      &@      2@      D@      @      P@      P@     �G@      2@     �F@      (@      0@     �E@      $@     �N@             �E@      &@     �I@      6@      &@      @      0@      >@      @     �L@      I@     �@@      2@      9@      @      ,@     �C@      "@      D@             �A@      $@      B@      2@      @      �?      (@      4@      @     �C@     �C@      <@      2@      4@      @       @      @      �?      5@               @      �?      .@      @      @      @      @      $@      �?      2@      &@      @              1@      @      $@      1@       @              @      ,@       @      @       @      @      @       @      $@      �?      @      ,@      ,@              �?      @       @       @                      @       @       @       @                              �?                      �?              �?              0@      @       @      .@       @                      (@              @       @      @      @      �?      $@      �?      @      ,@      *@              D@      0@      @      F@       @     �H@             �A@      �?     �I@       @       @      �?      @      =@      0@      B@      =@     �D@      *@      @@      $@      �?      4@       @     �@@              6@      �?      :@      @      @               @      2@      0@      >@      .@      6@      &@      :@      $@      �?      1@      �?      ;@              .@      �?      6@      @                              0@      &@      =@      ,@      4@       @      @                      @      �?      @              @              @              @               @       @      @      �?      �?       @      @       @      @       @      8@              0@              *@              9@      �?      @      �?      @      &@              @      ,@      3@       @      �?                      @               @                              $@      �?                              �?                      @      @              @      @       @      5@               @              *@              .@              @      �?      @      $@              @      &@      .@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��wlhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@��,�ܲ@�	           ��@       	                   �0@DwH��@~           ��@                            �?���@�             l@                           @4����@P             a@������������������������       ���:�/�@?            @Y@������������������������       �ڀ�Xw@            �A@                           @,��
@:             V@������������������������       �j`����
@)             O@������������������������       ����@             :@
                            @���"�@�           |�@                            �? >�c_@%           ��@������������������������       ��=�;�@�           �@������������������������       �K�{C}
@y            @f@                           �?�"
��@�            �t@������������������������       ��G�e�@i            `e@������������������������       �`I�Ho�@f             d@                           @	Qj<�`@A           ��@                          @A@��̎l@�           �@                            �?�@[�:�@�           ��@������������������������       �\~ɦ�@)            }@������������������������       �_{3R#�@�           P�@                           @*O
���@             ?@������������������������       ��8$��?             *@������������������������       �.Q���"@             2@                          �4@kX:&��@]           (�@                           �? �?P
@n            �e@������������������������       ��H*��@4            �S@������������������������       �3�e[G�
@:             X@                          �9@
Ғ�k0@�           ��@������������������������       ��j�D�O@]           ��@������������������������       ��%���@�            �l@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@      a@     �U@     �v@     �A@      |@      "@      n@      D@     �|@     �Z@      K@      >@     �Q@     @n@     @Q@     �w@      q@     P{@     �T@     �Y@      9@      ?@     �b@      @     @i@       @     @U@      @     `e@      :@      4@      @      *@     �U@      ,@     @a@     �W@     @j@      6@      3@      �?      @      5@             �F@       @      &@              ,@      @      �?              @      1@       @      2@      2@     �E@              .@                      0@              4@              "@              @              �?                      *@       @      (@      &@      @@              ,@                      @              2@              @               @              �?                       @       @      &@      @      <@              �?                      $@               @               @              @                                      @              �?      @      @              @      �?      @      @              9@       @       @              "@      @                      @      @              @      @      &@               @              @       @              .@       @       @              @       @                      @      @              @      @      &@               @      �?              @              $@                              @       @                              �?                      @                     �T@      8@      <@      `@      @     �c@             �R@      @     �c@      6@      3@      @       @     �Q@      (@      ^@     @S@     �d@      6@      E@      2@      1@     @W@       @      ^@              E@      @     @`@      &@      ,@      @      @     �H@      @     @V@      M@     ``@      2@      >@      0@      ,@     �S@      �?      U@              ;@      @      \@      &@      "@      @       @      E@      @      R@     �I@     �W@      1@      (@       @      @      .@      �?      B@              .@              2@              @      �?      �?      @              1@      @     �B@      �?     �D@      @      &@      B@       @     �B@              @@              ;@      &@      @              @      5@       @      ?@      3@      B@      @      .@      @      $@      2@       @      6@              .@              @      @      @              @      (@              4@      *@      0@      @      :@       @      �?      2@              .@              1@              5@      @      �?              �?      "@       @      &@      @      4@             �n@     �[@     �K@      k@      ?@      o@      @     `c@      A@     0r@      T@      A@      :@     �L@     `c@     �K@      n@      f@     `l@     �N@     �c@     �T@     �E@     �]@      5@     �`@      @     �\@      =@     �c@      J@      8@      4@     �B@      Y@     �E@     �`@     �X@     @_@     �E@      c@      S@      C@     @]@      5@     �`@      @     �[@      =@     �c@     �H@      5@      2@      B@      Y@     �E@     �`@     �X@     @_@     �E@     �E@      =@      $@     �B@      @      D@       @     �@@      (@     �E@       @       @       @      ,@     �J@      @      8@      >@      H@      (@     �[@     �G@      <@      T@      0@     �W@      @     �S@      1@     �\@     �D@      *@      $@      6@     �G@      B@     �[@      Q@     @S@      ?@      @      @      @       @                              @              �?      @      @       @      �?                                                              @      @                                      �?                              �?      �?                                                              @       @               @                               @              �?      @       @      �?      �?                                                      V@      <@      (@     @X@      $@     �\@       @     �D@      @     �`@      <@      $@      @      4@     �K@      (@     �Z@     �S@     �Y@      2@      (@       @      �?      @              =@               @       @      <@      @               @              &@              ,@      7@     �@@       @      @      �?              �?              1@               @              @      @              �?              @               @      *@      7@              @      �?      �?      @              (@              @       @      5@      �?              �?              @              (@      $@      $@       @      S@      :@      &@     @W@      $@     @U@       @     �@@      @      Z@      8@      $@      @      4@      F@      (@      W@      L@     @Q@      0@     �M@      7@      @     @Q@       @     �N@              8@       @     @T@      .@      @      �?      *@      B@      @     �Q@     �D@      A@      $@      1@      @      @      8@       @      8@       @      "@      �?      7@      "@      @      @      @       @      @      6@      .@     �A@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�|PUhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�.�@�	           ��@       	                    @�VZ	@n           P�@                           �?�f��Z@           ��@                           �?5�M��@�            Ps@������������������������       �h�×>�@b            `d@������������������������       ��"[��@[            @b@                            �?y�ټ�@Y           ��@������������������������       ���g ��@r            �d@������������������������       �����@�            pw@
                           �?v&�4�R@X           �@                          �1@3b��:
@�            `w@������������������������       ������r@]            �c@������������������������       �aw�6�I
@�             k@                           @p�VX@t           X�@������������������������       �NJ��
@�            s@������������������������       ���0�*4@�            �q@                          �<@H��f"�@P           j�@                          �5@Ya^)@u           ��@                            �?����@�            �s@������������������������       ���Vͧ�@8             U@������������������������       ������O@�            �l@                           �?մ]F�>@�           ��@������������������������       ���ݢ�@�            �@������������������������       �F�[f;@�           (�@                           �??�M��N@�            @u@                           @�=�o�@�            �g@������������������������       ��IeU�@J            @[@������������������������       ��Z��(�@6            �T@                          �>@�z�P�N@[            �b@������������������������       ���v<��@0             T@������������������������       �*�Xr�
@+            @Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       @t@     �Z@     �R@     �t@      C@     �~@      (@      m@      ?@     �|@     �Z@      N@     �F@     @Q@     `m@      P@      w@     `t@     �{@     @W@     @`@      3@      5@     �c@      $@      q@       @      Z@      @     �o@     �B@      ?@      &@      0@     �Z@      7@     @d@      d@      o@      E@      Q@       @      ,@     @Q@      "@      [@       @     �G@      @     �W@      :@      1@      @      *@     �K@      1@     �R@     �U@      Y@      @@      5@      @       @      7@      @     �B@              4@      �?      F@      @      @      @              :@       @      4@      >@     �H@       @       @              �?      "@              7@              .@              :@      @       @      @              &@              "@      1@      :@      @      *@      @      �?      ,@      @      ,@              @      �?      2@       @      @                      .@       @      &@      *@      7@       @     �G@      @      (@      G@      @     �Q@       @      ;@       @      I@      3@      $@       @      *@      =@      .@     �K@     �L@     �I@      8@      @              @      ,@              >@              $@              0@      @      @       @      �?       @      @      .@      *@      9@      ,@      E@      @      "@      @@      @     �D@       @      1@       @      A@      .@      @              (@      5@      &@      D@      F@      :@      $@      O@      &@      @      V@      �?     �d@             �L@      @      d@      &@      ,@      @      @     �I@      @     �U@     �R@     �b@      $@      @@                      A@      �?     �S@              9@      @      H@      @                      @      :@       @      ?@      =@      L@      @      @                      @      �?      C@              @              ;@                               @      *@       @      ,@      .@      <@      �?      :@                      <@              D@              5@      @      5@      @                      �?      *@              1@      ,@      <@       @      >@      &@      @      K@             �U@              @@              \@       @      ,@      @              9@      @      L@     �F@      W@      @      &@      @       @      D@             �F@              2@             �K@      �?      &@       @              &@      @      ;@      2@      J@      @      3@      @      @      ,@             �D@              ,@             �L@      @      @       @              ,@              =@      ;@      D@      @     @h@      V@     �J@     �e@      <@      k@      $@      `@      9@      j@     @Q@      =@      A@     �J@      `@     �D@     �i@     �d@     �h@     �I@      e@      P@     �A@     �c@      6@     �g@      @      \@      8@      g@     �H@      8@      0@      C@     �[@      =@     �f@     ``@     �e@      H@      :@      0@              =@             �A@              5@      @      ?@      @      &@      @      @      0@      �?      F@      8@      >@      @      @      "@              &@              @              @      @      @              @      @      @      @      �?      @      @       @       @      7@      @              2@              >@              0@              9@      @      @      �?      @      (@             �B@      2@      6@      @     �a@      H@     �A@     �_@      6@     �c@      @     �V@      3@     @c@      E@      *@      (@      @@     �W@      <@      a@     �Z@     �a@      E@      K@      9@      =@     �L@      (@      O@      @     �L@      @      Q@      4@      @      @      6@     �C@      1@     @P@      L@     �S@      3@     @V@      7@      @     �Q@      $@     �W@              A@      (@     �U@      6@      @      @      $@     �K@      &@     �Q@     �I@     �O@      7@      9@      8@      2@      2@      @      :@      @      1@      �?      8@      4@      @      2@      .@      3@      (@      :@      A@      9@      @      &@      5@      $@      0@      �?      $@      �?      *@      �?      (@      @      @      ,@      @      $@       @      $@      8@      &@              @      *@      "@      @      �?      @      �?      @      �?      @      @      @      @      @      @      @       @      (@      @              @       @      �?      *@              @              @              @      �?       @       @              @       @       @      (@      @              ,@      @       @       @      @      0@      @      @              (@      ,@              @       @      "@      @      0@      $@      ,@      @       @      @      @      �?      @      @              @               @      (@              @      @      @      @      @      "@       @      @      @              @      �?      �?      (@      @                      @       @                      @      @      �?      *@      �?      (@        �t�bub�s     hhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ/n:phG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?,d;�]�@�	           ��@       	                    �?\<��@           ܙ@                          �5@��Ǎ�@^           �@                           �?�~Y�@�            @q@������������������������       ��X��@M             _@������������������������       ��&q& �@]             c@                           @}Q�a�@�            �p@������������������������       ��d��@~            `g@������������������������       �+�)��>@6            �S@
                           �?�S�?q@�           h�@                            @ĔT'A@�            Px@������������������������       �=B^_>�@|            �i@������������������������       � ��eQ�@s            �f@                           @����,@�           ��@������������������������       �.�m(@�            @y@������������������������       �*oY��@�            t@                          �3@�6/�n@�           ��@                           �?$��W�@n           ��@                           @;y�5i@S           Ѐ@������������������������       ���0�,q
@           �{@������������������������       �Ŵ�yi
@;             X@                           @�Ft�@           @z@������������������������       �}�kw�
@m            �d@������������������������       ��"���@�             p@                          �;@��e!�1@A           P�@                           @�gz�W�@�           ��@������������������������       ��U`,5@�           X�@������������������������       ��X\���@            |@                           @D�H|#�@l             e@������������������������       �jI]�;@8            �U@������������������������       ����'v@4            �T@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       pr@     �b@     @X@     Pv@      B@     P~@      (@      m@      ?@     Pz@     �Y@      P@      E@     �N@     �m@     @S@     �w@     ps@     �|@     @Q@     �[@      U@     �M@      c@      <@     @a@      $@     �^@      5@      c@      D@      ?@      =@     �C@     @Z@     �E@      b@     �`@     �e@     �B@      C@      3@      4@     �I@      �?     �P@      @      =@      �?     �F@      4@       @      @      "@      =@      2@     �F@      D@     �R@      0@      >@       @       @      @@      �?      >@              *@              ;@      @                      �?      (@      &@      7@      :@      C@      "@      0@      @      @      *@              (@              "@               @      @                      �?      @      �?      @      *@      5@      @      ,@      @      @      3@      �?      2@              @              3@       @                              @      $@      1@      *@      1@      @       @      &@      (@      3@              B@      @      0@      �?      2@      *@       @      @       @      1@      @      6@      ,@     �B@      @      @      @       @      ,@              9@      @      (@      �?      $@      *@       @      @      @      ,@      @      $@       @      7@      @      �?      @      @      @              &@              @               @                       @      @      @              (@      @      ,@             @R@     @P@     �C@     @Y@      ;@      R@      @     �W@      4@     �Z@      4@      7@      7@      >@      S@      9@     �X@     �W@     �X@      5@      8@      0@      2@      :@      @      <@              B@      @     �J@      @      (@       @      *@      A@      @      @@      A@     �@@      $@      *@      (@       @      ,@      @      $@              0@             �C@      @      $@       @      �?      1@      �?      5@      (@      3@      @      &@      @      $@      (@              2@              4@      @      ,@      @       @              (@      1@      @      &@      6@      ,@      @     �H@     �H@      5@     �R@      7@      F@      @      M@      0@      K@      ,@      &@      5@      1@      E@      5@     �P@     �N@     �P@      &@     �@@      <@      @     �C@      .@      9@      @      ;@      (@      7@      ,@       @      (@      &@      5@      @      E@     �E@      A@      @      0@      5@      ,@      B@       @      3@              ?@      @      ?@              "@      "@      @      5@      .@      9@      2@      @@      @      g@      P@      C@     �i@       @     �u@       @     �[@      $@     �p@     �O@     �@@      *@      6@     �`@      A@     @m@      f@     �q@      @@     �H@      4@      &@     @U@             �e@              O@              ]@      :@      *@       @      @      H@      (@     �Z@      K@     �d@       @      =@      $@      @     �I@             �X@              B@             �M@      @      "@      �?      @     �A@       @      J@     �@@     @Z@      @      5@      @      �?     �B@             �S@              >@             �J@      @      "@      �?      @      ;@       @     �H@      4@     @X@      @       @      @      @      ,@              4@              @              @                                       @              @      *@       @      �?      4@      $@      @      A@             �R@              :@             �L@      7@      @      �?      @      *@      $@     �K@      5@      O@      �?      @       @       @      1@              =@              @              3@      $@                       @      @      @      ?@      @      6@              *@       @      @      1@             �F@              4@              C@      *@      @      �?      �?      @      @      8@      1@      D@      �?     �`@      F@      ;@      ^@       @     �e@       @      H@      $@      c@     �B@      4@      &@      0@      U@      6@     �_@     �^@     �\@      8@      \@     �D@      .@     @]@      @     �d@              E@      $@     �`@      =@      3@      @      $@     �Q@      1@     �Z@     �\@     �W@      6@      S@      8@      @      Q@       @      \@              ?@             �W@      .@      @      �?      @      D@      @      M@      P@      P@      1@      B@      1@      "@     �H@       @      K@              &@      $@      D@      ,@      .@      @      @      ?@      ,@      H@      I@      >@      @      7@      @      (@      @      @      "@       @      @              2@       @      �?      @      @      *@      @      5@       @      5@       @      ,@      �?      @      @      @      @              @              &@      @               @       @      @      @      "@      @       @       @      "@       @      "@              �?      @       @                      @      @      �?       @      @      @              (@      @      3@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�j�KhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@ī����@�	           ��@       	                    @���P�k@�           ̕@                           �?1+�N@	           `�@                            �?'0 @            {@������������������������       �Pi�:@�            �i@������������������������       �H�g���@�            �l@                           �?;���@�            �w@������������������������       ���͗	@b             c@������������������������       ������@�            @l@
                            @��Y�S
@|           8�@                          �2@�\W�x+
@@           0~@������������������������       ��[>�	@           @y@������������������������       �`/���j	@5            �S@                           @�cg6@<             Y@������������������������       ���c�D�@&            @P@������������������������       �-H�.��@            �A@                          �;@\l #m@/           ��@                           @���A�@*           n�@                           @��7�-�@�           �@������������������������       ��S��@           ��@������������������������       ��2�a��@�           P�@                           @&/|/	@x             f@������������������������       ���@�A@]            @`@������������������������       �Q�T�_@             G@                           @�	��@           �y@                           �?t��>Q@�            �i@������������������������       �(_;��@5            �T@������������������������       �f��<p@T            �^@                            �?V.,�\@|            `j@������������������������       ��԰!@#             P@������������������������       �������@Y            `b@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        v@     �a@      Y@      u@      C@     �~@      @     �m@      :@     �|@     @\@      J@      >@     @Q@      i@      P@     pu@     Ps@     �|@      V@      [@      @@      7@      _@      @      k@      �?     �S@      @     @h@      ;@      1@      @      @     �O@      1@      a@      X@      l@      2@     �J@      3@      .@     �U@      @     �X@      �?     �B@      @      [@      :@      *@      �?      @      D@      .@     �T@     �N@     �_@      0@      @@      (@      (@     �E@      @     �J@      �?      9@      @     �B@      *@      "@      �?      @      7@      @      C@     �D@     @Q@      "@      (@      @      @      =@      �?      5@              $@      @      0@      @      @      �?              @       @      .@      1@      E@      @      4@       @      @      ,@      @      @@      �?      .@              5@      @      @              @      1@       @      7@      8@      ;@      @      5@      @      @     �E@             �F@              (@             �Q@      *@      @               @      1@      &@     �F@      4@     �L@      @      (@                      4@              ?@               @              :@      @      @              �?      @      �?      3@      @      4@      @      "@      @      @      7@              ,@              $@             �F@      $@      �?              �?      &@      $@      :@      0@     �B@      @     �K@      *@       @      C@      �?     �]@             �D@             �U@      �?      @      @              7@       @     �J@     �A@     �X@       @     �@@      &@      @      C@      �?     �Y@              ;@             @R@      �?      @      @              5@      �?      H@      ;@     �T@      �?      3@      @      @     �@@      �?     �U@              9@              P@      �?      @      @              0@      �?     �B@      :@      S@      �?      ,@      @      @      @              1@               @              "@              �?                      @              &@      �?      @              6@       @      �?                      0@              ,@              *@                                       @      �?      @       @      .@      �?      $@                                      .@              ,@              @                                                       @      @      &@      �?      (@       @      �?                      �?                               @                                       @      �?      @      �?      @             �n@     �[@     @S@     �j@      ?@      q@      @     �c@      7@     �p@     �U@     �A@      9@      P@      a@     �G@     �i@     �j@      m@     �Q@     �k@     @U@      H@     �g@      :@     @o@      @     �`@      5@      l@     �O@      @@      1@      G@     @]@     �@@     �e@     �f@     �f@      L@     �h@     �Q@     �G@      g@      6@     `m@      @     �^@      5@     @i@     �L@      <@      ,@     �D@     @X@      9@     �d@     @d@      f@      L@     �_@     �A@      =@     @Y@      "@     @f@      @     �U@      (@     �`@     �G@      3@      "@      8@     @P@      .@      [@     �[@      ^@     �E@     �Q@     �A@      2@      U@      *@     �L@             �A@      "@     �P@      $@      "@      @      1@      @@      $@      M@      J@      L@      *@      7@      .@      �?      @      @      .@              (@              6@      @      @      @      @      4@       @      "@      2@      @              5@      "@      �?      @      �?      *@              $@              1@      @      @              @      *@      @      @      &@       @               @      @                      @       @               @              @                      @              @       @      @      @      @              8@      9@      =@      6@      @      8@       @      9@       @     �D@      7@      @       @      2@      4@      ,@      @@     �@@     �I@      ,@      ,@      3@      2@      $@      @      ,@              @       @      ,@      &@      @      @      $@      &@      "@      8@      *@      *@      @      @      @      "@      @      �?       @              @       @       @      "@              �?      @      @      @      @      @      �?      �?      $@      .@      "@      @       @      @               @              @       @      @      @      @       @      @      1@       @      (@      @      $@      @      &@      (@       @      $@       @      3@              ;@      (@               @       @      "@      @       @      4@      C@      $@       @      �?      @      @               @              @                       @              �?      @      �?      @       @      ,@       @      @       @      @      @       @       @       @       @      ,@              ;@      $@              �?      @       @              @      @      >@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�{?hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @���k��@�	           ��@       	                   �4@�m�Ky@           6�@                            @Q@wj��@           �@                           �?�|�.��@;           ��@������������������������       �����>/@j           ��@������������������������       ���m�@�            @v@                           @	$��g@�            s@������������������������       ��*i�Y�@�             p@������������������������       �^�7�@"            �G@
                            @��-T��@           T�@                            �?����@*           h�@������������������������       �FZ�W@�            �@������������������������       �b���n@l             e@                          �:@!qh3.@�            �v@������������������������       ���c$ �@�             o@������������������������       �T�N�@=            �[@                           @��D��@�           ��@                           �?a���['@�           ��@                           �?��x��@�           P�@������������������������       ����O
@�             k@������������������������       �O�X"@            {@                          �1@�J�k@@>           �}@������������������������       ������6
@;            @Z@������������������������       �	>*Җ@           `w@                          �9@�� ��@�            Pt@                          �4@��j�j@�            Pq@������������������������       �hX���e
@`            �b@������������������������       �;>/ ��	@P            �_@                          �;@�Kw���@             H@������������������������       ����v��@             5@������������������������       ����v�	@             ;@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        r@      ^@     �U@     �v@      B@     `|@      "@     �n@      >@     �~@      [@     @Q@      C@     �S@     �n@     �P@     �w@     �r@     �z@     �T@      f@     @Q@     �N@     �j@      0@     �r@       @     �c@      5@     0u@     @R@     �@@      1@      G@     �c@      =@     �l@     �e@     `q@     �P@     �R@      3@      8@     �^@      "@      g@      �?     �P@      @     �f@      4@      &@      @       @     @R@      @     �\@     @V@      f@      >@     �I@      .@      .@     �X@      @     �a@             �D@      @     �b@      $@      "@      @      @     �O@      @     @T@     �O@     �a@      2@      :@      @       @      O@      @      X@              5@      �?     �R@      @      @       @      @      D@              I@      F@      Z@      "@      9@      $@      @     �B@             �F@              4@       @      S@      @      @       @              7@      @      ?@      3@     �C@      "@      7@      @      "@      7@      @     �E@      �?      9@      @      ?@      $@       @      @      @      $@      @      A@      :@     �@@      (@      7@      @       @      6@      @     �A@      �?      4@      @      4@      $@       @      @      �?       @      @     �@@      2@      ;@      &@                      �?      �?               @              @              &@                              @       @              �?       @      @      �?     �Y@      I@     �B@     �V@      @      \@      @     �V@      .@     �c@     �J@      6@      $@      C@     �T@      6@     �\@     �U@     �Y@     �B@     @T@      >@      4@      N@       @     �W@      @     �J@      @      `@     �A@      0@       @      2@     �N@      0@     �W@     �J@     �R@      7@      R@      =@      0@     �G@       @      P@      @     �G@      @     �U@      A@      @      @      0@     �G@      *@     �S@      G@     �P@      3@      "@      �?      @      *@              >@              @             �D@      �?      "@      �?       @      ,@      @      0@      @       @      @      5@      4@      1@      ?@      @      2@      �?     �B@      $@      >@      2@      @       @      4@      6@      @      5@     �@@      <@      ,@      0@      &@      @      1@       @      ,@              =@      $@      7@      ,@      @       @      0@      .@              1@      6@      3@      *@      @      "@      *@      ,@      @      @      �?       @              @      @      �?              @      @      @      @      &@      "@      �?      \@     �I@      :@     �b@      4@     �c@      �?      V@      "@     @c@     �A@      B@      5@     �@@      V@     �B@     �b@      _@     @b@      0@     �U@     �D@      4@     �]@      3@     �Y@              U@      @      ^@      A@      <@      1@      <@      J@     �B@      \@     �Y@     �Z@      ,@     �M@      8@      &@     �O@      .@      I@              I@      @     �O@      *@      1@      ,@      5@      >@      1@      L@     @Q@     �N@      (@      0@      $@      @      9@      �?      5@              (@              4@       @              @      @      *@      @      7@      <@      ;@      �?     �E@      ,@      @      C@      ,@      =@              C@      @     �E@      &@      1@      &@      2@      1@      $@     �@@     �D@      A@      &@      <@      1@      "@      L@      @     �J@              A@             �L@      5@      &@      @      @      6@      4@      L@     �@@      G@       @       @      @              .@              0@               @              &@      �?                              @              .@       @      ,@      �?      4@      (@      "@     �D@      @     �B@              :@              G@      4@      &@      @      @      3@      4@     �D@      9@      @@      �?      9@      $@      @      ?@      �?     �K@      �?      @      @      A@      �?       @      @      @      B@             �B@      6@     �C@       @      0@      $@      @      =@      �?      K@              @      �?      @@              @      �?      @      >@              B@      1@     �@@      �?       @      @       @      @              A@              @      �?      2@              @      �?              0@              4@      &@      4@      �?       @      @       @      9@      �?      4@                              ,@              �?              @      ,@              0@      @      *@              "@               @       @              �?      �?              @       @      �?      @      @      �?      @              �?      @      @      �?       @                      �?                                      @      �?              @      @              @                       @              �?      @               @      �?              �?      �?                      �?      �?                      �?       @              �?      @      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�OhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?Rd)���@�	           ��@       	                    �?N���S�@           ��@                          �:@��[s0@O           x�@                          �2@ѹ�!*k@           �z@������������������������       ��	���@S            `a@������������������������       ���k��@�            @r@                            �?أG�i@=             X@������������������������       �<CVA�@)             P@������������������������       �T���5@             @@
                            @*"L��@�           L�@                           @�@�i�]@�           @�@������������������������       �;�U�&�@�            �q@������������������������       ����w�@�            �v@                           �?����#�@+           �|@������������������������       �h���@L            @^@������������������������       ��+[�@�             u@                          �3@_�h`@�           Ρ@                           @t��u�_@g           ��@                           @L�bh�
@�           p�@������������������������       ��u�Y	@-           �|@������������������������       ����?�@�            0r@                            �?��9�X@�             m@������������������������       �N�#@�@X            �b@������������������������       ���7tF@2            �T@                           @�8t2\@X           @�@                          �5@�)C��@�           X�@������������������������       �<��WN@�            �n@������������������������       ��V���U@I           P@                           @���/�@d           (�@������������������������       ��_����@�            �r@������������������������       ��Q�B=@�            �n@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �`@     �U@     �t@      B@     �~@      (@     `g@      ?@     ~@     �Y@     �R@      E@      K@     �k@     �T@      w@     `t@     �{@     �S@      a@     �R@      N@     �`@      6@     �^@      "@     �T@      6@      d@     �I@      E@      3@     �A@     �V@     �G@     �c@     �a@     �g@      @@      A@      .@      8@      ;@       @     �J@              @@      @      N@      .@      *@      "@      @      A@      ,@     �N@      F@      O@      &@     �@@      &@      3@      3@      @      J@              =@       @     �K@      &@      "@       @      @      ;@       @      H@      ?@     �J@      "@      $@       @      @      @       @      .@              @       @      ,@                                      .@       @      (@      1@      <@      �?      7@      "@      (@      (@      @     �B@              8@             �D@      &@      "@       @      @      (@      @      B@      ,@      9@       @      �?      @      @       @      �?      �?              @       @      @      @      @      @      �?      @      @      *@      *@      "@       @      �?      @      @      @      �?                      �?              @      @              @              @      @      &@      @      @       @              �?      �?      @              �?               @       @                      @              �?      �?      @       @      @      @             �Y@      N@      B@      [@      ,@     @Q@      "@     �I@      2@      Y@      B@      =@      $@      <@     �L@     �@@     �X@     �X@      `@      5@      J@      C@      ,@     �P@      @     �F@      @      :@      .@     �P@      $@      1@      @      $@      C@      <@      I@      N@      U@      (@      7@      *@      @      =@      �?      :@      @      (@      &@      A@      @      @       @      @      $@      $@      ;@      ;@      6@      @      =@      9@      @      C@      @      3@              ,@      @     �@@      @      $@       @      @      <@      2@      7@     �@@      O@      @     �I@      6@      6@     �D@      "@      8@      @      9@      @     �@@      :@      (@      @      2@      3@      @      H@      C@     �F@      "@      3@      @      *@       @      �?      @      �?      @      @      $@      @      @               @      @       @      ,@      $@      &@      �?      @@      1@      "@     �@@       @      4@       @      5@              7@      7@       @      @      0@      *@      @      A@      <@      A@       @     �h@     �L@      :@      h@      ,@      w@      @      Z@      "@     t@      J@      @@      7@      3@     @`@     �A@     `j@      g@     �o@     �G@     �O@      1@      @     �W@      �?     �f@              L@       @     �d@      &@      (@      @      @      N@      (@     @S@      P@     �a@       @     �F@      @      @     �T@      �?     �b@             �D@              _@      @      @      �?      @      H@      $@     �P@      G@      Z@      @     �@@              @      H@      �?     �Y@              9@             @V@      @      �?      �?      �?      6@      @     �A@      4@     �P@      @      (@      @      @      A@             �G@              0@             �A@       @      @              @      :@      @      @@      :@      C@      �?      2@      *@              *@             �@@              .@       @      E@      @      @       @       @      (@       @      $@      2@     �B@      @      (@      "@              $@              .@              @       @      ?@      �?               @              @       @      $@      &@      =@       @      @      @              @              2@               @              &@      @      @               @      @                      @       @      �?     �`@      D@      4@     �X@      *@      g@      @      H@      @     `c@     �D@      4@      4@      *@     �Q@      7@     �`@      ^@     �\@     �C@     �T@      =@      &@     �N@       @      [@              C@      @     �U@      3@      &@      ,@      @     �C@      5@     @Q@     �L@      L@      <@      (@       @      @      <@              B@              &@              <@       @      $@      @              @      @      ;@      ;@      5@      ,@     �Q@      5@      @     �@@       @      R@              ;@      @      M@      1@      �?       @      @      A@      ,@      E@      >@     �A@      ,@     �I@      &@      "@     �B@      @     @S@      @      $@      @     @Q@      6@      "@      @      @      ?@       @     @P@     �O@      M@      &@      A@      &@      @      ,@             �I@              "@              B@      0@      @      @      @      ,@             �C@      <@      <@      @      1@              @      7@      @      :@      @      �?      @     �@@      @      @       @      @      1@       @      :@     �A@      >@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJYj�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@a>b�@�@�	           ��@       	                    �?�)V�P�@7           Z�@                           �?dn�t�@�           h�@                            @��@�            0q@������������������������       �o���!w@t            `f@������������������������       ���n�i@<             X@                           @0[��J@           �y@������������������������       ���rj@�            0p@������������������������       �a���@e            �b@
                          �2@T�u �@z            �@                           @)����@�           p�@������������������������       ���
@�            �r@������������������������       ��ʳ�$�@0           ~@                           �?'yy�=�@�           ��@������������������������       ���=���@�             o@������������������������       ���}��@�            �w@                           �?�7�來@�           p�@                           �?�����g@�           H�@                           �?��ol{&@�            0s@������������������������       �1z�i�@�            �o@������������������������       ��8�!�@$             J@                           �?����\J@�            `s@������������������������       �[���@c            �d@������������������������       ��0F�5@Z            @b@                          �6@[�&uw�@�           ̒@                           �?CqO�	@�            �i@������������������������       �-P���
@=            �Z@������������������������       ��;��R@E             Y@                            �?(�r[Ç@{            �@������������������������       ����w�@M           ��@������������������������       �n���@.           �|@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@      a@     �W@     �u@      B@     �~@      @     �l@      =@     �{@      \@     �R@      A@     �R@     �m@     @P@      x@     �p@      z@      T@     @g@      G@      B@     �h@      $@     �s@             �[@      @     �p@     �J@      J@      3@      7@     @^@      <@     �j@     �a@     �n@      >@     @R@      0@      6@     @Q@      "@      W@              C@      @     �M@      5@      1@               @      G@      @     �L@      P@     �Q@      0@      A@      @       @      >@      @      C@              "@      �?      2@      "@      �?               @      ,@      �?      ;@      7@     �C@      $@      4@      @      @      6@      @      =@              @              "@      @      �?               @      @      �?      2@      ,@      ;@      $@      ,@      �?      @       @       @      "@              @      �?      "@      @                              @              "@      "@      (@             �C@      $@      ,@     �C@      @      K@              =@      @     �D@      (@      0@              @      @@      @      >@     �D@      ?@      @      4@      @      @      =@      @      A@              2@       @     �@@      @      @              @      2@       @      2@      ;@      <@      @      3@      @      @      $@      �?      4@              &@      �?       @      @      *@              �?      ,@      �?      (@      ,@      @      @     @\@      >@      ,@     �_@      �?     �k@             @R@       @     �i@      @@     �A@      3@      .@     �R@      8@     �c@     @S@     �e@      ,@      N@      *@      @     �S@      �?     @^@              I@             @a@      "@      ,@      "@      $@      ?@      (@      V@     �@@     �Y@      @      7@       @      �?      A@              B@              @              P@      @      @              @      ,@       @     �H@      "@     �@@      @     �B@      &@      @     �F@      �?     @U@             �E@             �R@       @      "@      "@      @      1@      @     �C@      8@     @Q@       @     �J@      1@      @      H@             @Y@              7@       @     �P@      7@      5@      $@      @      F@      (@      Q@      F@      R@      "@      9@      @       @     �@@              F@              @      �?      ;@      &@       @              @      *@              5@      ,@     �B@      @      <@      ,@      @      .@             �L@              0@      �?      D@      (@      3@      $@       @      ?@      (@     �G@      >@     �A@      @     @d@     �V@      M@     �b@      :@     @f@      @      ^@      7@     �f@     �M@      7@      .@     �I@      ]@     �B@     �e@     �_@     �e@      I@      F@      3@      3@      A@      "@     �Q@      �?     �E@      @     �P@      =@      @      @      *@     �I@      &@      L@      K@     �J@      :@      .@      1@      "@      3@      @      9@      �?      7@      @      8@      2@      @      @      (@      6@      @      >@     �A@      3@      (@      &@      .@       @      1@      @      5@              5@      @      6@      2@       @      @      @      4@      @      =@      7@      0@      @      @       @      �?       @       @      @      �?       @       @       @               @              @       @              �?      (@      @      @      =@       @      $@      .@      @      G@              4@              E@      &@      @      �?      �?      =@      @      :@      3@      A@      ,@      1@      �?       @       @      @      5@              ,@              6@      "@      @      �?              ,@      @      *@      @      (@       @      (@      �?       @      @      �?      9@              @              4@       @                      �?      .@              *@      *@      6@      @     �]@     �Q@     �C@     @]@      1@     �Z@      @     @S@      1@     @]@      >@      0@      $@      C@     @P@      :@     @]@     @R@     �]@      8@      5@      @      &@      .@      @      D@              *@      @      8@      @       @       @       @      "@      @      6@      "@      $@       @      .@              @      @      @      =@                      @      0@      @      �?              �?      @      @      @      @       @              @      @       @       @      �?      &@              *@      �?       @      �?      �?       @      �?      @      �?      .@      @       @       @     @X@      Q@      <@     �Y@      (@     �P@      @      P@      (@     @W@      8@      ,@       @      B@      L@      4@     �W@      P@     @[@      6@      L@      F@      *@      K@      @      F@      @      <@      @     �M@      ,@       @      �?      1@      ?@      (@      C@      D@      O@      @     �D@      8@      .@      H@      @      7@       @      B@      "@      A@      $@      @      @      3@      9@       @     �L@      8@     �G@      .@�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ���"hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@N��@�	           ��@       	                     �?����n:@c           ��@                           @E�.?T�@�            �@                           �?GQɾ+{@0           |@������������������������       ��>I� �@n             d@������������������������       �j����@�            r@                           @*E��	@W           �@������������������������       ���덵g	@Q            @_@������������������������       ���*��@           `x@
                           @�V�Wy@�           �@                          �2@��"@�            �w@������������������������       ��fzf��@�             k@������������������������       ��%��@i            �d@                          �1@����j�
@�            Pv@������������������������       �ft�_7@Y            �a@������������������������       �T;O���	@�             k@                           �?g�Wl�@g           H�@                           @�)w<�@�           D�@                          �<@�.���@�           ��@������������������������       �m�M"�@D           �@������������������������       ��&$��c@E             Y@                          �;@ff8�,�@            {@������������������������       �W��)6h@�            �r@������������������������       ��%/S�@R            �`@                           @ΑwS�O@�           L�@                          �7@7�iX�X@H            �@������������������������       ��0��A@�            @n@������������������������       �ͯn�w@�            �r@                            �?�4v،�@�           ��@������������������������       ��p��P@�            v@������������������������       ��A�G6�@�             q@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@      b@     @T@     �v@     �D@     �}@      &@     @o@      <@      z@     �V@     �Q@     �A@      S@     �n@      P@     �v@     �s@     �{@      S@      \@     �@@      ?@     �d@      "@     �m@      �?     �Y@      "@      i@      ?@      >@      @      (@      Y@      9@     �c@     @a@     �p@     �@@      L@      6@      (@     �Z@      �?      ]@             �J@      "@     ``@      ,@      (@      @      @     �K@      1@     �U@     @S@     �c@      9@      ?@      @       @      L@              F@              :@      @      M@      &@      @              @      ;@      &@     �B@     �A@     �P@      .@      ,@      @              0@              1@              2@              4@      �?       @                      (@      @      "@      (@      ;@      @      1@      @       @      D@              ;@               @      @      C@      $@      @              @      .@      @      <@      7@     �C@      $@      9@      0@      @     �I@      �?      R@              ;@      @     @R@      @      @      @              <@      @      I@      E@      W@      $@      @      @              $@              .@              @              >@               @      �?              &@       @      .@              6@      @      6@      (@      @     �D@      �?     �L@              6@      @     �E@      @      @      @              1@      @     �A@      E@     �Q@      @      L@      &@      3@     �L@       @      ^@      �?     �H@             �Q@      1@      2@      �?      @     �F@       @      R@     �N@     �[@       @     �B@      $@      (@      6@       @      H@      �?      9@              A@      ,@      @      �?       @      <@      @      H@      <@     �E@      @      @      @      @      .@      @      9@      �?      (@              :@      "@      @      �?              3@      @      ;@      3@      ;@      @      >@      @      @      @      @      7@              *@               @      @      @               @      "@       @      5@      "@      0@       @      3@      �?      @     �A@              R@              8@              B@      @      &@              @      1@      @      8@     �@@     �P@      �?      @      �?      @      ,@              <@              $@              5@              @              @      @               @      (@      3@      �?      .@                      5@              F@              ,@              .@      @      @              �?      $@      @      0@      5@      H@             �i@      \@      I@     @i@      @@      n@      $@     �b@      3@     �j@      N@      D@      <@      P@     @b@     �C@      j@      f@     �e@     �E@      P@      M@      C@     �W@      3@      V@      @     �U@      ,@     �U@      :@      <@      3@     �G@     �J@      2@     �Z@     @V@     @T@      3@     �@@      =@      9@     �I@      &@     �P@      @     �L@      @      I@      7@      3@      "@      :@      5@      &@      M@     �F@     �H@      &@      9@      0@      .@     �G@      $@      N@      @      F@      @      F@      4@      3@      @      8@      1@      "@     �H@     �C@     �E@      &@       @      *@      $@      @      �?      @      �?      *@              @      @              @       @      @       @      "@      @      @              ?@      =@      *@      F@       @      5@              >@       @      B@      @      "@      $@      5@      @@      @      H@      F@      @@       @      ;@      *@      &@      @@       @      5@              3@       @      2@      �?       @      @      .@      6@      @     �D@      8@      2@       @      @      0@       @      (@                              &@              2@       @      �?      @      @      $@       @      @      4@      ,@      @     �a@      K@      (@     �Z@      *@      c@      @     �N@      @      `@      A@      (@      "@      1@     @W@      5@     �Y@      V@      W@      8@      N@      8@      @     �A@      @      T@              C@             �P@      &@      @      @      @     �K@       @     �G@      9@     �L@      .@      >@      &@      @      0@              C@              $@              8@      @              @       @      :@              ;@      @      =@      "@      >@      *@       @      3@      @      E@              <@              E@      @      @      �?       @      =@       @      4@      2@      <@      @     @T@      >@      @      R@      "@     @R@      @      7@      @     �O@      7@       @      @      *@      C@      *@     �K@     �O@     �A@      "@      I@      5@      @      C@      @     �@@              ,@              9@      2@      @       @       @      9@      @     �B@      A@      4@      @      ?@      "@       @      A@       @      D@      @      "@      @      C@      @       @      @      @      *@      @      2@      =@      .@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJt\BhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�I���@�	           ��@       	                   �4@X�,�@           �@                           �?KQ[�Y@g           �@                          �3@P��w�@r           ��@������������������������       �N0�]�@           �|@������������������������       ��l	)�>@V            �`@                            @mp�+=@�           В@������������������������       ��aJ�A�@`           8�@������������������������       �5I�6�T@�            �m@
                            �??6>�@�           8�@                           @��`�M�@o            @f@������������������������       �����[�@9            �W@������������������������       ��^D��@6            �T@                           �?�����@,           P}@������������������������       �uEFD�8@v            �e@������������������������       ��s����@�            `r@                           �?Ti5�@�           ��@                           @Ԗ�_!@�           0�@                          �?@8�ه�@�           0�@������������������������       ���r��@�           Ђ@������������������������       �����V�@.             S@                          �;@w�[:Ȇ@@             X@������������������������       �6-��]@$            �M@������������������������       �+ķ�K
@            �B@                          �7@B	��4@�           ��@                           @G��O�i@R            @_@������������������������       ����fg
@0            �R@������������������������       �?ؓ��u@"            �I@                           @,[�_7@l           ؁@������������������������       ���O��@�            �u@������������������������       ���4��@�            �k@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �_@     @U@      v@     �G@     �@      @     @k@      A@     @}@     �W@      M@     �F@     @Q@     �m@     �J@     pv@      u@     @y@     @V@     �i@     �M@      F@     `k@      9@     �x@             �_@      :@     �r@     �H@      C@      7@      8@     `a@      ;@     �l@     �h@     �p@     �G@     @c@     �B@     �A@      d@      3@     �p@             �W@      $@     �k@      =@      5@      0@      (@      [@      1@     �d@     �c@     @m@      C@      L@       @      5@     �J@      2@     @Q@             �A@       @     �H@      2@      "@      @      @      A@       @      E@     �N@     @S@      7@      D@      @      ,@     �F@      "@     �K@              :@      @      B@      *@       @      @      @      9@              >@     �L@     @Q@      .@      0@      �?      @       @      "@      ,@              "@      @      *@      @      �?      �?      �?      "@       @      (@      @       @       @     �X@      =@      ,@     �Z@      �?      i@             �M@       @     `e@      &@      (@      (@      @     �R@      .@      _@     �W@     �c@      .@     @Q@      9@      "@     �U@              d@             �H@       @      a@      "@      $@      (@      @     @P@      @      [@     @R@     �`@      $@      =@      @      @      4@      �?     �D@              $@              A@       @       @               @      "@      $@      0@      6@      9@      @      I@      6@      "@     �M@      @      `@             �@@      0@     @S@      4@      1@      @      (@      ?@      $@     @P@      D@     �A@      "@      *@      &@       @      9@              :@              @      &@      &@      @      "@      @      @      @      @      $@      *@      2@      �?      "@       @       @      4@              1@               @      @      @      @      �?      @      @       @      �?      @              &@              @      "@              @              "@              �?      @      @               @      �?       @      @      @      @      *@      @      �?     �B@      &@      @      A@      @     �Y@              >@      @     �P@      1@       @       @      @      8@      @     �K@      ;@      1@       @      *@      @      @      "@      @     �@@              0@              8@      @      @              @      @      @      >@      &@      @              8@      @      @      9@      @     �Q@              ,@      @      E@      (@      @       @      @      3@              9@      0@      (@       @     �\@      Q@     �D@     �`@      6@      \@      @     �V@       @     `e@     �F@      4@      6@     �F@      Y@      :@      `@     �a@     �`@      E@      H@     �C@      >@     �Q@      *@      B@      @     �N@       @      R@      8@      1@      &@      9@     �L@      0@     �P@     �R@     �Q@      >@      F@      9@      :@     @P@      @      =@      @      M@      @     �P@      7@      ,@      "@      4@     �I@      *@     �N@     �P@      P@      >@      C@      0@      2@     �O@      @      9@      @     �J@      @      O@      7@      ,@      @      2@     �H@      "@     �L@     �H@      O@      :@      @      "@       @       @              @              @              @                      @       @       @      @      @      1@       @      @      @      ,@      @      @      $@      @              @       @      @      �?      @       @      @      @      @      @       @      @              @      "@      @              @      @               @       @      @              @              @      @      @      @       @                              @              @      @       @              �?               @      �?               @              �?               @      @      @             �P@      =@      &@     �O@      "@      S@      �?      >@             �X@      5@      @      &@      4@     �E@      $@     �N@     �P@      P@      (@      3@      @      @      2@              (@              �?              *@      @                               @       @      "@      5@       @      @      1@      @      @      @              &@              �?              @       @                               @              @      (@      @      @       @       @      �?      *@              �?                              $@      @                                       @      @      "@      @      �?      H@      8@      @     �F@      "@      P@      �?      =@             �U@      0@      @      &@      4@     �D@       @      J@     �F@      L@      @      7@      $@       @      >@      "@      G@              :@              N@      ,@       @      @      $@      7@      @      9@      =@      :@      @      9@      ,@      @      .@              2@      �?      @              :@       @      �?      @      $@      2@      @      ;@      0@      >@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?@�0�e�@�	           ��@       	                    �?�/�i(@�           ��@                          �:@Gg���@r            �@                           �?|m�˳.@3            ~@������������������������       ��8���@           �z@������������������������       �#6�
�e@"            �K@                            �?����@?             Y@������������������������       ���B�@$            �N@������������������������       �֤�$^@            �C@
                           �?�_uz+p@            �@                          �3@l_r��X@�           p�@������������������������       �|�w��~
@�            �v@������������������������       ������@�            �y@                           �?t�����	@5            �U@������������������������       ���鴄@             8@������������������������       �vu���p@$             O@                          �6@ZC,�%@           B�@                            �?	��!N@�           �@                           �?�V��%@           ��@������������������������       �{�IZ�@�            @u@������������������������       �"
4�{�@3           �}@                           @��Tr��@�           `�@������������������������       ��j��M@m           ��@������������������������       ���ҋF
@6             V@                          �?@G}z�C�@m           (�@                           �?�$�S�@1           (�@������������������������       �ר��V�@�             u@������������������������       �[&�4��@d           ��@                            �?Zkv�M@<             X@������������������������       �����@             @@������������������������       ��XS�R�@*             P@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@     `b@      [@     �u@      B@      |@      @     �m@      B@     �z@      [@     @R@     �C@     �N@     �l@     @Q@     �v@     @r@     @|@      T@      _@      ?@     �D@      `@      $@     �i@      �?     @U@      @     �d@      D@      :@      0@      9@     �R@      ,@      a@      Y@     �f@      D@      G@      4@      =@     �H@      @      M@      �?     �B@      @      J@      9@      1@      ,@      1@      >@      @      H@      H@      N@      ,@     �E@      1@      :@     �B@      @     �L@      �?      B@      @      H@      .@      *@      @      .@      7@      @     �E@      ?@     �H@      (@      D@      .@      6@      >@      @     �G@             �A@      @     �G@      .@      "@      @      $@      6@      @      D@      7@      G@      $@      @       @      @      @              $@      �?      �?              �?              @              @      �?              @       @      @       @      @      @      @      (@       @      �?              �?              @      $@      @      &@       @      @       @      @      1@      &@       @      �?      �?       @       @       @      �?                              @      $@      �?      &@              @              @      @       @       @       @       @      �?      @                              �?                              @               @      �?       @      �?      &@      "@             �S@      &@      (@     �S@      @     `b@              H@      �?     @\@      .@      "@       @       @     �F@      "@      V@      J@     @^@      :@      S@      $@      &@      Q@      @      `@             �G@      �?     @Y@      ,@      @               @     �E@      "@     @T@      E@      [@      :@      :@      @      @      C@       @     @S@              ;@      �?     �F@      �?      @                      4@      @      B@      &@     �O@       @      I@      @      @      >@       @      J@              4@              L@      *@                       @      7@       @     �F@      ?@     �F@      8@       @      �?      �?      &@              2@              �?              (@      �?      @       @               @              @      $@      *@                                      �?               @              �?              @      �?      @                                      @              @               @      �?      �?      $@              0@                              @               @       @               @               @      $@      @              l@      ]@     �P@      k@      :@     `n@      @     @c@      ?@     �p@      Q@     �G@      7@      B@      c@     �K@     �l@      h@     �p@      D@     �\@      H@      A@      _@      1@      g@       @     �T@      ,@     `f@     �E@      8@      (@      ,@     �T@      ;@      b@     �_@     `f@      0@     �O@      =@      5@     @P@      �?     �W@              A@      $@      Z@      8@      *@      (@      @      F@      2@     @R@     �R@     �]@      *@      <@      ,@      *@      7@             �C@              ,@              J@      &@      @      &@      @      8@      @      @@      8@      D@      @     �A@      .@       @      E@      �?     �K@              4@      $@      J@      *@      "@      �?      @      4@      *@     �D@      I@     �S@      $@     �I@      3@      *@     �M@      0@     �V@       @      H@      @     �R@      3@      &@               @     �C@      "@      R@     �J@     �N@      @      F@      1@      *@     �L@      ,@     @S@       @      E@      @     @Q@      1@      $@              @     �B@      @      F@      H@      K@       @      @       @               @       @      *@              @              @       @      �?              �?       @      @      <@      @      @      �?     �[@      Q@     �@@     @W@      "@     �M@      @      R@      1@     �U@      9@      7@      &@      6@     �Q@      <@     �U@     @P@      W@      8@     �X@     �K@      >@      V@      "@      L@       @     �M@      1@     �T@      8@      5@       @      4@      Q@      5@      S@     �M@      U@      6@      G@      *@      ,@      E@       @      2@      �?      0@      .@     �B@      @      @      @      @      6@      @      9@      ;@     �@@      @     �J@      E@      0@      G@      @      C@      �?     �E@       @      G@      3@      1@      @      1@      G@      2@     �I@      @@     �I@      .@      &@      *@      @      @              @      �?      *@              @      �?       @      @       @       @      @      $@      @       @       @       @      @      �?      �?              @              (@                                      @                      @                       @              "@      "@       @      @                      �?      �?              @      �?       @               @       @      @      $@      @      @       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ`�jhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@G8���@�	           ��@       	                    �?�X�lPo@k           ��@                           @j�JH��@x           ��@                           �?��T��@`           ��@������������������������       �5�ےɎ@�             n@������������������������       ���CZ@�             t@                           �?�'#��C@            �B@������������������������       �.��Zz�?             ,@������������������������       ��Zf�Ke@             7@
                          �3@e��Y�]@�           d�@                            @~��I��@\           ��@������������������������       ����]�F@�           8�@������������������������       ��r���@s             g@                           @�n���@�            @o@������������������������       ������@O            �_@������������������������       �A��/@�
@H             _@                           �??}�%�@;           ��@                          �:@�+��)@           Ȋ@                           @���=�%@�           ��@������������������������       ��ހoJ�@�            �s@������������������������       �3s0���@�             u@                            �?)��P�@             i@������������������������       �s�����@K             ]@������������������������       �ˀ�[�W@4             U@                          �<@>���ɭ@"           �@                           @�x��y@�           �@������������������������       � K"��@S           0�@������������������������       ��0���e@V            �_@                            @��wl��@y            �g@������������������������       ���/�;Q@Q            �_@������������������������       �\�;���@(            �O@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       0r@     �a@      `@     �v@      D@     �}@      @     �k@      8@     �z@      [@      R@      G@      Q@     �l@      H@      v@     �u@      {@     @V@     �X@      A@      H@     �d@      (@     �n@      �?     �V@      @     `m@     �G@      >@      (@      "@     @[@      4@     �b@     @f@     �n@     �B@     �B@      (@      8@      P@      $@     �O@      �?      ?@      @     @Q@      1@      &@      @      @      E@      @      H@      L@     @P@      :@      ?@      "@      8@      N@      $@      O@      �?      ;@      @     �O@      1@      &@      @      @     �D@      @      D@     �J@     @P@      :@      "@      @      (@      >@      �?      <@              (@      �?      7@      @       @              @      ,@      @      1@      6@      A@      3@      6@      @      (@      >@      "@      A@      �?      .@      @      D@      $@      "@      @      @      ;@       @      7@      ?@      ?@      @      @      @              @              �?              @              @                              �?      �?               @      @                      @                      @                               @                                                                       @                                      @                              �?               @              @                              �?      �?              @      @                      O@      6@      8@      Y@       @     �f@              N@      �?     �d@      >@      3@      "@       @     �P@      .@     �Y@     �^@     `f@      &@     �G@      ,@      1@     �T@              c@             �K@             �a@      8@      ,@      @       @     �H@      "@     �V@     �S@     �a@       @     �A@      $@      $@     �P@             �`@             �C@              \@      ,@      *@      @       @     �C@      @     �S@      O@     @]@      @      (@      @      @      0@              4@              0@              <@      $@      �?                      $@      @      (@      1@      7@       @      .@       @      @      2@       @      >@              @      �?      :@      @      @      @              2@      @      *@     �E@     �C@      @      �?       @      @      @       @      (@              @              2@      �?      @      @              @      @      @      5@      6@       @      ,@              @      (@              2@              �?      �?       @      @       @      �?              *@              @      6@      1@      �?      h@     �Z@      T@      i@      <@     �l@      @     ``@      1@      h@     �N@      E@      A@     �M@     �^@      <@      i@      e@     �g@      J@     �V@      ?@      E@     �S@      1@      Z@      @     �F@      @     �U@      =@      $@      &@      ,@      I@       @      Q@      R@     �Q@      5@     �Q@      :@      ;@      Q@      @      X@      �?      B@      @     @R@      3@       @       @      $@     �B@      @      K@      K@     �G@      1@      ?@      2@      (@      9@      �?     �J@      �?      ;@             �D@      &@      @       @      @      @      �?      8@      5@      8@      ,@     �C@       @      .@     �E@       @     �E@              "@      @      @@       @      @              @      ?@      @      >@     �@@      7@      @      5@      @      .@      $@      ,@       @       @      "@       @      ,@      $@       @      "@      @      *@       @      ,@      2@      8@      @      0@       @      *@      @      @      @      �?      @       @       @      "@               @      @      @       @       @      @      *@              @      @       @      @       @      �?      �?      @              @      �?       @      @      �?      @              @      *@      &@      @     @Y@     �R@      C@     �^@      &@     �_@       @     �U@      (@     �Z@      @@      @@      7@     �F@      R@      4@     �`@      X@     �]@      ?@     @U@     �J@      9@      [@      $@     @\@       @     @S@      (@      X@      =@      ?@      &@     �A@     �N@      1@     �\@     �S@     �Z@      =@     �P@      G@      8@     �W@      $@      [@       @     @S@      (@     @U@      =@      ;@      $@      ?@     �I@      1@     @Y@      O@     �U@      ;@      2@      @      �?      ,@              @                              &@              @      �?      @      $@              ,@      0@      4@       @      0@      6@      *@      ,@      �?      *@              "@              $@      @      �?      (@      $@      &@      @      2@      2@      *@       @      $@      0@      @      "@              (@              "@              @      �?      �?      &@       @      @      �?      &@      @      &@      �?      @      @      @      @      �?      �?                              @       @              �?       @      @       @      @      (@       @      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ���3hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?~��\�@�	           ��@       	                   �:@[y��@           �@                           �?��ǈw�@,           ��@                            �?���G��@4           �@������������������������       �D����@d            �c@������������������������       ���Wu�@�            Pv@                           �?����F@�           p�@������������������������       ��~`�B@�            Pp@������������������������       ��<;6@Z           H�@
                           @	�X�O�@�            0u@                          �?@���v�@�             j@������������������������       ��O��F�@e             d@������������������������       �`b�Q@"            �H@                          �@@�B$��P@P            @`@������������������������       ���'��@G            @\@������������������������       �?�{]�X@	             1@                           �?8k	[@�           ��@                          �1@��X�@+           ��@                            �?�5�r	@~            @g@������������������������       �nE����@G            @X@������������������������       �GNRݬ@7            @V@                          �9@X}��j@�            �@������������������������       �E�C-*�@Z           �@������������������������       �l�Y�@S            @`@                           @�@���@l           ��@                           @eZ���@�           @�@������������������������       ���<c�@)           0}@������������������������       �Q@cf@�            Ps@                          �6@ֆ�P*T@{           �@������������������������       ��j��q�@�            y@������������������������       ��wr!@�             j@�t�b�/     h�h5h8K ��h:��R�(KKKK��h��B`       �t@      `@     @V@     u@      G@     �|@      $@     �k@     �B@     @|@      \@      P@      >@     �Q@     �p@     �P@     �w@      s@     0z@     �U@     @_@      P@      M@     �a@     �@@     �a@      "@     @^@      ?@      a@     �L@      B@      *@     �J@     @[@     �C@      c@     ``@     `e@      E@      Z@      D@      G@     �[@      <@      a@       @     �V@      ;@      ^@     �F@      =@      @      G@     @S@      ?@      `@     �Y@      _@      B@     �A@      &@      5@      O@      �?     �L@      �?      ?@      @      C@      5@      $@              1@      7@      2@     �E@      D@      Q@      (@      @      @      @      <@              ,@      �?      &@              "@      @       @               @      @      @      @      (@      @@       @      =@       @      2@      A@      �?     �E@              4@      @      =@      2@       @              "@      1@      ,@     �B@      <@      B@      @     @Q@      =@      9@      H@      ;@      T@      �?     �M@      7@     �T@      8@      3@      @      =@      K@      *@     �U@      O@      L@      8@      @@      @      @      (@      @     �@@              2@      @      7@      @      @      �?       @      1@      @     �A@      ,@      <@      "@     �B@      6@      5@      B@      4@     �G@      �?     �D@      4@     �M@      1@      *@      @      ;@     �B@      $@     �I@      H@      <@      .@      5@      8@      (@     �@@      @      @      @      ?@      @      0@      (@      @      "@      @      @@       @      8@      =@     �G@      @      ,@      4@      @      9@      @       @      @      2@      @      @      &@      @      @      @      7@      @      1@      ,@      1@      �?      "@      "@      @      8@      �?              @      1@      @      @      "@      @      @       @      2@      @      ,@      &@      .@      �?      @      &@      @      �?       @       @              �?                       @      �?       @       @      @      @      @      @       @              @      @      @       @       @      @              *@              &@      �?      �?      @      @      "@       @      @      .@      >@      @      @              @      @       @      �?              (@              &@              �?              @      "@       @      @      *@      >@      @              @       @      �?               @              �?                      �?              @                                       @                     @j@      P@      ?@     @h@      *@      t@      �?     @Y@      @     �s@     �K@      <@      1@      1@     `c@      <@     �k@     �e@      o@     �F@     �S@      *@      @      P@      "@     �c@             �D@      �?     �a@      5@      @       @       @     �O@      @     �Q@      O@     �W@      7@      @                      "@      @     �K@              @              =@      �?      @              �?      ,@              ,@      4@      4@      @      @                      @      @      6@              @              4@              �?                      ,@              @      @      $@      �?       @                      @      �?     �@@              �?              "@      �?       @              �?                      @      .@      $@       @      R@      *@      @     �K@      @     �Y@              A@      �?      \@      4@      @       @      �?     �H@      @     �L@      E@     �R@      4@     �M@      *@      @     �H@             �T@              >@      �?      V@      1@      �?       @      �?     �C@              J@     �@@      O@      &@      *@               @      @      @      4@              @              8@      @      @                      $@      @      @      "@      (@      "@     �`@     �I@      8@     @`@      @     @d@      �?      N@      @     �e@      A@      5@      .@      .@      W@      7@      c@     @\@     @c@      6@      R@      @@      0@      S@             �U@              E@      @     �X@      2@      ,@      @      $@     �F@      4@     @W@      O@     �Q@      $@     �B@      *@      "@     �H@              O@              ;@      �?      J@      @      *@      @      "@      8@      (@      L@      @@      K@      @     �A@      3@      @      ;@              9@              .@      @      G@      *@      �?      �?      �?      5@       @     �B@      >@      1@      @      N@      3@       @      K@      @     �R@      �?      2@      �?     @S@      0@      @      "@      @     �G@      @     �M@     �I@     �T@      (@     �A@      @      @      B@      �?     �O@              0@      �?     �N@      $@      @       @              ?@             �F@      >@      H@      @      9@      ,@       @      2@      @      (@      �?       @              0@      @       @      @      @      0@      @      ,@      5@     �A@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�vB5hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���J�@�	           ��@       	                   �:@�� �
@#           @�@                          �3@#���@O           ؔ@                            �?�0l�@)            }@������������������������       ��I�M�:@�             n@������������������������       ��U��@�             l@                           @���7'@&           0�@������������������������       �C"�j
@�           ��@������������������������       �Ba-���@8            �T@
                          �<@�<�ͯ�@�            �u@                           �?�L�W*@W            `c@������������������������       �,���7@             L@������������������������       ���3�@;            �X@                           �?�#r�@}            �g@������������������������       �x��/&@(            �N@������������������������       �}:����@U            @`@                           �?�	�G�u@�           r�@                           @;(���@�           Ȉ@                            �?��Z�]@u           ��@������������������������       �^ܧן;
@�            �w@������������������������       �/���@�            �k@                           �?�"�h@}             h@������������������������       �Ɲ�k�@C            �Y@������������������������       �-$1�
@:            �V@                            �?��0+R@�           ��@                           @��2�#@*           ؊@������������������������       ����W@�           ��@������������������������       �持f�@?            �X@                           @�IYo{@x           (�@������������������������       �������@�            `u@������������������������       ����@�            �m@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �r@     @_@     �W@     �v@     �F@     �}@      "@     `j@      C@     �z@      Z@     �Q@     �C@      Q@     �p@     �Q@     �w@     Ps@     �{@     �T@      `@      I@     @P@      d@      >@     �`@      "@     �W@      >@      a@     �J@      G@      7@      G@     �^@      ;@     �a@     `c@     �f@     �F@      [@      =@     �F@     @_@      9@     �_@      @      Q@      8@     �]@     �F@     �@@      &@     �C@     �Y@      4@     �]@      [@      b@     �D@      ?@      @      .@      E@       @     �M@      �?      2@      @      C@      .@      *@      �?      @      @@      @      E@     �G@     @R@      ,@      ,@       @      $@      8@              9@              @      @      8@      @      @      �?      @      3@      �?      .@      1@      I@      &@      1@      @      @      2@       @      A@      �?      (@              ,@       @      @              @      *@      @      ;@      >@      7@      @     @S@      8@      >@     �T@      7@     �P@      @      I@      3@     @T@      >@      4@      $@      @@     �Q@      0@      S@     �N@     �Q@      ;@     �P@      1@      <@     �S@      6@     �O@      @     �E@      1@      R@      >@      ,@       @      ?@     �N@      "@     @Q@      M@     �Q@      ;@      &@      @       @      @      �?      @              @       @      "@              @       @      �?      "@      @      @      @                      5@      5@      4@      B@      @       @      @      :@      @      2@       @      *@      (@      @      4@      @      7@     �G@     �C@      @      $@      @      @      2@      @      �?      @      0@      @      @      @      "@               @      @      �?      $@      5@      :@       @      @       @      @       @              �?      @      @       @      @      @      @                      @               @      @      ,@      �?      @      @       @      0@      @                      (@      �?      @              @               @       @      �?       @      2@      (@      �?      &@      .@      ,@      2@              @              $@      @      (@      @      @      (@      @      .@      @      *@      :@      *@       @      �?      �?      @      @              �?               @      @      @      @              @      @      "@      @      @      @      @              $@      ,@      &@      *@              @               @              @       @      @      @      �?      @      @      $@      6@      $@       @      e@     �R@      =@     @i@      .@     �u@             @]@       @      r@     �I@      8@      0@      6@     �a@     �E@     �m@     @c@     0p@      C@     �P@      .@      $@      N@      @     �_@              F@             �\@      (@      @              @      I@       @     �W@      K@     @[@      .@      H@      "@      @      F@      @     �[@              >@             �U@      "@      @              �?     �C@      @     �S@     �E@     �R@      "@      :@      "@       @      7@       @     �P@              3@             @P@      @                              9@      �?      H@      6@     �N@      @      6@               @      5@       @      F@              &@              6@      @      @              �?      ,@      @      >@      5@      ,@      @      3@      @      @      0@              1@              ,@              <@      @                      @      &@      �?      1@      &@      A@      @      "@      @       @      $@              ,@              @              .@      �?                       @      @              @      @      0@      @      $@              @      @              @               @              *@       @                       @      @      �?      &@      @      2@             @Y@      N@      3@     �a@      &@      k@             @R@       @     �e@     �C@      5@      0@      1@      W@     �A@     �a@      Y@     �b@      7@     �M@     �E@       @     �T@      @     �_@              A@      �?      X@     �@@      *@      *@      ,@     �O@      .@     �T@     �P@     @V@      .@     �G@      D@      @      T@      @     @\@              =@      �?     �V@      :@      (@      "@      ,@      I@      .@     @S@     �I@      S@      .@      (@      @      �?       @              *@              @              @      @      �?      @              *@              @      .@      *@              E@      1@      &@      N@      @     �V@             �C@      @     @S@      @       @      @      @      =@      4@     �N@      A@     �N@       @      ;@      &@      �?     �D@      @      K@             �A@      @      B@      @      @                      ,@      4@      E@      0@      6@      @      .@      @      $@      3@      �?     �B@              @      @     �D@      �?      @      @      @      .@              3@      2@     �C@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ]�3PhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@���2�@�	           ��@       	                   �4@kˏC��@�           ��@                           �?�^K�%V@_           ��@                           @�_Bh�@k           P�@������������������������       ��tM"�@�            �v@������������������������       �~��Z�@y            `g@                           @=\��@@�           P�@������������������������       ��񉉻S@�           P�@������������������������       �i���uv@X           P�@
                          �5@��o��|@s           x�@                           �?Y����a@�            Ps@������������������������       �;�e�T�@T             _@������������������������       ���|��@t             g@                            �?���m*c@�            �q@������������������������       ��e��	'@c            �c@������������������������       ��@Tpl@H            �^@                            @[eWs�@�           �@                            �?8��dpF@�           p�@                           @Z�+�-K@           �z@������������������������       �a�d��@�            Ps@������������������������       �sH��@Q            �^@                           �?_~(U+�@�           h�@������������������������       ��n�*8s@�             o@������������������������       �����EE@�            @w@                           �?�'�MB@1            ~@                          �7@�U�"�e@b            �b@������������������������       �b�����@             ;@������������������������       �w�`ħ+@R            �^@                           @-����@�            �t@������������������������       �7D�Y@�            @r@������������������������       ����7�M@            �C@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@     �`@     @V@     �u@      @@     `|@      @     @l@      7@     @z@     �Y@      N@     �D@     @R@     �o@     @T@     �w@     �t@      z@     �X@     �g@      Q@      H@     �l@      &@     �t@      �?     �`@      (@     r@      O@     �B@      "@      =@     �a@      ?@     �m@     �h@     0q@     �J@     �a@      A@     �@@     �e@      $@     �n@      �?      Y@      @     �k@     �F@      7@      @      1@     @Z@      8@     @f@     �d@     @l@      E@     �Q@      &@      5@     �H@       @      K@      �?      :@       @     �J@      1@      *@      �?      (@      C@      @     �E@     �H@      N@      3@     �G@      $@      *@      >@      �?     �D@      �?      (@      �?      F@       @      @      �?       @      6@      @      ?@      >@     �F@      &@      7@      �?       @      3@      @      *@              ,@      �?      "@      "@      "@              @      0@              (@      3@      .@       @     �Q@      7@      (@     @_@       @     �g@             �R@      �?      e@      <@      $@      @      @     �P@      1@     �`@     �\@     �d@      7@     �A@      3@      @     @W@      �?     �W@              :@             @T@      2@      @       @      @      =@      .@     �U@      O@     @V@      .@      B@      @      @      @@      �?     �W@              H@      �?     �U@      $@      @       @       @      C@       @      H@     �J@     @S@       @     �G@      A@      .@      L@      �?     @V@              @@      "@      Q@      1@      ,@      @      (@     �A@      @      M@     �@@     �H@      &@      =@      6@      @      >@             �@@              5@      @      8@      @      @      @       @      5@      �?      B@      <@      9@      @      ,@       @       @      *@              1@              $@      @       @                              @      @      �?      1@      (@      @      @      .@      ,@      @      1@              0@              &@              0@      @      @      @       @      2@              3@      0@      4@       @      2@      (@      $@      :@      �?      L@              &@      @      F@      (@      @              @      ,@      @      6@      @      8@      @      1@      @      $@      3@              @@              @      @      2@      �?      @              �?      @      @       @      @      5@      �?      �?      @              @      �?      8@              @       @      :@      &@      @              @      "@              ,@       @      @      @     `d@     �P@     �D@     �]@      5@     @^@      @     �W@      &@     ``@      D@      7@      @@      F@     @\@      I@     �a@     ``@     �a@      G@     �\@      G@      4@     �V@      &@     �W@      @     �N@       @      Z@      <@      ,@      4@      5@     �R@     �B@     �X@     @U@     �Y@      8@     �H@      8@      "@     �D@      "@      A@      @     �@@              =@      @      �?      (@      ,@      B@      (@      A@     �A@      D@      "@      9@      0@      @      :@      "@      2@      @      >@              7@      @      �?      (@      "@      ?@      "@      4@      ;@      ?@      "@      8@       @      @      .@              0@              @              @       @                      @      @      @      ,@       @      "@             @P@      6@      &@      I@       @      N@       @      <@       @     �R@      5@      *@       @      @     �C@      9@      P@      I@      O@      .@     �A@      @      @      *@       @      <@       @      0@       @      9@      (@       @      @      �?      0@       @      6@      1@      <@      $@      >@      2@       @     �B@              @@              (@              I@      "@      &@      @      @      7@      1@      E@     �@@      A@      @     �H@      4@      5@      <@      $@      ;@             �@@      "@      ;@      (@      "@      (@      7@      C@      *@      E@      G@     �C@      6@      0@      @      "@      @      @      @               @      @      (@      @      @       @      �?      @      @      *@      0@      4@      (@      �?      �?      @                      @              �?       @       @                                                              $@      @              .@      @      @      @      @      �?              @      @      $@      @      @       @      �?      @      @      *@      @      1@      (@     �@@      ,@      (@      6@      @      7@              9@      @      .@      "@      @      $@      6@      A@       @      =@      >@      3@      $@      <@      (@      (@      *@      @      7@              9@      @      &@      @      @      $@      6@      :@      @      :@      >@      1@      "@      @       @              "@                                              @      @                               @       @      @               @      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ;�khG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?��9P��@v	           ��@       	                   �?@�u�=��@�           ��@                            @��#��n@�           L�@                           �?D�^f�@            ��@������������������������       �K9ԓ�+@�            s@������������������������       ���M�@k           (�@                           @��)�@x           �@������������������������       �Ϭ8�$@�            @q@������������������������       ��ߨ���@�            �t@
                           �?��MCd@:            @V@������������������������       ��§�?@             2@                           @g�/���@/            �Q@������������������������       ��C�Y }@            �C@������������������������       �|R��>
@             @@                           @��4J�@�           :�@                           �? ���+@;           ܔ@                           @"o��Q@           �|@������������������������       �ߜQ�@�            �j@������������������������       �����@�            �n@                          �3@�_���&@            `�@������������������������       ��\�'@�            �t@������������������������       ��@���@Y            �@                           @�փ��@i           0�@                            �?�DR��
@            |@������������������������       ��f��X@?             Z@������������������������       ��BE른	@�            �u@                            @��Mv@T            �@������������������������       ��z�?z6@           �{@������������������������       �U �:��@F             Z@�t�bh�h5h8K ��h:��R�(KKKK��h��B        �r@      a@      Z@     pw@      H@     P}@      @     @n@      ;@     0z@      X@     �K@      A@      R@     Pp@     �T@     �u@     �r@     �}@      Q@      ^@     �P@     @P@      a@     �@@     ``@      @     �^@      6@     `b@     �E@      >@      0@     �D@     @[@      =@      \@      `@     �h@      =@     �[@      H@      M@     ``@      ?@     �_@      @     �\@      6@      b@     �E@      <@      $@      C@     �Z@      8@     @[@     @_@      h@      9@      L@      ?@      >@     �V@      ,@     @R@      �?      P@       @     �V@      0@      4@       @      3@      Q@      3@      P@      Q@      a@      .@      (@      $@      @      8@      @      =@              :@             �C@       @       @       @      @      4@      �?      1@      7@      P@      @      F@      5@      7@     �P@      &@      F@      �?      C@       @      J@       @      (@              *@      H@      2@     �G@     �F@      R@      "@     �K@      1@      <@      D@      1@      K@       @     �I@      ,@     �J@      ;@       @       @      3@     �C@      @     �F@     �L@      L@      $@      7@      "@      *@      9@      �?      :@             �@@      @      4@       @      @      �?      *@      .@      @      5@      >@      3@      @      @@       @      .@      .@      0@      <@       @      2@      "@     �@@      3@      @      @      @      8@      �?      8@      ;@     �B@      @      "@      2@      @      @       @      @               @              @               @      @      @       @      @      @      @      @      @                              �?              @              @                              �?              �?               @      �?              �?      @      "@      2@      @      @       @                      @              @              �?      @       @       @      @       @      @      @              �?      .@      @       @       @                      @              �?                              �?       @       @      �?      @                       @      @      �?       @                               @               @              �?      @      �?              �?      �?      �?      @             `f@     �Q@     �C@     �m@      .@      u@      �?     �]@      @      q@     �J@      9@      2@      ?@      c@     �J@     `m@      e@     �q@     �C@     �Z@     �F@      5@     �c@      ,@     �e@              P@      @     �c@     �A@      0@      $@      .@      U@      I@     ``@     @U@      a@      =@     �D@      @      @     �F@      @      O@              9@              N@       @      @       @      &@      A@      @     �M@      @@      C@      0@      ;@      �?       @      8@      �?      2@              (@              ?@      @      @       @              4@      @      ;@      ,@      ,@       @      ,@      @      @      5@      @      F@              *@              =@      @                      &@      ,@      �?      @@      2@      8@       @     �P@      D@      0@      \@      "@     @\@             �C@      @     @X@      ;@      "@       @      @      I@      G@      R@     �J@     �X@      *@      .@      &@      @     �I@              B@              *@              G@      @      �?                      8@      3@     �A@      &@      M@             �I@      =@      "@     �N@      "@     @S@              :@      @     �I@      6@       @       @      @      :@      ;@     �B@      E@      D@      *@      R@      :@      2@     �T@      �?     `d@      �?     �K@      �?     �\@      2@      "@       @      0@      Q@      @      Z@     �T@      b@      $@      ?@               @     �B@      �?     �W@              :@              L@      @      @      @       @      9@              C@      D@     �R@      @      (@              @      @              0@              @              0@      �?      @      �?       @      @              0@      @      $@              3@              @     �@@      �?     �S@              4@              D@      @       @       @              2@              6@     �A@      P@      @     �D@      :@      $@     �F@              Q@      �?      =@      �?     �M@      *@      @      @      ,@     �E@      @     �P@     �E@     �Q@      @      A@      4@      $@      =@              O@      �?      7@      �?     �G@      *@      �?      @      (@      ?@      @      M@      =@      O@      @      @      @              0@              @              @              (@              @               @      (@               @      ,@      "@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ� �UhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�p%j@�	           ��@       	                    @E�8h	@           H�@                           �?���b��@t           L�@                           �?��5��/@�           \�@������������������������       ���m�>@�            �v@������������������������       ���2q�L@�           P�@                          �6@4�<$+@�           ��@������������������������       �rJ�*�@*           �}@������������������������       ��1Ej^H@�            �q@
                           �?���c�2@�           D�@                          �2@�c���]@�            �w@������������������������       �ɒ�!'@              L@������������������������       ��e��Mf@�             t@                           �?Ґ@!Dk@�           Ȅ@������������������������       ��μOj@�            �r@������������������������       �o�ɝ�/@�            �v@                          �6@�v�p�	@�           ��@                          �5@bɥ��@�           �@                           �?�����@\           ��@������������������������       ��sIlB@�            @r@������������������������       ���cl׸@�            @o@                           �?k���@6            �W@������������������������       �o�Cs�4@            �B@������������������������       �p�I	J;
@!             M@                           �?IR���@           �z@                           @�@��@)            @P@������������������������       ��S��vH@            �E@������������������������       ���7��@             6@                           @H�$���@�            pv@������������������������       ���]��@�            �s@������������������������       ��J'P"@            �E@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �r@     �^@     @V@     Pw@      <@      ~@      "@     �l@      4@     @}@     @Y@     �P@     �B@     �M@     @o@      O@      w@     t@     @|@     �R@     `j@     �V@     �M@     `q@      $@     �v@      @     `b@      0@     �v@     �Q@      H@      ?@      @@      h@     �B@     Pp@     �k@     �v@      L@     �a@     �I@      B@      c@      @     �m@      @     �U@      $@     �p@      G@      =@      7@      0@      Z@      5@     �e@     �a@     `l@      D@     �Q@      8@      8@      V@      @     �b@             �H@      @     �b@      2@      .@       @      $@      M@      @      Z@     �U@     �b@      =@      0@      .@      1@     �@@       @      <@              9@       @      D@      *@      $@      @       @      <@      @     �@@      >@      F@      &@      K@      "@      @     �K@       @      ^@              8@      @     @[@      @      @      @       @      >@       @     �Q@      L@     �Z@      2@     �Q@      ;@      (@      P@             �V@      @     �B@      @      ^@      <@      ,@      .@      @      G@      ,@     @Q@      K@     @S@      &@     �A@       @      @      H@              P@              :@      @     �U@      &@      @      $@              9@      "@     �G@     �B@      I@      @     �A@      3@      @      0@              :@      @      &@      �?     �@@      1@      @      @      @      5@      @      6@      1@      ;@      @     �Q@      D@      7@     �_@      @     �^@             �N@      @     �W@      9@      3@       @      0@      V@      0@      V@     @T@     �`@      0@      9@      6@      &@     �H@      @      1@              B@      �?      >@      @      $@      @      @      =@      &@      ;@     �B@      I@      @      @      �?      �?      $@               @               @                              @              �?      �?      �?       @              ,@              4@      5@      $@     �C@      @      "@              <@      �?      >@      @      @      @      @      <@      $@      9@     �B@      B@      @      G@      2@      (@     @S@       @     �Z@              9@      @     @P@      5@      "@      @      (@     �M@      @     �N@      F@     �T@      (@      4@      @      @      C@      �?     �I@              �?      @      9@      (@      @      �?              @@      @      :@      <@     �A@      "@      :@      *@       @     �C@      �?     �K@              8@              D@      "@      @       @      (@      ;@      �?     �A@      0@      H@      @     �V@      ?@      >@     �W@      2@     �]@      @      U@      @      Z@      >@      3@      @      ;@      M@      9@     �Z@      Y@      W@      2@      O@      ,@      *@     �I@      (@     �W@      �?      M@       @     @Q@      *@      (@      �?      @      D@      @     �O@     �K@     �K@       @      M@       @      "@     �G@      &@      S@      �?      I@       @     �K@      &@      $@      �?      @      :@      @     �K@     �H@     �K@      @      =@      @      @      ;@      $@      D@      �?      0@       @      3@       @       @      �?      @      0@      �?     �B@     �@@      9@      @      =@      @       @      4@      �?      B@              A@              B@      @       @              �?      $@      @      2@      0@      >@      @      @      @      @      @      �?      2@               @              ,@       @       @               @      ,@      �?       @      @              �?       @       @      �?                       @               @              @                               @      "@              @      �?              �?       @      @      @      @      �?      0@                               @       @       @                      @      �?      @      @                      =@      1@      1@      F@      @      9@       @      :@       @     �A@      1@      @      @      4@      2@      2@      F@     �F@     �B@      $@      @      @      @      &@              @       @       @              @      @                      @       @              $@      @      @      �?       @      �?      @      &@              @       @       @              @      @                               @              @       @      @               @       @      �?                       @                                                              @                      @       @      @      �?      9@      ,@      &@     �@@      @      4@              8@       @      @@      ,@      @      @      1@      0@      2@      A@     �D@      ?@      "@      1@      *@      &@      <@      @      4@              7@      �?      :@      *@      @      @      ,@      (@      *@      A@     �D@      ;@      "@       @      �?              @       @                      �?      �?      @      �?       @              @      @      @                      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJN�mhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�;��Bw@�	           ��@       	                    @a���z�@*           �@                            �?NR]Ť@           ��@                          �:@���R��@>           �~@������������������������       ���\��@�             x@������������������������       �b����@B            �Y@                           �?���4�@�           ��@������������������������       ���;�<�@           0y@������������������������       �Vף.�@�           P�@
                             @�'�@P�@             =@������������������������       �
`��	�@
             *@������������������������       �>��_�@
             0@                           @�8��;@           ��@                            �?'I�T@W           ��@                           �?.��I�@d           p�@������������������������       ��?Ϝ�@�            @i@������������������������       �@B�؃$@�            @v@                          �:@���h@�            �x@������������������������       �
u�ǧf@�             u@������������������������       ��Ћ�m@             K@                           �?U.2��@(           @�@                           @!7�6�@�           �@������������������������       �J�N��
@^            �a@������������������������       ����t�@K           x�@                           @�^�Ē@           ��@������������������������       �� ��D@�             v@������������������������       �h|��_�@�            0q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�       �t@     @`@     @U@     pw@      >@     �}@      @     �m@      >@     @|@     �\@      I@      >@      O@     �p@     �O@     Pv@     Pr@     0|@     �R@     @b@     �R@      J@      e@      6@     ``@      @      ]@      4@     �c@     �K@      ?@      5@      C@     �\@      =@      b@     �`@     `e@     �B@     �a@     @Q@      J@     �d@      4@     ``@      @     �[@      4@     �c@     �K@      ?@      5@      C@     @\@      <@     �a@     �`@     �d@     �B@     �@@      3@      @      M@      @      D@       @      D@      $@     �H@      $@      @      $@      $@     �C@      @      =@     �C@     �P@      (@      ?@       @      @      H@      @      C@       @      <@      @     �F@      @      @      �?      @      <@      @      :@      :@     �M@      @       @      &@      �?      $@      �?       @              (@      @      @      @      �?      "@      @      &@       @      @      *@      @      @     �[@      I@     �G@      [@      *@     �V@      @     �Q@      $@     @[@     �F@      9@      &@      <@     �R@      7@     �\@     @W@      Y@      9@      E@      &@      ,@      ;@      @     �F@      �?      2@      @      >@      8@       @       @      "@      <@      "@     �F@     �B@      G@      @      Q@     �C@     �@@     @T@      $@      G@       @      J@      @     �S@      5@      7@      "@      3@      G@      ,@     @Q@      L@      K@      2@      @      @               @       @                      @              �?                                       @      �?       @              @                      @                      �?                       @              �?                                              �?      �?              @              @       @               @      �?                      @                                                       @              �?              �?             `g@      L@     �@@     �i@       @     `u@       @     �^@      $@     Pr@     �M@      3@      "@      8@     �b@      A@     �j@      d@     �q@      C@     �P@      >@      .@      W@      @     @b@              H@      �?      a@      8@      @      @      $@     �Q@      0@      Y@     �P@     @U@      ;@     �@@      .@      @     �L@      @     @U@              3@      �?      R@      0@      @       @      @      G@      $@     �P@     �E@     �O@      *@      (@       @      �?      .@              @@              (@              ;@      �?                      @      8@              7@      0@      9@      "@      5@      *@      @      E@      @     �J@              @      �?     �F@      .@      @       @      @      6@      $@     �E@      ;@      C@      @      A@      .@      $@     �A@      @     �N@              =@             @P@       @      @       @      @      8@      @      A@      7@      6@      ,@      <@      .@       @     �@@       @      G@              8@             �K@      @      @       @      @      8@      @      A@      4@      6@       @      @               @       @      �?      .@              @              $@      @                                      �?              @              @      ^@      :@      2@     �\@       @     �h@       @     �R@      "@     �c@     �A@      *@      @      ,@     �S@      2@      \@     �W@     `h@      &@     �J@      ,@      @     �P@       @     �]@       @      :@      @      T@      8@      @      @       @     �F@      @     �J@     �F@     @]@      �?      *@      @      �?      .@      �?      1@              @      �?      0@      @      �?              �?      @       @      1@       @     �A@              D@      $@      @     �I@      �?     @Y@       @      5@       @      P@      1@       @      @      �?     �D@      @      B@     �E@     �T@      �?     �P@      (@      &@     �H@             �S@             �H@      @      S@      &@      $@       @      (@      A@      *@     �M@      I@     �S@      $@     �E@      @       @      C@             �I@             �B@      �?      E@      @       @      �?      @       @      $@      ?@      >@     �A@      @      8@       @      "@      &@              ;@              (@      @      A@       @       @      �?      "@      :@      @      <@      4@     �E@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ(�KMhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @4p��@�	           ��@       	                   �7@��]�@l           �@                           �?����@T           ̔@                           �?��N%
T@B           �~@������������������������       �� ��@_            �`@������������������������       ����S��@�            `v@                            @�6B�H@           8�@������������������������       ��G���@g           ��@������������������������       ���8a��@�            `q@
                           �?���D@           ��@                            @�G)�X@�           @�@������������������������       �qQ>2,@�            �w@������������������������       �%!��8@�            �r@                          �:@̔���y@s             f@������������������������       �E�F�@D            �Y@������������������������       ��s~]@/            @R@                           �?��w��@E           ��@                           @)�K�@l           ��@                          �6@bQ_RWU@S            �`@������������������������       ��mҸ>
@C            �Z@������������������������       ����]�@             =@                            �?%�taQ@           �|@������������������������       ��Z(c��
@<            �X@������������������������       �N/颷�
@�            �v@                           @D��+?@�           ��@                           �?���ݓ�@�            �@������������������������       �M�H0��@�            @w@������������������������       �K�Z+˱@�             y@                           �?E#�
�@�            `v@������������������������       �E�L�@c            �a@������������������������       �q�[��@�             k@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@      `@     @W@     �t@     �@@     �}@      @     �k@      A@      {@      ]@     �R@     �A@     �Q@     �p@      P@     `w@     �r@     �{@     �R@     �h@     @T@     �P@     `h@      :@     �j@      @     @b@      9@      g@     �T@     �H@      ?@      L@      e@      C@     �h@     �d@     �j@      H@     �`@      @@     �@@      a@      "@      c@      �?      R@      .@     �]@     �I@      =@      @      =@     �V@      3@     �`@     @Z@     �`@      <@      L@      "@      @      E@      @      N@              ;@       @      J@      2@      @      @      @      C@       @     �I@     �G@     �L@      @      1@              @      &@       @      0@              @              *@      @       @              @      @              @      ,@      7@      @     �C@      "@      @      ?@      @      F@              5@       @     �C@      *@      @      @              ?@       @      F@     �@@      A@       @     �S@      7@      :@     �W@      @     @W@      �?     �F@      *@     �P@     �@@      6@      @      9@     �J@      1@     �T@      M@      S@      7@     �G@      &@      0@     @R@      @     �M@              6@      @     �H@      ,@      1@      @      3@      C@       @      L@      D@     �O@      0@      ?@      (@      $@      6@      �?      A@      �?      7@      @      2@      3@      @      �?      @      .@      "@      ;@      2@      *@      @      O@     �H@      A@      M@      1@     �M@      @     �R@      $@     �P@      ?@      4@      8@      ;@     @S@      3@      O@      O@     �T@      4@     �D@     �D@      A@      G@      *@      C@      @      L@      @     �K@      7@      4@      6@      ;@     �J@      0@     �L@     �J@      O@      *@      2@      8@      *@      B@       @      9@      @     �@@      �?      G@      (@      $@      &@       @      ;@      "@      ?@      :@      @@      @      7@      1@      5@      $@      @      *@              7@      @      "@      &@      $@      &@      3@      :@      @      :@      ;@      >@      @      5@       @              (@      @      5@              2@      @      &@       @               @              8@      @      @      "@      4@      @      *@      @              (@               @              1@      @      @      @              �?              ,@              @      @      "@      @       @      �?                      @      *@              �?              @      @              �?              $@      @       @      @      &@      @     �b@      H@      :@      a@      @     Pp@      �?     @S@      "@     �n@      A@      9@      @      .@     @X@      :@     @f@     �`@     @l@      :@      L@      &@      *@     �G@      @     �[@             �A@      �?     @P@      @      @              @     �B@       @     �N@     �F@     @U@      $@      @      @      @      @      �?      @@              @              .@      �?      @              @      $@      �?      0@      "@      *@      @              @      @      @              =@              �?              .@      �?      @              @      @      �?      0@      @      $@      @      @              �?      @      �?      @               @                                                      @                      @      @      �?     �I@      @      @      D@       @     �S@              @@      �?      I@      @                      @      ;@      �?     �F@      B@      R@      @       @              @      *@              1@               @      �?      .@       @                       @      $@      �?      @       @      (@             �E@      @       @      ;@       @     �N@              >@             �A@       @                       @      1@              E@      <@      N@      @      W@     �B@      *@     @V@      @     �b@      �?      E@       @     �f@      =@      6@      @       @      N@      8@     @]@     �V@     �a@      0@      O@      3@      @     @Q@      �?      ]@              <@      @     @_@      .@      1@       @      @      D@      7@     �P@     �N@      X@      ,@      ;@      "@      @     �D@      �?      O@              1@      @     �M@      @       @       @       @      3@       @      ?@      >@     �E@      @     �A@      $@      @      <@              K@              &@             �P@      $@      "@               @      5@      5@     �A@      ?@     �J@      &@      >@      2@      @      4@      @     �A@      �?      ,@      �?     �L@      ,@      @       @      @      4@      �?     �I@      =@     �F@       @      "@      @      @      $@      @      .@      �?      @              ?@      @      �?      �?              @      �?      5@       @      .@              5@      (@      @      $@              4@               @      �?      :@      "@      @      �?      @      ,@              >@      5@      >@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�\%hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �3@Gl��@�	           ��@       	                    @��ڕ��@f           8�@                          �0@�䢉�m@�           ��@                           �?)4�D�	@g            �d@������������������������       �Q���+�@9            �V@������������������������       �"s�c	@.            �R@                            �?!��@J           �@������������������������       �
˯�q�@�            �p@������������������������       ��!k�y@�           ��@
                            �?���s�K@�            pr@                          �2@��Pt�@v            �h@������������������������       �H��H�f@X            �b@������������������������       �w48#(@            �G@                          �1@)�U�B@?            @X@������������������������       �Y�?q��@%            �L@������������������������       �.���eA@             D@                          @A@��
FK�@>           v�@                            @��@&           2�@                           �?r��A@T           �@������������������������       �r�i8��@�           Є@������������������������       ���9y'�@�           |�@                          �6@�u��	@�            �@������������������������       ��
�Ae@�            �p@������������������������       �4��1x;@&            }@                           @��ݞ�	@             A@                            @c���@             5@������������������������       �u�&-�?             "@������������������������       �C8iY�o @             (@������������������������       ��s�|�@	             *@�t�bh�h5h8K ��h:��R�(KKKK��h��B         u@      `@     �Z@     �u@      C@     0{@      @     `j@     �A@     �|@     �[@      M@      F@     �S@     �m@      K@     0w@     �s@     |@     �U@     �Z@      :@      :@     �]@       @     �k@             �S@      @      k@     �@@      5@       @      &@     �S@      (@     @`@      ]@      h@      3@     �Q@      3@      1@     �V@       @      f@             @Q@      @     �f@      =@      3@       @      @     �P@       @      X@     @V@     @d@      ,@      @      @      @      @      �?      H@              .@              8@      @      �?              �?      @              1@       @      6@      �?      �?      �?       @      @              <@              @              ,@      @      �?                      �?              $@      @      1@      �?      @       @       @      �?      �?      4@              (@              $@                              �?      @              @      @      @             @P@      0@      *@      U@      @      `@              K@      @     �c@      :@      2@       @      @     �N@       @     �S@     @T@     �a@      *@      .@      @      �?      @@              6@              @      @      J@      (@      "@      �?              1@              8@      6@     �D@      @      I@      (@      (@      J@      @     �Z@             �H@             �Z@      ,@      "@      �?      @      F@       @     �K@     �M@     �X@      @      B@      @      "@      =@             �G@              "@              A@      @       @              @      (@      @      A@      ;@      ?@      @      0@      @      @      5@              ?@              @              3@      �?       @              @      @      �?      ?@      6@      8@      �?      *@      @      @      5@              .@              @              1@      �?       @              @      @              7@      2@      2@              @              �?                      0@              @               @                                       @      �?       @      @      @      �?      4@       @      @       @              0@              @              .@      @                              @      @      @      @      @      @      .@      �?      @      @              @              �?              .@      �?                              @              @       @              @      @      �?              @              $@               @                       @                               @      @              @      @             �l@     �Y@     @T@     @l@      >@     �j@      @     �`@      @@     �n@     �S@     �B@      E@     �P@     �c@      E@      n@     `i@      p@      Q@     �l@      X@     �R@      l@      >@     �j@      @     �`@      @@     `n@     �R@     �A@     �C@     �P@     �c@      E@     �m@     `i@     �o@      Q@     `d@     @P@      H@      d@      2@     `c@      @     �V@      ,@     �f@      M@      4@      8@     �C@     �[@      @@     �d@     �_@     @h@     �I@     �R@      :@      @@      N@      "@      D@       @     �H@      @     @Q@      5@      @      "@      5@      I@      3@     �G@      B@     �Q@      2@     @V@     �C@      0@     @Y@      "@     �\@       @      E@       @     @\@     �B@      *@      .@      2@     �N@      *@     @]@     �V@     �^@     �@@     �P@      ?@      ;@     �O@      (@     �L@       @     �D@      2@     �N@      1@      .@      .@      <@     �G@      $@     �R@      S@      M@      1@      ;@      *@      @      0@       @      @@              2@      @      :@      @      @      �?      @      2@      �?      ?@      ;@      9@      @     �C@      2@      6@     �G@      @      9@       @      7@      .@     �A@      *@      &@      ,@      5@      =@      "@      F@     �H@     �@@      *@       @      @      @       @                              �?               @      @       @      @                               @              @               @      @      @                                                              @               @                                              @              �?      @      �?                                                                                                                              @              �?      �?      @                                                              @               @                                                                      @               @                              �?               @               @      �?                               @                        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��dIhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �3@ �4���@�	           ��@       	                     @�&/.��@�           d�@                           @8��8�@�           D�@                           @T�͘�@X           ��@������������������������       �ݞ�v@           �y@������������������������       �Z9�2:	@K            �^@                          �1@^zj��
@>           �@������������������������       �k���8
@�            Pr@������������������������       ��(	��
@�            @k@
                           �?c��@�            �x@                           �?�V���r@j            �f@������������������������       �Kb�h�@4            �U@������������������������       �t�����	@6            @W@                          �1@��JX�|@�            �j@������������������������       �dZ�8�/@:             W@������������������������       �Q�j:޹@J             ^@                           �?=�<
�@3           `�@                           @�b��Q:@�           0�@                           �?���/@�           ؑ@������������������������       ���ρ-~@�            �t@������������������������       � �L$�7@           @�@������������������������       ��\�u�@             6@                          �4@��/M�N@>           ��@                            �?�{q`�@�            �l@������������������������       ���S��@.            @U@������������������������       �Y��d�@c            @b@                          �>@���g:@�           ��@������������������������       ��Y䫄@�           ��@������������������������       ����&y@-            @Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B         s@      a@     �U@     Pw@      B@     �@       @     @m@     �A@     �{@     �Y@      O@      I@     �S@     �m@      L@     �v@     �q@     �z@     �U@     �T@      A@      ;@      c@      "@     �j@              V@      @      h@      >@      1@      @      (@      V@       @     �b@     @W@     @i@      4@      H@      ;@      &@     �]@      @      d@             �H@      @      b@      .@      (@      @      @     �N@      @     �^@     �P@     �d@      (@      8@      $@      @     �R@      @      O@              6@      @      N@      (@      @       @      @      A@      @     �Q@      C@     �T@      $@      .@      "@      @     �I@      @      F@              0@      @      J@      $@      @       @      @      ?@      @     �H@      9@     �P@      $@      "@      �?              8@              2@              @               @       @                       @      @              5@      *@      .@              8@      1@      @     �E@      @     �X@              ;@      �?      U@      @      @      @              ;@      �?      J@      =@     �T@       @      (@      @      �?      2@      @      K@              .@              M@      @      @                      3@      �?      8@      4@      J@      �?      (@      &@      @      9@              F@              (@      �?      :@              �?      @               @              <@      "@      ?@      �?     �A@      @      0@      A@       @     �K@             �C@              H@      .@      @      �?      @      ;@      @      <@      :@     �B@       @      4@      @              0@      �?      >@              .@              8@      "@              �?      @      @      �?      ,@      $@      2@      @      *@      �?              @      �?       @              "@              @      @              �?      @      @              "@      "@      @      @      @      @              "@              6@              @              2@       @                              @      �?      @      �?      (@      @      .@      @      0@      2@      �?      9@              8@              8@      @      @               @      4@      @      ,@      0@      3@      �?      &@              "@      @      �?      &@              $@              ,@       @      @                       @              @      @      @      �?      @      @      @      &@              ,@              ,@              $@      @                       @      (@      @      $@      &@      .@             �k@     �Y@      N@     �k@      ;@     r@       @     @b@      <@     �o@     @R@     �F@      F@     �P@     �b@      H@     �j@      h@      l@     �P@      Y@      N@     �G@     �X@      5@     �W@      @     �V@      4@      Y@      ?@      4@      :@      D@      L@      =@     @Y@     �V@     �X@     �A@      Y@     �L@     �G@     �X@      .@     �W@      @     �U@      4@      Y@      >@      4@      :@      D@     �J@      <@     �X@     @V@     �X@     �A@      6@      1@      .@     �@@              A@      �?      7@      �?      ?@      *@      @      @      &@      5@      "@      9@      1@      C@      (@     �S@      D@      @@     �P@      .@     �N@      @      P@      3@     @Q@      1@      ,@      5@      =@      @@      3@     @R@      R@      N@      7@              @                      @                      @                      �?                              @      �?      @      �?                     �^@      E@      *@     �^@      @     @h@      @     �K@       @     `c@      E@      9@      2@      :@     �W@      3@     �[@     �Y@     �_@      ?@      @       @       @      7@              B@              @      @      8@      @      $@       @              (@      @      ?@      <@      9@      @      @               @      @              *@              @              @      �?      $@      @               @              *@      "@      @      �?       @       @              3@              7@                      @      1@      @              @              @      @      2@      3@      4@      @     @]@      D@      &@     �X@      @     �c@      @      I@      @     ``@     �A@      .@      $@      :@     �T@      0@      T@     �R@     @Y@      9@     �[@      C@      "@     @X@      @     @b@              I@      @     @^@      A@      .@      $@      8@     @T@      ,@     @Q@     @R@     �V@      6@      @       @       @       @              (@      @                      $@      �?                       @      �?       @      &@       @      $@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@&����@�	           ��@       	                     @���5�@c           ��@                           @"�L
�@p           ��@                            �?�Y����@�           h�@������������������������       �Oe@H            �@������������������������       �,d;�ֿ	@g            �a@                           �?-�'mw�@�             s@������������������������       �PWܜs	@N            �_@������������������������       ���o��@s            �f@
                           @1`h[_|@�            @x@                           @�P�T~:@�             u@������������������������       ���W�(�@�            �p@������������������������       �Š�2G�@0            �Q@                           �?J>�=��@"             J@������������������������       �z�>�@             8@������������������������       �:*/);q@             <@                           �?�8�J(k@?           ̣@                          �9@�d.#@�           ��@                           @��oT�@�           `�@������������������������       ��n��۬@	           �z@������������������������       �ۓq[�@�            �s@                           @`�S��@           |@������������������������       �}�ϭ"�@�             n@������������������������       �/��3�@�             j@                           �?��ڕ�L@C           �@                           @G���@�           p�@������������������������       ��ȉ-�y@w            `i@������������������������       �|�xT�2@           0|@                           @�q��.�@�           X�@������������������������       �
F�gn�@9           0@������������������������       ��H�2�@u             g@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@      `@      X@     @u@     �E@     �|@      @     �j@      ;@     �}@     @[@      T@      =@      Q@     `m@     �O@     �x@     �q@     �z@     �T@     �X@      :@      ;@      `@      "@      i@      �?     @Q@      @     �i@      ?@      4@      @      $@     �Q@      0@     `b@      W@     `i@      4@     �P@      2@      3@     @X@      @      d@             �F@      @      c@      $@      0@      @       @      H@      $@     @W@     �N@     `d@      ,@      F@      (@      *@     �O@      @     �Z@              A@      @      _@      @      &@      @       @     �D@      @     �L@      C@      [@      *@      B@      "@      *@     �J@      @     �R@              <@      @     �X@      @      "@       @             �B@      @     �C@      ?@      V@      (@       @      @              $@      �?      @@              @              :@               @      �?       @      @              2@      @      4@      �?      6@      @      @      A@             �J@              &@              =@      @      @              @      @      @      B@      7@     �K@      �?      @      �?       @      0@              @@              @              &@      �?      @                      @              (@      $@      6@      �?      0@      @      @      2@              5@               @              2@      @                      @      @      @      8@      *@     �@@              @@       @       @      ?@      @     �D@      �?      8@             �I@      5@      @               @      7@      @      K@      ?@      D@      @      =@       @      @      8@      @      A@      �?      2@              B@      5@      @                      7@      @      K@      <@      B@      @      7@      @      @      1@      @      8@      �?      .@              8@      1@      @                      4@       @     �G@      6@     �A@       @      @      @      @      @              $@              @              (@      @                              @      @      @      @      �?       @      @               @      @              @              @              .@              �?               @                              @      @       @       @               @      @              @               @              �?                                                                       @       @      �?                      �?                              @              ,@              �?               @                              @       @             �o@     �Y@     @Q@     �j@      A@      p@      @      b@      8@     �p@     �S@      N@      :@      M@     �d@     �G@      o@      h@     `l@     �O@      \@     �L@     �E@     @Y@      8@     @W@      @     �V@      0@     �[@     �D@     �A@      *@     �C@      P@      :@      [@      U@      Y@      B@     �S@      ;@      9@     �K@      4@     @R@       @     �J@      ,@     �T@      <@      "@      @      9@      A@      ,@     �R@      C@      O@      ;@      C@      "@      &@      =@      @     �J@       @     �A@      @     �E@      7@      @      @      3@      4@      &@     �D@      3@     �@@      9@      D@      2@      ,@      :@      ,@      4@              2@      @      D@      @      @      @      @      ,@      @     �@@      3@      =@       @      A@      >@      2@      G@      @      4@      �?      C@       @      <@      *@      :@      @      ,@      >@      (@      A@      G@      C@      "@      ,@      8@      (@      9@               @      �?      8@       @      $@      &@      .@              @      .@      @      :@      8@      3@              4@      @      @      5@      @      (@              ,@              2@       @      &@      @      $@      .@      @       @      6@      3@      "@     �a@      G@      :@     �[@      $@     �d@              K@       @     �c@     �B@      9@      *@      3@      Y@      5@     �a@     @[@     �_@      ;@      V@      6@      $@      I@      @     �U@              8@      @      S@      5@      "@      @      @      I@      0@      G@     �P@     �I@      0@     �@@       @              .@      @      5@              ,@              :@      @      �?      @              6@       @      @      4@      3@      @     �K@      4@      $@     �A@      @     @P@              $@      @      I@      ,@       @      @      @      <@       @      D@     �G@      @@      *@     �J@      8@      0@     �N@      @     �S@              >@      @     @T@      0@      0@      @      .@      I@      @     �W@      E@      S@      &@     �C@      2@      @     �G@      @     �P@              =@      �?      N@      *@      &@      @      @     �C@      @      Q@      ?@     �F@       @      ,@      @      $@      ,@              *@              �?      @      5@      @      @              &@      &@              ;@      &@      ?@      @�t�bub��     hhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�x�^hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�U�Wޥ@�	           ��@       	                     @Cu��n@�           h�@                            �?�����@M           ��@                           �?@ΨY@L           (�@������������������������       �K{��@*           �|@������������������������       �&�6�]�@"           ��@                           �?�*H�
@           �y@������������������������       �4���,�	@g            �d@������������������������       ��i|$m
@�            `n@
                           �?�map�@�           ��@                           �?3�L
?~@�            �v@������������������������       �C��M@a            �c@������������������������       ��H��}@x            �i@                           �?y��"ȧ@�            Pr@������������������������       ���q�
@c             c@������������������������       ��k�ao�
@Z            �a@                            @X��&u�@�           T�@                           �?x���_1@�           Ԑ@                           @'M3O�@)           p~@������������������������       ��ӢB@           `{@������������������������       ���hE�@            �H@                          �?@�1���@q           p�@������������������������       �7�X�@R           ��@������������������������       �A�@             L@                           @��Dq�R@A            ~@                           �?��=�,@�            �t@������������������������       �ņ=��@J            @[@������������������������       ���%� @�            �k@                           @��i��%@`            �b@������������������������       �7����@S             `@������������������������       ��	�o��@             4@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     @\@      V@     �v@      C@     �~@       @     `n@      B@     @|@      Z@     �M@      A@     �O@     @m@      M@     �v@      t@     �z@     �Y@     `e@      G@     �I@      l@      3@      v@             �a@      7@     0s@      G@     �@@      *@      3@     �\@      8@     @n@     �g@     r@     �H@     @[@     �A@      ?@     �g@      @      p@             �V@      2@     �n@      7@      ?@      (@      @      U@      ,@     @d@     @`@     `k@     �A@     @U@     �@@      <@     �b@      @     @e@             @P@      $@     �f@      6@      7@      (@      @      Q@      ,@      ]@     �Y@     �e@      =@     �B@      &@      @     �K@      @     @Q@             �@@      @     �Q@      @      @               @      =@      �?     �@@      =@      P@      @      H@      6@      9@     @W@      �?     @Y@              @@      @     �[@      3@      3@      (@      @     �C@      *@     �T@     @R@      [@      6@      8@       @      @      E@      �?      V@              9@       @      O@      �?       @               @      0@              G@      <@     �G@      @      @      �?      @      (@             �B@              @              7@              @              �?      @              :@      5@      4@      @      5@      �?              >@      �?     �I@              2@       @     �C@      �?      @              �?      (@              4@      @      ;@      �?      O@      &@      4@      A@      (@      X@             �I@      @     �O@      7@       @      �?      (@      ?@      $@      T@      N@     �Q@      ,@      C@      @      1@      *@      &@      F@              =@      @      8@      4@       @      �?      &@      0@      @      J@     �A@      =@       @      =@      @      $@      @      �?      9@              @               @      (@              �?       @      $@      �?      2@      .@      (@      @      "@      @      @      $@      $@      3@              8@      @      0@       @       @              "@      @       @      A@      4@      1@      @      8@      @      @      5@      �?      J@              6@             �C@      @                      �?      .@      @      <@      9@     �D@      @      &@      �?       @      .@      �?      ;@              .@              ,@                                      $@      �?      @      *@      >@      @      *@      @      �?      @              9@              @              9@      @                      �?      @      @      5@      (@      &@             �a@     �P@     �B@      a@      3@     @a@       @     �Y@      *@      b@      M@      :@      5@      F@     �]@      A@      _@     @`@     `a@      K@     �[@      E@      0@     �Y@      &@     @\@      @      P@      @      Z@     �@@      .@      *@      5@     �V@      ;@      V@      T@     @Y@      B@     �J@      (@      &@      H@      @     �M@      @      ?@      @      I@      .@       @      @      @     �K@      $@     �C@      ;@      ;@      6@     �D@      &@      $@      H@      @      M@      @      =@      @      F@      .@       @      @      @     �C@      $@     �@@      9@      :@      6@      (@      �?      �?              �?      �?               @              @                                      0@              @       @      �?             �L@      >@      @     �K@      @      K@      @     �@@              K@      2@      *@      @      .@     �A@      1@     �H@     �J@     �R@      ,@     �K@      4@      @      I@      @     �E@      @     �@@             �J@      2@      $@      @      .@     �A@      .@      E@     �H@      P@      ,@       @      $@              @              &@                              �?              @      �?                       @      @      @      $@              @@      9@      5@      A@       @      9@       @      C@      "@     �D@      9@      &@       @      7@      =@      @      B@      I@      C@      2@      0@      ,@      2@      <@      @      1@       @      =@      @      6@      4@      $@       @      .@      0@      @      <@      D@      6@      2@      @      @      @      &@      �?      @              &@      @      (@      @      @              @      @       @      $@      "@      @      @      "@      $@      (@      1@      @      ,@       @      2@      @      $@      *@      @       @      (@      (@       @      2@      ?@      .@      *@      0@      &@      @      @      @       @              "@       @      3@      @      �?      @       @      *@      @       @      $@      0@              0@      &@      @      @      @       @              "@       @      &@      @      �?      @       @      (@      �?      @       @      ,@                                       @                                               @       @                              �?       @      �?       @       @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJDbyhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @�i�S@�	           ��@                            @;�i.@�           ��@                           @�K�^Q�@x           l�@                            �?�gm~k�@i           �@������������������������       ��~��@�           ��@������������������������       �g�7,�	@{             i@������������������������       ��X�1R�@             6@                           �?��{y�@           ��@	       
                   �?@U�aqv}@�           p�@������������������������       ��@/�ZH@�           Ѓ@������������������������       ��/�Ѩ�	@             J@                           @�M���
@Y            �`@������������������������       �rt��4@$             L@������������������������       ����2i@5            �S@                          �4@�Tw�_�@           �@                          �2@��bi@9           `�@                           @�I^0�
@q           �@������������������������       ��(,$
@�            �s@������������������������       ������
@�            `r@                            �?���Ր@�            �r@������������������������       �bw@Ș@n             d@������������������������       ��H-z
@Z            @a@                          �8@8�@lT�@�           h�@                           �?���/�@            |@������������������������       �=̔�.�@�            `k@������������������������       ��5��@�            �l@                            �?b�J��@�            �r@������������������������       ���Y�A�
@2             T@������������������������       �>?3(�@�            `k@�t�bh�h5h8K ��h:��R�(KKKK��h��B        Pv@     �a@     �W@      v@     �D@      �@      @     �k@      ;@     �}@     @W@      L@      A@     �L@     �j@     �L@     �w@     �r@     �z@     �Q@     �h@     @X@     �Q@      k@      A@      o@      @     �b@      8@     `m@     @P@      ?@      8@     �A@      `@      C@     `i@      h@     @j@     �I@     �^@      M@      @@     @c@      3@     �b@      @     @V@      *@     �d@     �@@      2@      (@      1@     �V@      8@     @^@     �_@     �b@      C@     �^@     �J@      @@     @c@      .@     �b@      @      U@      *@     �d@     �@@      2@      &@      1@     @V@      8@     �]@     �_@     `b@      C@     �Y@      H@      >@      a@      &@     �_@      @     �R@      *@     ``@     �@@      0@      &@      *@     @R@      8@     @X@      [@      `@     �A@      4@      @       @      2@      @      7@              "@             �A@               @              @      0@              6@      2@      3@      @              @                      @                      @              �?                      �?              �?               @      �?       @             @S@     �C@      C@     �O@      .@     �X@              O@      &@      Q@      @@      *@      (@      2@     �C@      ,@     �T@     @P@     �N@      *@     �P@      :@      A@     �I@      .@     �S@              H@      $@     �K@      :@      $@      "@      2@      C@      @     @R@      L@      K@      &@      O@      1@      >@     �F@      .@     @S@             �G@      $@     �H@      5@      $@      @      0@      C@      @     @R@      G@      K@      &@      @      "@      @      @               @              �?              @      @              @       @                              $@                      &@      *@      @      (@              4@              ,@      �?      *@      @      @      @              �?      @      "@      "@      @       @      @              �?      @               @               @              @      @      @                              �?       @      @      �?       @      @      *@      @      @              (@              @      �?      @                      @              �?      @      @      @      @             �c@     �E@      9@      a@      @     �p@              R@      @     �m@      <@      9@      $@      6@     @U@      3@      f@     �Z@     `k@      3@     @Q@      0@      "@     �P@      �?     @c@             �I@             �a@      &@      ,@      @             �B@      &@     @Y@     �M@     `b@      (@     �H@      (@      "@      A@      �?     �X@             �A@             �]@       @       @      @              5@      $@     �Q@      B@     �X@      @      >@      @      �?      8@      �?      M@              (@              I@      �?      @                      &@      @     �A@      .@      M@      �?      3@      @       @      $@              D@              7@              Q@      �?       @      @              $@      @     �A@      5@     �D@      @      4@      @             �@@              L@              0@              9@      "@      @      @              0@      �?      ?@      7@      H@       @      *@      @              ,@              ?@              $@              3@      @      �?      @              (@              *@      1@      1@      @      @      �?              3@              9@              @              @      @      @                      @      �?      2@      @      ?@      @     @V@      ;@      0@     �Q@      @     �[@              5@      @     �W@      1@      &@      @      6@      H@       @      S@      H@      R@      @      L@      8@      "@     �D@             @R@              0@       @      J@      @      @              (@      @@      @     �K@      9@      @@      @      5@       @      �?      9@              F@              @       @      =@      @                      @      6@      @      :@      &@      &@      @     �A@      0@       @      0@              =@              (@              7@      @      @              @      $@       @      =@      ,@      5@             �@@      @      @      =@      @     �B@              @      �?      E@      $@      @      @      $@      0@      @      5@      7@      D@      @      @               @      @              5@               @              @       @                      @      @      �?       @      @      (@       @      <@      @      @      8@      @      0@              @      �?     �B@       @      @      @      @      &@       @      *@      2@      <@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ2��-hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@^��Y�@�	           ��@       	                    @�v9Ps@0           f�@                          �3@5"yk��@p           H�@                           �?k��ii@]           Ȍ@������������������������       ��RE��@�            0s@������������������������       ��؊q�
@�           0�@                           �?��d��@           �{@������������������������       ��-%@�            �p@������������������������       � �%�Ԋ@k            �e@
                           @S��yR@�           �@                            @ܐ���+@�           (�@������������������������       ��a̡@.           `@������������������������       ��C.@            �i@                           @f�a�1@             <@������������������������       ���.�@             1@������������������������       �lofON@             &@                          �:@�K�&x�@�           X�@                            @!Τ�A@           ��@                           @���@           �@������������������������       ���"�
�@p           h�@������������������������       �O ����@�            �n@                           �?>0����@�            �x@������������������������       �8$�(*@a             b@������������������������       ��kA��@�            `o@                           �?��I��@�           8�@                          �?@���5�@v             g@������������������������       ����^$�@[            �a@������������������������       �5�:W�9@            �E@                           �?�{)e�@           �z@������������������������       ���'G9�@_            @b@������������������������       ��RWˍ@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       `t@     �`@      U@     �u@      A@      �@      @     @m@      @@      z@     @Z@     �M@      ?@     �O@     �m@     �U@     �u@     �s@     �{@     �V@     �c@      M@      ?@      j@      @     �t@      �?     @]@      &@      m@     �B@      D@      &@      .@     @Z@      E@     �h@     �f@     �p@      H@     �Y@      =@      2@      c@      @     �l@      �?      S@      @     �e@      4@      $@      @      &@     �L@      0@     @_@     �\@     �e@      A@     �N@      6@      ,@     �W@      @     �b@      �?     �I@      @     �`@      2@       @      @      @     �D@      @     �T@     @Q@      a@      2@      2@      @       @      ?@       @      ?@      �?      5@      @      9@      (@      @              @      4@      @      0@      ?@     �M@      "@     �E@      .@      @      P@      �?     @]@              >@      �?     �[@      @       @      @      �?      5@      @     �P@      C@     @S@      "@     �D@      @      @     �L@      �?     �T@              9@      @      C@       @       @      @      @      0@      "@     �E@      G@     �C@      0@      9@      @      @      A@      �?      H@              2@              0@      �?       @              @       @      �?      ;@      <@      ?@      (@      0@      �?              7@              A@              @      @      6@      �?              @               @       @      0@      2@       @      @      K@      =@      *@      L@      @      Y@             �D@      @      N@      1@      >@      @      @      H@      :@     @R@     �P@     �W@      ,@      H@      <@      *@     �K@      @      Y@              A@      @      M@      1@      >@      �?      @      H@      :@     �Q@      P@      W@      ,@      5@      6@      @      E@             �Q@              7@      @      E@      $@      0@      �?      @      D@      3@      J@      F@      S@      $@      ;@      @      @      *@      @      >@              &@      �?      0@      @      ,@                       @      @      2@      4@      0@      @      @      �?              �?                              @               @                      @                              @      @       @              @      �?                                              @              �?                      @                              @                              @                      �?                              �?              �?                                                              @       @             @e@     @S@     �J@     �a@      ;@     @g@      @     @]@      5@     �f@      Q@      3@      4@      H@     �`@      F@      c@     ``@      f@      E@     �\@      K@      @@     �W@      .@     �a@       @     @R@      .@     @b@      G@      @      @      @@     �U@      :@     �Y@     �Q@      Z@      ?@     �T@     �A@      5@     �P@      $@     �Z@       @      B@      @     @Y@      <@       @              (@     �M@      2@     @R@      C@      V@      4@      M@      1@      2@     �G@       @     @T@       @      8@      �?      S@      ,@      �?               @     �A@      &@      J@      9@     �M@      4@      9@      2@      @      3@       @      9@              (@      @      9@      ,@      �?              @      8@      @      5@      *@      =@              ?@      3@      &@      =@      @      B@             �B@      $@     �F@      2@      @      @      4@      <@       @      >@     �@@      0@      &@      (@      @      $@      $@       @      @              &@      @      4@      @      �?              @      @      @      $@      .@      (@      �?      3@      *@      �?      3@      @      =@              :@      @      9@      (@      @      @      0@      5@      @      4@      2@      @      $@      L@      7@      5@     �F@      (@      F@      @      F@      @     �B@      6@      *@      .@      0@     �G@      2@     �H@      N@     @R@      &@      @      @       @      0@      @      *@              ,@              @      @      @      "@      @      4@      �?      *@      @@      (@      @      @       @       @      &@      �?      $@              (@              @      @      @      "@      �?      .@              (@      8@      (@      @      �?      @      @      @      @      @               @                      �?                      @      @      �?      �?       @                     �H@      1@      *@      =@       @      ?@      @      >@      @      ?@      0@      @      @      (@      ;@      1@      B@      <@     �N@      @      <@      @       @      @      @       @       @       @      @      $@       @       @      @      @      "@      @      1@      @      (@      @      5@      ,@      &@      9@       @      7@      �?      6@              5@       @      @       @       @      2@      (@      3@      7@     �H@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJF.�dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�#> ^z@�	           ��@       	                    �?��[�ػ@           \�@                           �?���r�x@[           �@                          �:@�@M3�@�            @j@������������������������       ��~
M@v            �f@������������������������       �����H�@             >@                           �?��@�             u@������������������������       �|im'�@G             ^@������������������������       ����|�@�             k@
                           @�투�@�           Ԑ@                            @�z��@j           p�@������������������������       ��D��0�@I           H�@������������������������       �7og�@!           P|@                           @I�-A{@@            �Y@������������������������       �`ޗZ�[@3            �S@������������������������       ���H+-@             8@                            @�+2:r*@�           �@                          �4@�yg%��@z           ܜ@                           �?kv���o@W           x�@������������������������       ��s��<)
@(           �}@������������������������       �P���j @/           @                           �?\��G�@#           @�@������������������������       ��Ĵ��@           z@������������������������       �ɂ��&�@           p|@                           @G��+8@           �{@                           @*l�� @�            @j@������������������������       �B-XL}�@Z            ``@������������������������       ��_6�2@-            �S@                          �5@#���@�             m@������������������������       ��
�͏n@`            @c@������������������������       �~����d@7            �S@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        t@      a@     �V@     �v@     �C@     �|@      @     �m@      6@     P}@     �\@     �K@      >@     @P@      n@      M@     `w@      r@      }@      S@     �_@     �Q@      M@     @a@      >@     @]@      @     �[@      .@     `c@     �J@     �A@      ,@      E@     �X@      A@     @b@     �`@      i@      D@     �G@      4@      5@     �F@      �?     �I@      @      A@      @     �H@      0@      @       @      (@      <@      (@     �G@     �B@     @X@      *@      .@      @      *@      *@      �?      9@      @      .@      �?      6@      @      @              @      (@      @      @      .@      E@      @      .@       @      &@      *@      �?      9@              $@              .@      @      @              @      &@      @      @      .@      B@      @              �?       @                              @      @      �?      @      �?                      �?      �?      �?      �?              @              @@      1@       @      @@              :@              3@      @      ;@      &@       @       @      @      0@       @      D@      6@     �K@      @      2@      @      @      ,@              &@              @      @      @       @       @              @       @      �?      (@      @      1@       @      ,@      ,@      @      2@              .@              *@              7@      @               @       @      ,@      @      <@      0@      C@      @     �S@     �I@     �B@     @W@      =@     �P@       @      S@      "@     �Z@     �B@      >@      (@      >@     �Q@      6@     �X@     �X@     �Y@      ;@     @Q@      E@      B@     �T@      9@      O@       @     �P@      "@     �V@     �A@      >@      (@      =@      L@      5@     �U@     @W@     @Y@      9@      <@      9@      (@      L@      "@      =@       @      =@      @     �L@      .@      1@       @      $@      B@      ,@      I@      E@     �P@      (@     �D@      1@      8@      ;@      0@     �@@             �B@      @      A@      4@      *@      @      3@      4@      @     �B@     �I@     �A@      *@      $@      "@      �?      $@      @      @              $@              .@       @                      �?      .@      �?      (@      @       @       @      @      @      �?       @       @      @              @              .@       @                      �?      &@      �?      "@      @      �?       @      @      @               @       @                      @                                                      @              @      �?      �?             �h@     �P@      @@      l@      "@     Pu@      �?     �_@      @     �s@      O@      4@      0@      7@     �a@      8@     �l@     `c@     �p@      B@     �c@      H@      8@     �f@      @     �q@      �?     �V@      @     �o@      F@      *@      *@      5@      ]@      .@      h@      `@     �l@      7@      I@      9@      $@      V@             �e@             �G@       @      c@      1@      $@      @      @     �K@      @     @Y@      Q@      c@      "@      7@      *@      �?     �F@             �W@              6@              R@      @      @      @              7@             �C@      C@     �V@      @      ;@      (@      "@     �E@              T@              9@       @      T@      *@      @      �?      @      @@      @      O@      >@     �O@      @     @[@      7@      ,@      W@      @     @\@      �?     �E@      @      Y@      ;@      @      @      1@     �N@      &@      W@     �N@     �R@      ,@      L@      (@      @      L@      @     �L@      �?      3@      @      E@      2@              @      @      ?@      @     �@@      ;@      9@      &@     �J@      &@      &@      B@              L@              8@              M@      "@      @      @      $@      >@      @     �M@      A@      I@      @     �B@      2@       @     �F@      @      K@             �B@      �?      O@      2@      @      @       @      :@      "@     �A@      :@      C@      *@      *@      &@       @      .@      @      =@              5@              9@      0@      @               @      *@       @      (@      $@      6@      $@      (@      @      �?      &@      @      5@              (@              0@      "@      @                      @       @      "@      @      @      @      �?      @      �?      @               @              "@              "@      @                       @      @              @      @      .@      @      8@      @      @      >@              9@              0@      �?     �B@       @      @      @              *@      @      7@      0@      0@      @      *@      @       @      (@              0@              *@              ;@      �?      @                      &@      @      1@      &@      ,@      �?      &@              @      2@              "@              @      �?      $@      �?              @               @       @      @      @       @       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJv�9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@����s@�	           ��@       	                     @}�����@�           �@                           �?Ec6�*)@d           ��@                           �?��l�t@G            @������������������������       �x�����@q            �e@������������������������       �8A��l'@�            Pt@                           @S�� eC@           4�@������������������������       �`���0�@>           �@������������������������       �h%��x@�           x�@
                          �4@�HWJܗ@�           ��@                           @�U��@)           �|@������������������������       ���[��@�            �u@������������������������       ��I�K0�@I            �[@                           �?��G,��@i            �d@������������������������       ��X��T@,             Q@������������������������       �^C��Z@=             X@                           �?�){W@�           `�@                           �?~�zTx@           �z@                            �?�$��@v             g@������������������������       �\e9)W
@$            �K@������������������������       �7�p��9@R            @`@                            @����@�            �n@������������������������       �O4,T�~@f            �d@������������������������       ����.��@0            �T@                           @��Y!0a@�           ��@                           �?Xֿۙ@�           �@������������������������       ��Az��)@�            �t@������������������������       ���W��@�            �s@                           @�E�hP@           pz@������������������������       �USs�d�@�            Pt@������������������������       �k)���(	@=            �X@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �`@     @V@     �t@     �E@     �~@      @     `k@      5@     �|@     �X@      M@     �A@     �R@      p@      P@     �w@     �r@     `}@     �M@     @d@      R@      I@     �k@      5@     Pv@      @     ``@       @      s@     �J@      B@      "@      @@     �b@      A@     �n@     �g@     pr@      D@     �\@      K@      ?@      e@      "@     �q@      �?     �U@      @     �l@      =@      7@      "@      9@     �[@      5@     �g@     �`@     �m@      ?@     �E@      2@      4@      J@      @     �L@      �?      8@      @      H@      @       @       @      @      >@      $@     �@@      E@     @R@      .@      7@       @      @      0@      @      6@              "@      �?      0@                              �?      &@              (@      "@      A@      @      4@      $@      .@      B@      @     �A@      �?      .@      @      @@      @       @       @      @      3@      $@      5@     �@@     �C@      (@      R@      B@      &@      ]@      @     @l@             �O@             �f@      9@      .@      @      3@     @T@      &@     `c@     �V@     �d@      0@      4@       @      @      J@      �?     @Q@              4@             �S@      *@      @      �?      .@     �A@      $@      R@      D@     �J@      &@      J@      <@      @      P@       @     �c@             �E@             �Y@      (@       @      @      @      G@      �?     �T@      I@     @\@      @     �G@      2@      3@      K@      (@     �R@       @      F@       @     @S@      8@      *@              @      D@      *@     �L@      M@      L@      "@     �C@      &@      ,@      G@      (@      L@       @      6@       @      G@      3@      $@              @      @@      (@      D@      D@     �H@      @      8@      @      "@      D@      $@     �G@       @      0@      �?      @@      *@      @               @      <@       @      =@      <@     �G@       @      .@      @      @      @       @      "@              @      �?      ,@      @      @              �?      @      @      &@      (@       @      @       @      @      @       @              2@              6@              ?@      @      @              @       @      �?      1@      2@      @       @      @      �?      @      @              @              "@              "@      �?      �?               @       @      �?      @      *@      @      �?      �?      @       @      @              *@              *@              6@      @       @               @      @              (@      @       @      �?     `c@     �O@     �C@     �[@      6@     �`@      @      V@      *@     @c@     �F@      6@      :@     �E@     @Z@      >@      a@      \@     �e@      3@     �A@       @      .@      D@       @     �G@              =@       @      F@      .@      @       @       @     �@@      @     �G@     �A@      F@      &@      2@       @       @      0@       @      5@              1@              8@      @       @       @              $@       @      "@      4@      1@       @      @      �?       @      "@       @      @              @              @                                      @                      �?      $@      @      *@      �?      @      @              .@              $@              3@      @       @       @              @       @      "@      3@      @      @      1@      @      @      8@              :@              (@       @      4@       @      @      @       @      7@      @      C@      .@      ;@      @      (@      @      @      $@              7@              @              0@      @      @      @       @      1@      @      9@      "@      2@       @      @      @      �?      ,@              @               @       @      @      @      �?                      @       @      *@      @      "@      �?      ^@     �K@      8@     �Q@      4@      V@      @     �M@      &@     �[@      >@      .@      2@     �D@      R@      7@     @V@     @S@     ``@       @     @R@      C@      (@      G@      (@      P@      @      B@      "@     �J@      ;@      &@       @      9@     �A@      "@      I@     �I@      R@      @     �@@      5@      &@      4@      @      3@      @      =@      @      1@      (@      $@      @      0@      2@      @      8@     �@@     �A@      @      D@      1@      �?      :@      @     �F@              @      @      B@      .@      �?      @      "@      1@      @      :@      2@     �B@       @     �G@      1@      (@      8@       @      8@              7@       @     �L@      @      @      $@      0@     �B@      ,@     �C@      :@     �M@      �?      ?@      0@      (@      4@      @      2@              6@       @      E@      @      @      $@      .@      8@      &@      A@      ,@     �C@      �?      0@      �?              @      �?      @              �?              .@                              �?      *@      @      @      (@      4@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�K�QhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @a�1A��@�	           ��@       	                   �3@��vN�:@�           F�@                           @[F�S@�           ��@                           @����@           @y@������������������������       ��	���@�            `s@������������������������       ��P<@;            �W@                            �?f-��u�
@�           ��@������������������������       ��m�@#           �|@������������������������       ���Դ�	@}            �h@
                           @b�M�^@Z           �@                           @�P��@�           ��@������������������������       �XΒH��@�           �@������������������������       �o�}6t@Z           (�@                           �?���#մ@\            �a@������������������������       ���b{%�@             8@������������������������       �L�|���@L            �]@                          �5@�ߘ��@�           ��@                          �1@qE�Tz@K           �@                          �0@-(&�2�@_            `b@������������������������       ��+���@             D@������������������������       ��*9kk�@F            �Z@                           @\4�r��@�            �v@������������������������       �ށB��@@�            �p@������������������������       ��+�q��@;            @W@                           @brŵ4@`           H�@                           �?u���=@A           �@������������������������       ��,��	@U            �`@������������������������       ���kO@�            Pw@                          �7@�B�X
@            �F@������������������������       ���@             0@������������������������       ��|�Ԏ@             =@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        s@     �a@      X@     �t@     �B@     @@       @     @m@      3@     P{@      `@     �P@      C@     �Q@     �k@     �M@     �u@     �s@     p|@     @Y@     �j@      X@     �O@     p@      6@     �y@      @     @d@      $@     �t@     �U@     �D@      9@      E@     @d@      C@     �o@     `k@     �u@     �P@     �F@      6@      &@     �[@       @     �f@             �O@      �?      a@      =@      .@      @      @     �O@       @     �W@      R@     @f@      3@      2@      @       @     �M@       @      C@              3@      �?      D@      3@      @              @      ;@      @      B@      A@     @Q@      *@      ,@      @      @      D@       @      =@              ,@      �?     �B@      ,@      @              @      :@      �?      ;@      9@      J@      *@      @              @      3@              "@              @              @      @      �?              @      �?      @      "@      "@      1@              ;@      0@      @     �I@              b@              F@             @X@      $@      &@      @      �?      B@      @      M@      C@     @[@      @      6@      .@       @     �C@              V@             �@@             @S@      "@      @      @              7@      @      E@      <@     �Q@      @      @      �?      �?      (@             �L@              &@              4@      �?      @       @      �?      *@              0@      $@     �C@      �?     �d@     �R@      J@     `b@      4@      l@      @     �X@      "@     �h@     �L@      :@      4@     �A@     �X@      >@      d@     `b@      e@      H@     `b@      P@     �I@     �a@      2@     �j@      @      W@      "@      g@     �J@      5@      4@     �A@     �V@      9@     �a@     @_@     �c@      H@     �W@     �H@      B@      U@      (@      d@      @     �Q@      @     �`@     �B@      ,@      0@      *@     �M@      ,@     @V@     �S@     �X@      <@     �J@      .@      .@      M@      @      K@      �?      6@      @      J@      0@      @      @      6@      @@      &@     �J@     �G@     �L@      4@      4@      $@      �?      @       @      $@              @              *@      @      @                       @      @      2@      6@      *@               @       @      �?      �?              @                              �?                                               @      @      @                      2@       @              @       @      @              @              (@      @      @                       @      @      *@      0@      *@             �W@      F@     �@@     �R@      .@      W@       @      R@      "@     �Y@     �E@      :@      *@      <@      N@      5@      X@     �W@      [@      A@      M@      0@      &@      C@       @     �N@      �?      =@       @     �L@       @      .@      @      @      7@      &@     �H@      G@     �K@      (@      ,@      @      @      (@      @      7@      �?       @              9@       @      @               @      @      @      .@      @      @       @       @       @               @               @      �?      @              &@      �?                               @              @              �?       @      (@      �?      @      $@      @      .@              @              ,@      �?      @               @      @      @      &@      @      @      @      F@      *@       @      :@      @      C@              5@       @      @@      @       @      @      @      1@      @      A@      D@     �I@      @      B@      "@      �?      5@      @      =@              (@       @      6@      @      �?      @      @      .@      @      9@      :@     �F@      @       @      @      @      @      �?      "@              "@              $@              @              �?       @      �?      "@      ,@      @              B@      <@      6@      B@      @      ?@      �?     �E@      @      G@     �A@      &@      $@      6@     �B@      $@     �G@     �H@     �J@      6@      A@      9@      6@     �@@      @      >@      �?     �E@      @     �C@      =@      &@      "@      6@      =@      $@      G@      G@     �G@      2@       @      @      @      @       @      @              .@              3@      @      @              @      &@      @      (@       @       @      &@      :@      6@      1@      :@      @      9@      �?      <@      @      4@      8@      @      "@      0@      2@      @      A@      C@     �C@      @       @      @              @              �?                              @      @              �?               @              �?      @      @      @                              @              �?                              @                                      @                      @      �?               @      @                                                               @      @              �?              @              �?              @      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�G�}hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@Ҥ@���@�	           ��@       	                     @g��8p�@�           Ƣ@                            �?T�L�+@d           ̛@                           @��w�e@p           ��@������������������������       ��NjQ�|@�           �@������������������������       ��9��@@�            @v@                          �0@�ԏ��@�            �x@������������������������       �;I�� @             E@������������������������       �Ws���@�            v@
                           �?s5\��@�           ��@                          �1@
��	 �@�            �q@������������������������       �E���@+            �O@������������������������       �*���@�             k@                           �?���PY�@�            �u@������������������������       ��~�{��	@             J@������������������������       ���~�w�@�            @r@                           @���z�@�           ��@                           �?�q�4�@           $�@                           �?��]~�B@�           �@������������������������       �td�ƈ�@�            �l@������������������������       ���]L�I@d           ȁ@                           �?~���z@           �z@������������������������       �� Z�M@|            �g@������������������������       ���3�u@�            �m@                           @d�Dk*@�            �q@                            �?C���<�
@R            �`@������������������������       ���Y0@             A@������������������������       ������	@>            �X@                           �?}m#&@e             c@������������������������       �&���
@+             Q@������������������������       ��W�. t@:             U@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     ``@     �U@     �v@     �H@      ~@      (@     `l@      >@     �{@     �X@      P@      ?@     �L@     @o@     @R@     �v@     �s@      z@     @T@      h@     @R@      F@     `k@      4@     �u@      @     @`@      *@     �r@     �J@      C@      ,@      5@      b@      C@     `m@      h@      r@      C@     �`@      I@      9@     �f@      @     Pp@              X@      $@     @l@      @@      >@      "@      &@      \@      7@     �e@     �`@     �m@      ?@     @Z@      G@      8@     �b@      @      f@             �R@      @     �f@      ;@      7@      @      @     �U@      7@     �`@     �[@     �f@      8@     �P@     �@@      3@     �_@       @     �_@             �I@      @      `@      0@      7@      @      @     @P@      5@     �Z@      S@     @`@      5@     �C@      *@      @      6@       @     �H@              7@      @     �I@      &@              �?              5@       @      :@     �A@      I@      @      ;@      @      �?      A@      @     @U@              6@      @      G@      @      @       @      @      :@              D@      7@      L@      @                               @              (@                              $@              �?              �?      $@               @              @              ;@      @      �?      @@      @     @R@              6@      @      B@      @      @       @      @      0@              C@      7@      J@      @      N@      7@      3@     �B@      *@     �T@      @      A@      @     �R@      5@       @      @      $@     �@@      .@     �O@      M@      K@      @      B@       @      @      ;@      @      B@              &@              A@      ,@       @      @       @      (@       @      8@      =@      7@      @      @       @      �?       @      �?      @               @              $@      @                               @       @      @      @              �?      =@              @      3@      @      =@              "@              8@      "@       @      @       @      $@              3@      9@      7@      @      8@      .@      (@      $@       @     �G@      @      7@      @     �D@      @      @       @       @      5@      *@     �C@      =@      ?@       @      @      @      �?      �?              @                       @      (@                                      �?      @      �?       @      @      �?      1@      (@      &@      "@       @     �D@      @      7@      �?      =@      @      @       @       @      4@      $@      C@      5@      9@      �?     �a@      M@      E@     �b@      =@     @a@      "@     @X@      1@     �a@     �F@      :@      1@      B@     @Z@     �A@      `@     �_@     �_@     �E@     �X@      I@     �B@      `@      ;@     @\@      @     @W@      1@     �Y@     �@@      8@      .@      <@     @T@      A@      W@     �Y@     �Y@     �C@      P@     �A@      A@     @U@      6@      J@      @      K@      @      O@      6@      6@      ,@      7@      J@      5@     �N@     @Q@     �Q@      5@      4@      *@      @      =@      @      6@      @      $@      �?      9@      @      "@       @      @      9@              1@      &@      3@      @      F@      6@      ?@      L@      3@      >@       @      F@      @     �B@      0@      *@      (@      3@      ;@      5@      F@      M@     �I@      1@     �A@      .@      @     �E@      @     �N@             �C@      $@     �D@      &@       @      �?      @      =@      *@      ?@     �@@     �@@      2@      3@      @      �?      4@       @      5@              0@      $@      2@      @       @              �?      ,@      @      .@      2@      @      ,@      0@      &@       @      7@      @      D@              7@              7@       @              �?      @      .@      @      0@      .@      :@      @      F@       @      @      4@       @      9@       @      @              C@      (@       @       @       @      8@      �?      B@      9@      7@      @      ,@       @      @      "@              ,@              @              9@      @      �?                       @              8@       @      (@      �?      @               @      @              @              @               @                                      �?                              @              $@       @      @       @               @                              1@      @      �?                      @              8@       @      "@      �?      >@      @              &@       @      &@       @      �?              *@      @      �?       @       @      0@      �?      (@      1@      &@      @      0@       @              @       @      @       @                      @      @      �?                      @      �?       @      (@      @              ,@      @               @               @              �?               @       @               @       @      "@              @      @       @      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJe9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?7%=��@�	           ��@       	                     �?*���t@A           h�@                          �8@` k���@�           ��@                           �?͸f.�@l           ��@������������������������       �B�`�|@v            �f@������������������������       ��`��V
@�            �x@                           �?�֫�Ȕ@^            �b@������������������������       ��n�7��@)            �M@������������������������       �&s��!@5             W@
                          �3@����@w            �@                           �?ݞ.�B@�            `m@������������������������       ����M�q
@             B@������������������������       �+��C�	@�            �h@                            @��]8"�@�            �u@������������������������       ��q(M�@W             a@������������������������       �0�Lο@�             j@                            @tۉ��(@v           ^�@                            �?9���O�@�           �@                           �?�K�Ym�@�           ��@������������������������       ��K$э�@u           ؂@������������������������       �?�n�`�@           h�@                           �?��;2q@           �y@������������������������       ��=V�^�
@f             c@������������������������       ���L!�U@�             p@                          �6@���g��@�           `�@                           �?��܋�@@            �x@������������������������       ���މ+@w            �f@������������������������       ���%(��@�             k@                           @��Ɇ�^@�             v@������������������������       �j2ј�'@�             k@������������������������       �/R��Z�@_             a@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       t@     @b@     @X@     �v@      C@     �|@      @     �n@      D@     �{@     @Z@     @Q@     �@@     �N@      l@      L@     �v@     �s@     |@      R@      [@      @@      A@      ]@      "@     �g@             �X@      @      d@      8@      3@      @      (@      U@      "@     @^@     �W@     �c@      <@     �M@      7@      3@     �R@      @      [@             �F@      @      [@      &@      @      @      @      D@      �?     �Q@     �E@     �W@       @     �I@      .@      @     @Q@      @     @X@             �C@      @      U@      @      @               @      8@              K@      ?@     �S@      @      0@      @       @      :@       @      6@              .@      �?      0@      @      @               @      (@              2@      @      <@             �A@      "@      @     �E@      @     �R@              8@       @      Q@      �?                              (@              B@      9@      I@      @       @       @      ,@      @      �?      &@              @              8@      @              @       @      0@      �?      0@      (@      0@      @      �?       @      @      @      �?      @               @              $@      �?               @              @              @      @      @      @      @      @      $@                      @              @              ,@      @              �?       @      "@      �?      *@      @      $@             �H@      "@      .@      E@       @     �T@              K@      @      J@      *@      *@               @      F@       @     �I@     �I@      O@      4@      4@       @      @      .@             �J@              1@              .@      @      �?               @      1@       @      0@      7@      D@      @      @       @      @       @              @               @               @                                      @      �?      @              @              0@                      *@              H@              .@              *@      @      �?               @      *@      �?      (@      7@      A@      @      =@      @      &@      ;@       @      >@             �B@      @     �B@      $@      (@              @      ;@      @     �A@      <@      6@      .@      &@              @       @              (@              "@              3@      @      @              @      (@       @      ,@      .@      @      $@      2@      @      @      3@       @      2@              <@      @      2@      @      @              �?      .@      @      5@      *@      0@      @     �j@     �\@     �O@     `o@      =@     �p@      @     �b@     �@@     �q@     @T@      I@      >@     �H@     �a@     �G@      n@     �k@     Pr@      F@      c@     �S@     �C@     �g@      3@     �g@      @      Y@      7@      k@      F@      B@      1@      :@     �[@      A@      e@     �b@     �m@      :@     @_@     �N@      @@     �a@      ,@      _@      @     �S@      0@     @c@      D@      <@      0@      6@      S@      =@     �a@      `@      h@      8@     �F@      ;@      6@     �O@       @      F@      @      F@      ,@      F@      (@      .@      @      (@      ?@      3@      J@      E@     �V@      &@      T@      A@      $@     �S@      @      T@              A@       @     �[@      <@      *@      &@      $@     �F@      $@     �V@     �U@     �Y@      *@      <@      1@      @      H@      @     �P@              6@      @     �O@      @       @      �?      @      A@      @      :@      3@     �F@       @      @      @              ,@      �?      C@              @      @      9@      �?       @              �?      &@       @      @      &@      2@      �?      8@      $@      @      A@      @      <@              .@      �?      C@      @      @      �?      @      7@      @      6@       @      ;@      �?      N@      B@      8@     �N@      $@     @T@      @      H@      $@     �P@     �B@      ,@      *@      7@      >@      *@     �Q@      R@      L@      2@      ?@      0@      $@      A@      @     �M@       @      7@             �H@      5@      $@       @      @      1@      @     �E@      B@      7@      @      7@      @       @      2@       @      <@              "@              4@      &@       @               @      $@      @      (@      (@      3@      @       @      *@       @      0@       @      ?@       @      ,@              =@      $@       @       @       @      @      �?      ?@      8@      @      @      =@      4@      ,@      ;@      @      6@       @      9@      $@      2@      0@      @      &@      3@      *@       @      <@      B@     �@@      &@      *@      "@       @      2@      @      .@       @      ,@       @      @      &@              @      *@      &@      @      7@      9@      1@      "@      0@      &@      @      "@       @      @              &@       @      *@      @      @      @      @       @      @      @      &@      0@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�ndhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @v���ª@�	           ��@       	                   �4@b��@�           ҥ@                            �?����@R           ,�@                          �3@U���@�           L�@������������������������       ���ǔ��@           ��@������������������������       ��f�~ �@�            `l@                           @A��2@�            �s@������������������������       ���X1�w@b            �c@������������������������       �'j��&C@b            @c@
                           �?�4���@�           x�@                            �?��N��@�           ��@������������������������       ��i+�Y�@�            `s@������������������������       ��ej�b@�            �q@                           @"���@           h�@������������������������       �^l�a�@�           ��@������������������������       �Ea}2�b@0            @T@                           �?�61��@�           ��@                          �:@�0*�V@�           �@                          �3@�7^Ŋ�@Y            �@������������������������       �	����@�            `j@������������������������       �)���s @�            u@                          �?@rsP|@c            �c@������������������������       �?��y�(@A            @Z@������������������������       ���z�WN@"            �J@                           @��ɲrc@           �y@                           �?�eg_z�@_            �c@������������������������       �&T��@.            �S@������������������������       �P���%@1            @S@                          �1@d!�Z�@�             p@������������������������       ��pjh��@            �D@������������������������       �<W�'r@�             k@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     ``@     �V@      u@      E@     �~@      @     `n@     �B@     @|@      X@     �L@      B@      M@     �o@     @Q@     @w@     �s@     z@     @T@      o@      U@      F@     @n@      5@     �v@      @     @c@      4@     �u@     �L@     �G@      9@      A@     �h@     �E@     0p@     �k@     @t@      J@      T@      ;@      0@     �a@      @     �j@             �R@      @      g@      8@      1@      @       @     �W@      3@      ]@      \@      g@      ;@      P@      7@      $@     �[@       @     �b@              H@      @     �b@      7@      *@      @      @     @R@      3@     @V@     �W@      a@      5@     �E@      4@      "@     �V@       @     @^@              A@      @     �^@      5@      (@      @      @      J@      (@     @R@     �N@      ^@      &@      5@      @      �?      4@              >@              ,@       @      :@       @      �?      @              5@      @      0@     �@@      0@      $@      0@      @      @      ?@      �?     �O@              :@             �A@      �?      @              @      6@              ;@      2@     �H@      @      (@      @              4@      �?      6@              6@              6@      �?      �?              @      @              &@      ,@      0@      @      @              @      &@             �D@              @              *@              @                      1@              0@      @     �@@       @      e@     �L@      <@     @Y@      2@     �b@      @      T@      ,@     �d@     �@@      >@      2@      :@     �Y@      8@     �a@     �[@     `a@      9@     �J@      <@      3@     �E@      *@      E@      @     �I@      "@     �P@      (@      2@      @      "@      D@      .@     �M@     �F@      J@      "@      <@      1@       @      6@      &@      0@      @     �A@      "@      A@      @      @      @      @      1@      @      0@      7@      B@      @      9@      &@      &@      5@       @      :@              0@              @@      @      (@      @       @      7@      "@     �E@      6@      0@      @      ]@      =@      "@      M@      @      [@      �?      =@      @      Y@      5@      (@      &@      1@     �O@      "@      U@     @P@     �U@      0@     �Z@      7@      "@     �L@      @     �Y@      �?      4@      @     @W@      2@      (@      @      1@     �K@      "@     @S@     �L@     �R@      0@      "@      @              �?              @              "@              @      @              @               @              @       @      *@              T@     �G@     �G@     �W@      5@     @`@       @     @V@      1@     �Y@     �C@      $@      &@      8@      L@      :@     @\@     �V@     @W@      =@     �E@     �@@     �E@      L@      2@     �R@       @     �G@      1@      H@      7@      @      &@      6@      ?@      0@     @S@     @Q@     �J@      1@      C@      1@      <@      B@      0@     �Q@              B@      ,@      C@      2@      @       @      1@      7@      $@     �Q@      J@      B@      ,@      &@      @      $@      *@      @      D@              $@              ,@      $@      �?              @      *@      @      9@      5@      4@      @      ;@      (@      2@      7@      $@      ?@              :@      ,@      8@       @      @       @      *@      $@      @      G@      ?@      0@      &@      @      0@      .@      4@       @      @       @      &@      @      $@      @      �?      @      @       @      @      @      1@      1@      @      @      @      $@      1@      �?               @      "@      @      @              �?               @       @      @      @       @      0@                      "@      @      @      �?      @               @              @      @              @      @                       @      "@      �?      @     �B@      ,@      @      C@      @      L@              E@              K@      0@      @               @      9@      $@      B@      5@      D@      (@      .@      $@      @      $@      �?      9@              :@              *@       @      �?                       @      @      $@       @      &@      @      "@      @       @      @              @              3@              @      @      �?                      @              @      �?      @      @      @      @       @      @      �?      3@              @              @      @                              @      @      @      �?      @      �?      6@      @              <@       @      ?@              0@             �D@       @      @               @      1@      @      :@      3@      =@      @      @                      �?      �?      ,@              �?              $@              �?              �?      �?               @               @       @      1@      @              ;@      �?      1@              .@              ?@       @       @              �?      0@      @      8@      3@      ;@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ(hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�W�>��@�	           ��@       	                    �?�o64.�@�           $�@                           @G�TDB@�           Ї@                           �?�ޒ�@           �{@������������������������       �E�Q&@           �y@������������������������       �����@             <@                            �?.�̝��
@�            t@������������������������       ����K�		@q            @g@������������������������       �t�̹<@S            �`@
                          �1@y�'�@�           x�@                          �0@,n-��o@T            `b@������������������������       ���/#z@             L@������������������������       �/�Qt~�
@6            �V@                           �?�P��@@�           ��@������������������������       �Ʋ��.@H           h�@������������������������       ���;lex@G            �[@                          �6@d�	0�@�           ��@                            �?�y���(@z           �@                           @���u @           Pz@������������������������       ��Tt���@�            @k@������������������������       �;��|�	@�            `i@                           @ɇH�;@j           ��@������������������������       ����u~`@�           ��@������������������������       ��n.��@�             v@                           @�7���l@_            �@                            �? ���@�           H�@������������������������       ���(���@           �{@������������������������       ��]0�@�            �t@                           �?-:�@n            `g@������������������������       ��5�~� 
@'            �R@������������������������       ���}��@G            @\@�t�b�?     h�h5h8K ��h:��R�(KKKK��h��B`       �t@     �a@     �S@     �t@     �I@     �}@       @     @h@      =@     �|@     @W@     �J@      G@      M@     �p@     �R@     �w@     @r@     p}@     �S@     �Y@      G@      :@     �_@      3@     `m@      �?     �T@      "@      i@      C@      &@      "@      3@     @Y@      5@      a@     �^@     �h@      E@      J@      3@      @     �O@      (@     �]@      �?     �D@       @     @\@      7@      @      @      @      G@      @      J@     �N@      [@      ;@      <@      .@      @      C@      @     �K@      �?      <@       @     �P@      1@      @      @      @      ?@      @      @@     �A@      I@      .@      :@      .@      @      :@      @     �H@      �?      <@       @     @P@      .@      @      @      @      ?@      @      ?@     �@@     �H@      .@       @                      (@              @                              �?       @                      �?                      �?       @      �?              8@      @              9@      @     �O@              *@             �G@      @      �?                      .@       @      4@      :@      M@      (@      1@      @              .@      �?     �D@              @             �A@      @      �?                      @              &@      ,@      ?@              @                      $@      @      6@              @              (@      @                              "@       @      "@      (@      ;@      (@      I@      ;@      5@     �O@      @     @]@              E@      @     �U@      .@      @      @      *@     �K@      0@      U@     �N@     �V@      .@       @              @      *@      �?     �B@               @      @      ,@              �?              @      (@      @      $@      1@      ,@       @      �?                       @              2@              @               @                              �?      @      @      "@       @      @              �?              @      &@      �?      3@              @      @      (@              �?               @      @              �?      .@       @       @      H@      ;@      1@      I@      @      T@              A@      @     @R@      .@      @      @      $@     �E@      $@     �R@      F@     @S@      *@     �E@      5@      (@     �G@      @     �J@              ?@      @      O@      .@      @      @      @     �B@      "@     �Q@      >@     �O@      &@      @      @      @      @       @      ;@              @      �?      &@              �?       @      @      @      �?      @      ,@      ,@       @     �l@     �W@     �J@     �i@      @@      n@      �?     �[@      4@     pp@     �K@      E@     �B@     �C@      e@      K@     @n@     @e@      q@     �B@     �\@     �E@     �A@      ^@      0@     �f@             �O@      @     �d@      A@      ;@      5@      (@      W@      8@      d@     @[@      d@      1@      2@      4@      ,@     �D@              N@              *@      @     �J@      @      @      &@      @      3@      �?      J@      8@     �P@      @      *@       @       @      :@              ;@              "@      @      (@      @      @      "@      @      ,@      �?      2@      0@      D@      @      @      2@      @      .@             �@@              @             �D@      @       @       @              @              A@       @      ;@              X@      7@      5@     �S@      0@     �^@              I@      @     @\@      ;@      4@      $@       @     @R@      7@     @[@     @U@     @W@      $@     @Q@      .@      1@     �K@      ,@     �P@              ;@      @     @U@      :@      $@      @      @      I@      4@      M@      L@     �F@      @      ;@       @      @      8@       @      L@              7@      �?      <@      �?      $@      @       @      7@      @     �I@      =@      H@      @     �\@      J@      2@     �U@      0@     �L@      �?      H@      *@     @X@      5@      .@      0@      ;@     @S@      >@     @T@     �N@      \@      4@     @Y@     �E@      (@     �T@      "@     �E@      �?      D@      (@     �R@      2@      *@      $@      4@      K@      4@     �L@     �J@      X@      2@      O@      ;@      @      G@      @      8@              4@       @     �B@      *@      (@      @      1@     �@@      1@     �@@      6@      L@      "@     �C@      0@       @     �B@      @      3@      �?      4@      $@     �B@      @      �?      @      @      5@      @      8@      ?@      D@      "@      ,@      "@      @      @      @      ,@               @      �?      7@      @       @      @      @      7@      $@      8@       @      0@       @      "@              @      �?      @      @                      �?      0@       @                              ,@      @      @      �?      @              @      "@      �?      @       @      $@               @              @      �?       @      @      @      "@      @      1@      @      $@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ���BhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�e���@�	           ��@       	                     @�8�E�x@?           z�@                           @$^&�z@�           �@                          �4@�x����@,           �@������������������������       �4��ӡa@�           �@������������������������       �h7$I,@h             d@                          �3@��N�Y�@�           �@������������������������       ��ף~F�
@9           P~@������������������������       ����K_@w            �g@
                           @���=��@c           ��@                          �3@:osn�@5           �~@������������������������       ��U)1@�             u@������������������������       �6���R@b            �b@                          �3@,`�W}�@.            �S@������������������������       ���E�@            �G@������������������������       ��8�R�@             @@                          @A@=r�kB�@x           0�@                          �?@
Va��@c           ��@                           �?��ګ!b@(           �@������������������������       ��|����@           ��@������������������������       ���p7�@           x�@                            �?�n���;@;            �X@������������������������       �ޟ��ij@             ;@������������������������       �D��S Q@*             R@                           @�7��r}@             C@������������������������       �P:&У@             8@������������������������       �����G@	             ,@�t�bh�h5h8K ��h:��R�(KKKK��h��B�       �s@     `c@      T@     u@      D@     �~@      @     @m@      3@     �}@     @`@      O@     �B@      S@     �o@     �N@     `v@     �r@     �y@      T@     `b@      R@     �A@     �g@      "@     �r@             @_@      @     p@      K@      A@      0@      2@     �^@      6@     @k@      e@     �q@      C@      U@     �I@      8@     �a@       @     @l@             �S@      @     �h@      >@      =@      *@      ,@     �V@      2@     �d@     �^@     �k@      <@     �F@      =@      .@     �V@       @     �W@             �F@       @     @[@      0@      7@      @      *@      L@      1@     �X@     �P@     �^@      3@     �C@      1@      .@     �R@       @     @R@              D@              V@      .@      0@      �?       @      I@      ,@     �R@      J@     �[@      2@      @      (@              1@              5@              @       @      5@      �?      @      @      @      @      @      7@      .@      (@      �?     �C@      6@      "@     �I@             �`@             �@@       @     @V@      ,@      @      "@      �?     �A@      �?     �P@     �K@     @Y@      "@      9@      2@      @     �F@             �W@              =@      �?     �Q@      @      @       @              :@      �?     �G@      @@     @S@      @      ,@      @      @      @              C@              @      �?      2@      $@      �?      @      �?      "@              4@      7@      8@      @     �O@      5@      &@     �H@      @     �Q@             �G@       @     �M@      8@      @      @      @      ?@      @     �J@      G@      M@      $@     �L@      2@      $@     �B@      @     �O@             �C@       @     �J@      8@      @      @      �?      3@      @     �H@      C@     �I@       @      D@      (@      $@      =@       @      H@              9@              >@      4@      �?      �?      �?      0@      @     �A@      7@     �B@      @      1@      @               @      @      .@              ,@       @      7@      @      @       @              @              ,@      .@      ,@      @      @      @      �?      (@              @               @              @                              @      (@              @       @      @       @      @       @      �?      @              @               @              @                              @       @                      @      @       @              �?              @              �?                              �?                                      $@              @      @      @             @e@     �T@     �F@     @b@      ?@      h@      @     @[@      *@     �j@      S@      <@      5@      M@     ``@     �C@     �a@      `@     �`@      E@     @e@     @R@      E@     �a@      ?@      h@      @     �Y@      *@     �j@      R@      ;@      1@     �L@      `@     �C@     �a@     �_@     �`@      E@     @d@     �M@      D@      a@      :@      f@       @      Y@      *@      j@      R@      ;@      ,@     �J@     �_@      B@     @`@     �]@     �_@      D@     �N@      9@      3@     �P@      *@     �Q@       @      N@      @     @Y@     �B@      5@      @     �D@     �N@      6@     @P@      N@      P@      4@     @Y@      A@      5@     �Q@      *@     �Z@              D@      @      [@     �A@      @      "@      (@     �P@      ,@     @P@      M@      O@      4@       @      ,@       @      @      @      .@       @      @              @                      @      @       @      @      $@      "@      @       @              @                              $@              @              �?                      �?      �?       @      �?              �?      @               @      $@       @      @      @      @       @                      @                       @      @               @      $@       @      @       @              $@      @      @                              @                      @      �?      @      �?       @                      �?      �?                      @      @      �?                              @                      @              @      �?       @                              �?                      @              @                               @                      �?      �?                                              �?                �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJMS/hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����@�	           ��@       	                   �2@�~z&
�@�           Ԗ@                           �?��򍽇@           �|@                           �?G�	��\@           �z@������������������������       �������
@�             o@������������������������       �y�� @t            �f@                           �? 	R�H@            �@@������������������������       �rD��*@             ,@������������������������       ���y�=� @             3@
                           �?�^�1b@x           0�@                           �?K.H��@           �y@������������������������       ��eH��@V            @a@������������������������       �E���U!@�            Pq@                          �<@��>�@q           8�@������������������������       ���~���@U           ��@������������������������       �"!&:?T@             J@                           @U9��I@           (�@                          @A@�S+:@v           �@                          �?@;l
���@a           `�@������������������������       ���X��@@           l�@������������������������       ����YU�@!            �N@                           @`�����@             A@������������������������       ����=�@             1@������������������������       �Ii��G@
             1@                            �?�a;��@�           h�@                           @r����w@�             r@������������������������       ��X]"{�@V             b@������������������������       �_�E�P@\             b@                           @'Al��@�           ��@������������������������       ��@Z�k*@w            `h@������������������������       ��&���@g           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@      ^@     �V@     �r@      H@     �@       @     �m@     �A@     P{@     �\@     �Q@      G@     �K@      o@      Q@     �w@     `s@     �z@     @V@     @Z@      =@     �C@      [@      *@     �l@             �\@      �?     �d@     �A@      8@      @      4@     �V@      3@     �_@     @_@     `e@      B@      <@      @       @      B@      @     @V@              @@              P@              �?       @      @      8@      @     �D@     �A@      R@      &@      <@      @       @      >@      @     �T@              >@             �L@              �?      �?      @      8@      @     �D@      ;@      R@      &@      ,@      @      @      ,@       @     �B@              7@              C@                      �?      �?      $@              ;@      (@      J@      "@      ,@      �?      @      0@       @      G@              @              3@              �?              @      ,@      @      ,@      .@      4@       @              �?              @              @               @              @                      �?       @                               @                              �?              �?               @               @                                               @                              @                                              @              @                              @                      �?                                       @                     @S@      7@      ?@      R@      "@     �a@             �T@      �?     �Y@     �A@      7@      @      *@     �P@      0@     @U@     �V@     �X@      9@      5@      (@      8@      @@      @      G@              G@      �?     �B@      .@      *@      @       @      9@      *@      =@      E@      =@      $@      &@      @      @      "@      @      5@               @              "@      $@      @      �?              *@      @      @      .@      "@      @      $@      @      2@      7@      @      9@              C@      �?      <@      @       @      @       @      (@      "@      8@      ;@      4@      @      L@      &@      @      D@       @     �W@             �B@             �P@      4@      $@              @      E@      @      L@      H@     �Q@      .@     �J@      "@      @      D@       @     �T@             �B@             �L@      4@      $@              @      C@             �K@     �C@     @P@      *@      @       @      �?                      *@                              "@                                      @      @      �?      "@      @       @     `j@     �V@      J@      h@     �A@     pq@       @     �^@      A@     �p@     �S@     �G@     �C@     �A@     �c@     �H@      p@      g@      p@     �J@     �\@     �M@      C@     �\@      <@     ``@      @     �T@      :@     �[@      K@     �@@      :@      8@     �X@      >@     ``@     �[@     �b@      A@     @\@     �K@     �A@      [@      <@     ``@      @     �T@      :@     �[@     �H@      ?@      2@      8@     �X@      >@     ``@     @[@     �b@      A@     @[@      J@      ?@      [@      <@      _@      @     @T@      :@     �Z@     �H@      ?@      0@      5@     �X@      ;@      _@     �Y@     �a@      :@      @      @      @                      @              �?              @                       @      @              @      @      @      "@       @      �?      @      @      @                              �?              �?      @       @       @              �?                       @                      �?      @      @                                                              @              @              �?                                                      �?              @                              �?              �?      �?       @      @                                       @                     @X@      @@      ,@     �S@      @     �b@      �?     �C@       @     �c@      9@      ,@      *@      &@     �M@      3@     @_@     �R@     �Z@      3@      7@      ,@       @      @@              B@              (@              I@       @              @       @      1@      @     �A@      ,@      =@       @      "@      @      @      8@              2@              @              ;@       @              @      �?      @       @       @      @      4@       @      ,@      @      @       @              2@              @              7@      @                      �?      ,@      �?      ;@       @      "@             �R@      2@      @     �G@      @      \@      �?      ;@       @     @[@      1@      ,@       @      "@      E@      0@     �V@      N@     �S@      1@      2@      @              1@      @      4@              @              H@      @      @                      @      "@      <@      $@      0@       @      L@      *@      @      >@      @      W@      �?      5@       @     �N@      (@      &@       @      "@     �B@      @      O@      I@      O@      .@�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�hhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���*.�@�	           ��@       	                   �:@T�|M�	@           D�@                           �?>s��@2           �@                            �?��\[S@*           �|@������������������������       �-ۙ��@d             d@������������������������       �!Z~uW�@�            �r@                           @����@           ��@������������������������       �<U��1�@�           �@������������������������       ��ߣR�x@             ;@
                           �?�|�s<@�            �t@                            @h>9eX�@7            �T@������������������������       ���ONH,@%            �M@������������������������       �7�u`\
@             7@                           @��Z���@�             o@������������������������       �k�,�@@            �Y@������������������������       �?��g�d@^            @b@                          �6@{�[t}@�           �@                          �4@�T�5��@�           �@                           �?Nmaf@�           ,�@������������������������       ��[N4�@x           ��@������������������������       �>5 BW�@�           h�@                          �5@��p��@�            �v@������������������������       ��0��?p@�            @j@������������������������       ���rT@d            �c@                           @Ui�2�@�           ��@                           @�~g+Y�@?           0~@������������������������       �z{�q4�@           y@������������������������       �`Y�H�@3            �T@                           �?���6�@�            `k@������������������������       �9�N�@:            @T@������������������������       ���]���@W            @a@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �`@     �V@     �v@     �I@     �}@      @     Pp@      A@     �{@      \@      K@      B@     �S@      n@      K@     Pv@     0r@     z@     �V@      a@      O@     �O@      b@      ?@      _@      @     ``@      9@     �c@     �K@      A@      :@      L@      V@      5@      a@     @`@     @c@     �B@     �\@      B@      I@     �[@      >@      \@       @     @W@      7@     �`@     �F@      :@      *@     �E@      S@      .@     �_@      X@     @[@      A@     �D@      &@      :@      H@       @      I@      �?      4@      @      E@      2@      @       @      $@      =@      @      D@     �@@     �I@      *@       @              "@      2@              1@      �?      (@              .@      @      �?       @      @       @      @      "@      0@      7@       @     �@@      &@      1@      >@       @     �@@               @      @      ;@      ,@      @              @      5@      @      ?@      1@      <@      @     @R@      9@      8@     �O@      <@      O@      �?     @R@      0@     �V@      ;@      3@      &@     �@@     �G@       @     �U@     �O@      M@      5@     �Q@      7@      8@     �O@      4@      O@      �?     �Q@      0@     �V@      ;@      3@      &@     �@@      F@       @     @S@     �O@      M@      5@      @       @                       @                       @                                                      @              "@                              6@      :@      *@     �@@      �?      (@      @      C@       @      9@      $@       @      *@      *@      (@      @      &@      A@     �F@      @       @      @      @       @              "@      @      "@              &@       @      @      @      @      @              @      @      *@                      @      �?       @               @              @              "@      �?      @      @       @      @              @       @       @               @      @       @                      �?      @       @               @      �?                      �?                              �?      @              4@      3@      $@      ?@      �?      @      �?      =@       @      ,@       @      @      $@      $@       @      @       @      ?@      @@      @      �?       @      @      5@              �?      �?      *@      �?      @      @       @               @       @      @      @      1@      *@      �?      3@      &@      @      $@      �?       @              0@      �?      &@      @      �?      $@       @      @       @      @      ,@      3@       @     �f@      R@      <@     �k@      4@     v@      �?     @`@      "@      r@     �L@      4@      $@      6@      c@     �@@     �k@      d@     pp@      K@     @V@     �D@      4@     `d@      "@      q@              Z@      @     �i@     �A@      2@      @      "@     @W@      5@     `c@     �[@     �i@     �A@     �Q@      ;@      $@     @_@       @     �j@             �T@      @      e@      >@      @      @      @     �Q@      1@     @Z@      V@     `e@      7@     �C@      0@      @     �L@      @     �Y@              D@             �T@      @      �?      @             �@@       @      I@      G@      Y@      1@      ?@      &@      @      Q@       @     �[@             �E@      @     �U@      9@      @      �?      @     �B@      .@     �K@      E@     �Q@      @      3@      ,@      $@      C@      �?      N@              5@       @      B@      @      &@      �?      @      7@      @      I@      6@     �@@      (@      (@      &@       @      1@              <@              &@              .@       @      $@      �?      @      *@       @     �A@      2@      5@      @      @      @       @      5@      �?      @@              $@       @      5@      @      �?                      $@       @      .@      @      (@      @     �V@      ?@       @      N@      &@     @T@      �?      :@      @      U@      6@       @      @      *@     �M@      (@     @P@     �I@     �M@      3@     �K@      6@      @     �E@      "@     �R@      �?      .@       @     �O@      ,@      �?      @      "@      B@      @     �C@      <@      E@      0@      G@      5@      @     �A@      @     �J@              *@      �?     �L@      &@      �?      �?      @     �A@      @      A@      :@      @@      ,@      "@      �?      �?       @       @      5@      �?       @      �?      @      @               @      @      �?      �?      @       @      $@       @      B@      "@      @      1@       @      @              &@       @      5@       @      �?              @      7@      @      :@      7@      1@      @      ,@      �?              "@       @      @              @       @       @      �?      �?                      @       @      "@      &@      @      @      6@       @      @       @              @               @              *@      @                      @      0@      @      1@      (@      (@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJB�UhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?g.���@�	           ��@       	                     @g4M�K�@           ��@                           @:����"@d           ��@                          �8@WLe�@�           p�@������������������������       �D�z�B�@?           ؀@������������������������       ��=ʞ�#@�            `j@                          �8@���χ@�            pp@������������������������       �/��Ә�@\             c@������������������������       ��Ns�Hj@B            �[@
                           �?	��6@�           ��@                          �9@�����@m             g@������������������������       ��1�vz�@Y            �b@������������������������       ���\�
�
@             A@                          �:@9�z��9@@           �@������������������������       ��vL�2@�            �x@������������������������       �}�\j�2@J             \@                           @ʖ"M�@�           F�@                          �4@�1G�l@           ��@                          �2@S�0�^�@�           Ȑ@������������������������       ��ۤ���@�           ��@������������������������       ��l_!�@�            �w@                           �?Q�lIQ�@c           ��@������������������������       �P�P��@�            �u@������������������������       ��5�h�@~           ��@                            �?��I���@t            �g@                           �?�%SFH@>            @X@������������������������       �E�4��@            �B@������������������������       ��s��b
@'             N@                          �7@ppJAF(@6            �W@������������������������       ��O�:@&             Q@������������������������       ���v��@             :@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       @t@     `a@     �T@     `x@     �E@     �}@       @     �i@      @@     �|@     �\@     �T@     �F@      O@     �m@     �O@     �u@     @q@     0|@      S@     `a@     �R@      M@      f@      ;@     �a@       @     �Z@      6@      d@     �J@      G@      7@      B@     @X@      A@     �a@     �`@     �f@      D@     @S@      J@      4@     �^@      .@      T@      @      K@      &@      ^@      4@      9@      &@      1@      K@      9@     �V@     @R@     �]@      7@      K@      <@      ,@     @X@      @      R@      @      D@      @     �V@      2@      4@       @       @      F@      .@      N@     �O@     �U@      2@     �C@      (@       @      R@      @      M@              8@      @     �Q@      &@      &@       @       @      =@      "@      F@     �C@     @S@      2@      .@      0@      @      9@      @      ,@      @      0@      �?      4@      @      "@      @              .@      @      0@      8@      "@              7@      8@      @      :@      "@       @              ,@      @      >@       @      @      @      "@      $@      $@      ?@      $@     �@@      @      1@      6@      @      @      @      �?              "@      @      ,@       @      @              @      "@      �?      4@      @      4@       @      @       @       @      3@      @      @              @              0@               @      @      @      �?      "@      &@      @      *@      @      O@      7@      C@      K@      (@      O@      @      J@      &@     �D@     �@@      5@      (@      3@     �E@      "@     �H@      O@      P@      1@      4@      @      0@      ,@       @      2@      @      @              (@      @      @               @      *@       @      *@      2@      4@       @      0@      @      0@      ,@       @      &@              @              $@      @      @              �?      "@       @      (@      0@      1@              @       @                              @      @                       @      �?                      �?      @              �?       @      @       @      E@      1@      6@      D@      $@      F@             �F@      &@      =@      :@      ,@      (@      1@      >@      @      B@      F@      F@      .@      @@      &@      ,@      6@       @      F@             �@@      $@      7@      :@      &@      "@      *@      7@      @     �@@      ?@      >@      .@      $@      @       @      2@       @                      (@      �?      @              @      @      @      @       @      @      *@      ,@              g@      P@      9@     �j@      0@     �t@              Y@      $@     pr@     �N@     �B@      6@      :@     �a@      =@      j@     �a@     �p@      B@     �e@     �J@      8@      j@      ,@     �r@              V@      $@     �q@      K@     �@@      2@      :@      _@      5@      g@      `@     `n@      B@     @R@      0@      "@     @\@      �?     @f@             �H@       @     �d@      2@      1@       @      @      N@      $@     �W@      S@     `d@      0@     �C@       @      @     �S@      �?     �Z@             �C@             @^@      &@      *@      @      @     �C@      @     �L@      D@     �Z@      @      A@       @      @      A@             �Q@              $@       @     �E@      @      @       @              5@      @      C@      B@      L@      $@     �X@     �B@      .@     �W@      *@      ^@             �C@       @      ^@      B@      0@      $@      4@      P@      &@     �V@     �J@      T@      4@     �C@      @      (@     �@@      @      H@              7@             �C@       @      @       @      @      <@      �?      A@      4@     �A@      @      N@      >@      @      O@       @      R@              0@       @     @T@      <@      (@       @      .@      B@      $@      L@     �@@     �F@      *@      *@      &@      �?      @       @      B@              (@              &@      @      @      @              0@       @      8@      (@      9@              "@      @               @              (@              $@               @      @              @              *@               @      @      .@              @                                       @              @               @                                      &@              �?      @      �?               @      @               @              @              @              @      @              @               @              @       @      ,@              @      @      �?      @       @      8@               @              @      @      @                      @       @      0@      @      $@              @                      @       @      7@                              �?      �?      @                       @      @      "@      @      @                      @      �?                      �?               @               @      @                              �?      �?      @              @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��3hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @.���@�	           ��@       	                   �?@��?.��@u           *�@                            �?�log�@+           `�@                            �?$�C��@�           ��@������������������������       �v��f�@�            �@������������������������       �I,���@=           �}@                            @Tay�f�@g           ��@������������������������       �/�!c
@q            `f@������������������������       �Uk���@�           ��@
                          �@@<���oe@J            @Y@                            @x�k_o@'            �J@������������������������       �,Q�o�@             8@������������������������       �e�t?@             =@                           �?z��'�@#             H@������������������������       ���H �@             1@������������������������       ���=��@             ?@                           �?�,4�@;           К@                          �4@C���f@t           x�@                            �?��)R
@�            �v@������������������������       ����3@0            @Q@������������������������       ��cǰ�	@�            `r@                           �?�6H@r_@�            �l@������������������������       ��mG��@O            �`@������������������������       �L�q�\�
@:            �W@                           @��tSu�@�           ��@                           @�(v��@�           ��@������������������������       �x��g��@�            �t@������������������������       ��~���@�            �x@                          �6@G*x�P@�            �x@������������������������       ��Ջ3@�            `o@������������������������       �4h�ۍ@Z            �b@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       pu@     �^@      V@     �t@     �B@      ~@      *@     �k@      >@      }@     @]@     �K@      =@     �N@     �m@     @T@     @x@     �r@      z@     �W@      f@     �T@      P@     �g@      <@     @j@      *@     `b@      ;@     �k@      V@     �D@      2@     �I@      a@     �O@      i@     �f@     �h@     �P@      e@     �Q@     �K@     �f@      8@     �i@      *@     @a@      ;@     @k@     �U@     �C@      ,@     �G@     �`@      K@      h@     @e@     @h@     @P@     �S@      G@      :@     �Z@      @     �W@      $@      L@      .@      ^@     �F@      8@       @      5@     �R@      6@     �V@      T@     �^@     �D@     �@@      6@       @     �O@      @      I@      @      E@      $@      N@      2@      3@      @      0@     �A@       @     �K@      H@     �R@      ?@      G@      8@      2@      F@              F@      @      ,@      @      N@      ;@      @      @      @      D@      ,@     �A@      @@      H@      $@     �V@      9@      =@     �R@      3@      \@      @     �T@      (@     �X@     �D@      .@      @      :@      M@      @@     �Y@     �V@     �Q@      8@      (@       @      �?      6@      @      7@              $@             �@@      @                      @      "@       @      4@      3@      &@       @     �S@      7@      <@      J@      ,@     @V@      @      R@      (@     @P@     �B@      .@      @      6@     �H@      >@     �T@     �Q@      N@      6@       @      &@      "@      @      @      @              "@               @       @       @      @      @      @      "@       @      &@       @       @      @      @       @      @       @      @              @               @                       @                      "@      @      "@       @       @              �?       @                       @              @              �?                                              "@       @      �?       @      �?      @      @              @       @      �?                              �?                       @                              @       @              �?      @      @      @      @       @      �?              @                       @       @       @      @      @               @       @                       @              @      �?                              @                       @                              �?                      �?                      @      @       @      @       @      �?              �?                               @       @      @       @               @      �?                     �d@     �D@      8@     �a@      "@      q@             �R@      @     �n@      =@      ,@      &@      $@      Y@      2@     �g@     �^@     �k@      ;@     �K@      @      $@      K@      @     �_@              <@      �?      Q@       @      @              @      ?@      @     �L@      F@     �S@      $@     �@@      �?       @      <@      �?     @V@              3@      �?     �D@       @      @              @      (@      @     �@@      9@     �O@      @      @              �?      @              &@              @      �?      "@      �?                               @       @      @      @       @              :@      �?      �?      6@      �?     �S@              .@              @@      �?      @              @      @      �?      <@      3@     �K@      @      6@      @       @      :@       @      C@              "@              ;@               @               @      3@      �?      8@      3@      0@      @      ,@      @      @      ,@       @      :@              @              2@                              �?      *@      �?      @      $@      @      @       @      �?      @      (@              (@              @              "@               @              �?      @              3@      "@      "@             �[@      A@      ,@     @V@      @      b@             �G@       @      f@      ;@       @      &@      @     @Q@      ,@     ``@     �S@     �a@      1@      M@      4@      &@     @Q@      @     �W@              :@      �?     @_@      5@      @      $@      @      G@      @      S@     �A@     �Y@      &@      2@      $@             �E@      @      I@              $@      �?     �F@      "@      @      @       @      9@      @      A@      ,@      H@      @      D@      $@      &@      :@      �?      F@              0@              T@      (@              @       @      5@              E@      5@     �K@      @     �J@      ,@      @      4@       @     �I@              5@      �?     �I@      @      �?      �?      �?      7@      "@     �K@     �E@      C@      @      0@       @      @      (@              G@              *@      �?     �C@       @      �?      �?              ,@      @     �B@      ?@      5@      @     �B@      @               @       @      @               @              (@      @                      �?      "@      @      2@      (@      1@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ&�U<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@x�F��@�	           ��@       	                    �?z��ib�@�           �@                           �?K�]2�@
            �@                           @}��E"�@�            Pu@������������������������       ��aiw�@�             p@������������������������       � ��<?@0            �T@                          �2@r�����@;           �~@������������������������       ���� 0@k            �d@������������������������       �H�@�            pt@
                          �2@�,��@�           Ș@                           �?�	L�@�           �@������������������������       �,)�r��
@�             t@������������������������       �u3��X@           |@                           �?��s�@�           x�@������������������������       ��6�Y�@�            `v@������������������������       ���ACX�@           �|@                            @S�ANR�@�           \�@                           �?b���Z@�           �@                          �<@��,�@           @x@������������������������       ��MrN�@�            �r@������������������������       �CRAR�@:             W@                           @=�#)M�@�           ��@������������������������       �嬘*�@           �|@������������������������       �h�f�_@q            �f@                           �?�T�lD@#           P}@                           �?�ȅ�i@^             d@������������������������       ���ADr@             H@������������������������       �A����@D            @\@                           @�na;�9@�            @s@������������������������       �MSH���@�            �j@������������������������       ���pJ�@7            �W@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       `t@     �c@     �U@     0v@      <@     @}@      "@     �l@      ?@     �z@      [@     @R@     �A@      M@     �p@     �O@     �w@     Pt@     �y@     �Q@     �f@      V@     �E@     �k@      ,@     w@      �?     �`@      (@     �q@     �H@     �I@      &@      5@     �a@      ;@     �n@     @i@     �q@      E@      S@     �E@      8@     �R@      "@     �W@      �?     �K@      @     �R@      3@      <@      @      $@     �H@      $@     @R@      T@     �T@      3@     �D@      0@      &@     �A@      �?      E@              6@      @      7@      "@      @              �?      "@      "@      ;@      =@     �G@      $@      ?@      &@      "@      >@      �?      =@              0@      @      2@      @      @                       @      "@      4@      1@      A@      "@      $@      @       @      @              *@              @              @       @                      �?      �?              @      (@      *@      �?     �A@      ;@      *@      D@       @     �J@      �?     �@@      @     �I@      $@      6@      @      "@      D@      �?      G@     �I@     �A@      "@      @       @      @      ,@       @      .@      �?      &@              0@       @       @      �?       @      7@      �?      @      3@      4@      @      >@      3@       @      :@      @      C@              6@      @     �A@       @      ,@       @      @      1@             �C@      @@      .@      @      Z@     �F@      3@      b@      @      q@             �S@      @     `j@      >@      7@       @      &@     �W@      1@     �e@     �^@     �h@      7@     �H@      4@      &@     �R@       @      `@             �E@             @]@      @      *@      @       @      :@      &@      U@      L@      [@      $@      9@      �?      @      =@       @      R@              *@             �A@       @      @              @      @       @     �@@      8@     �L@      @      8@      3@      @      G@             �L@              >@             �T@      @      "@      @      @      4@      "@     �I@      @@     �I@      @     �K@      9@       @     �Q@      @      b@             �A@      @     �W@      9@      $@      @      @      Q@      @     �V@     �P@     �V@      *@     �@@      .@              =@              Q@              ,@              I@      *@      �?       @      @      9@      @      :@      7@     �G@      @      6@      $@       @     �D@      @     @S@              5@      @      F@      (@      "@       @             �E@      @      P@     �E@     �E@      @     @b@     �Q@     �E@     �`@      ,@     �X@       @      X@      3@     �a@     �M@      6@      8@     �B@     �_@      B@     �`@     �^@     @`@      =@     @X@      G@      <@      Y@      $@      T@      @      O@      @      Z@      B@      *@      2@      4@     @X@      ;@     @W@      R@      X@      2@     �B@      &@      (@      I@      @      B@      @      4@      @      C@      .@      �?       @      �?      E@      $@      >@      >@      7@       @      ?@      @      "@     �G@      @      8@      �?      4@      @      @@      @      �?      @      �?      ?@      @      :@      8@      1@      @      @      @      @      @       @      (@      @              �?      @      $@              @              &@      @      @      @      @       @      N@     �A@      0@      I@      @      F@              E@             �P@      5@      (@      $@      3@     �K@      1@     �O@      E@     @R@      $@      ?@      ?@      $@     �D@      @     �@@             �B@              K@      ,@      $@      @      $@     �D@      &@     �B@      <@     �H@      $@      =@      @      @      "@              &@              @              (@      @       @      @      "@      ,@      @      :@      ,@      8@             �H@      9@      .@     �A@      @      3@      @      A@      ,@     �C@      7@      "@      @      1@      =@      "@      E@     �I@      A@      &@      2@      "@      @      (@              @      @       @       @      6@      @      @       @       @      @       @      .@      8@      .@      @      @       @               @              @      @      @              @      @      @                      @              �?      @      @      @      *@      @      @      $@                              @       @      3@       @       @       @       @      �?       @      ,@      1@      &@              ?@      0@      &@      7@      @      0@      �?      :@      (@      1@      2@      @      @      .@      7@      @      ;@      ;@      3@      @      .@      @      $@      1@      �?      *@      �?      2@      (@      @      .@      @       @      (@      2@      @      8@      5@      $@      @      0@      $@      �?      @      @      @               @              (@      @               @      @      @      @      @      @      "@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ6	<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��kuL�@�	           ��@       	                   �5@�7��̧@�           ī@                           �?|F�=g@�           D�@                          �1@�]<�+@�            �@������������������������       ��!n�	@�            �m@������������������������       �>dc�@`           ��@                            �?bҬ!G�@�           4�@������������������������       �����CG@�             v@������������������������       �O�
�}�@           h�@
                           �?tJ ��@           D�@                            @���,�P@�           �@������������������������       ��k�QE@           z@������������������������       �[)�	�@{             h@                           �?���=�@�           ��@������������������������       ���L:��@d            �c@������������������������       ��I0��@!           ��@                           @����^@�            pv@                           �?�z�N@�             r@                          �6@�u�ݨ@>             [@������������������������       �B-j�	@$             O@������������������������       �m�3,d	@             G@                           �?����@s            �f@������������������������       �Jf�¸^@;             W@������������������������       ��D	�<�@8            �V@                           �?qi�Q�a@,            @Q@                            �?�t�l7@            �D@������������������������       �J�g�W��?             ,@������������������������       ��F���@             ;@                          �3@�1�g:�@             <@������������������������       �=��,@	             $@������������������������       �����w@             2@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �r@     �c@     �V@      u@     �D@     �~@      @     `k@      5@     0}@     @]@     �Q@     �E@     �P@      j@     �R@     0v@     Pr@     �}@      U@      p@     �`@     �U@     �s@      A@     P|@      @     �h@      5@     �z@      X@     �P@      C@      O@     �g@      N@     Pt@      p@     �{@     �T@     �`@     �G@      B@     �f@      $@     Pq@             �^@      @     �o@      D@     �G@      *@      1@      W@      8@     �d@     �b@     �q@     �D@      Q@      0@      1@     �P@      @     @_@             �K@      �?     @]@      *@       @      �?      @     �A@       @      N@      J@     �\@      $@      &@              @      4@       @      G@              ,@             �D@       @      �?              �?      ,@       @      *@      6@     �E@      �?     �L@      0@      ,@      G@      @     �S@             �D@      �?      S@      &@      @      �?      @      5@             �G@      >@     �Q@      "@     @P@      ?@      3@     �\@      @      c@             �P@      @      a@      ;@     �C@      (@      $@     �L@      6@     @Z@     @X@     @e@      ?@      (@      .@      @      >@             �H@              .@      @      H@      @      "@      @      �?      (@       @      ?@      6@      O@      2@     �J@      0@      ,@      U@      @     �Y@              J@       @     @V@      5@      >@      @      "@     �F@      ,@     �R@     �R@      [@      *@     �^@     �U@     �I@     `a@      8@      f@      @     �R@      .@      f@      L@      4@      9@     �F@      X@      B@      d@     �Z@     �c@      E@     �G@      2@      9@      D@      @     �R@              9@      @     @P@      :@      $@      (@      .@      H@      $@     �R@     �E@     �D@      7@     �C@      (@      0@      @@      @      O@              ,@             �E@      "@      @      (@      @      A@      @     �H@      =@     �@@      *@       @      @      "@       @      @      *@              &@      @      6@      1@      @              $@      ,@      @      :@      ,@       @      $@      S@      Q@      :@     �X@      2@     @Y@      @     �H@      $@     �[@      >@      $@      *@      >@      H@      :@     @U@      P@     �]@      3@      "@      $@      &@       @              1@       @      @              1@      @       @      �?       @      @      @      3@      &@      :@      @     �P@      M@      .@     �V@      2@      U@      @     �E@      $@     �W@      ;@       @      (@      <@      E@      7@     �P@     �J@      W@      0@     �D@      7@      @      3@      @     �C@              7@             �B@      5@      @      @      @      5@      ,@      >@     �B@      >@      �?      @@      2@      @      0@      �?      C@              *@              ?@      3@      @      @      @      3@      ,@      7@      =@      5@      �?      4@      @       @       @      �?      ,@              @               @      "@      @              �?      @      @      @      .@       @              @                      @              &@              @              @       @      @                       @       @      @      .@      �?              .@      @       @       @      �?      @                              @      �?                      �?      @      @      @              �?              (@      *@      �?       @              8@              $@              7@      $@      �?      @      @      *@      "@      1@      ,@      3@      �?      @      @      �?      @              0@              @              &@              �?      @      @      @      @      "@      "@      @      �?       @      @               @               @              @              (@      $@                              $@      @       @      @      (@              "@      @              @      @      �?              $@              @       @              �?               @              @       @      "@              @      @              �?      @                      $@              �?       @                                              @       @      @                      @                       @                      @                                                                                       @              @                      �?      @                      @              �?       @                                              @       @      @              @                       @              �?                              @                      �?               @              @      @      @                                       @              �?                               @                                                      �?       @       @              @                                                                      @                      �?               @               @      @       @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��X@hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@	/J��@�	           ��@       	                    �?�}gr@s            �@                           �?� `Tn@           P�@                          �1@Ai��O�@L            �Y@������������������������       ��}��S(@$             G@������������������������       �|B8��	@(            �L@                            @ j��
@�           �@������������������������       �K ���@
@O           ��@������������������������       ��+�
n@u            �e@
                           @�@Y��@c           ��@                           �?���Ҩ�@�           ��@������������������������       ��|��B9@�            �u@������������������������       ��kj��@�            �o@                           �?)J��vd@�            pt@������������������������       ���B#�@Q            @^@������������������������       �e�08�@�            �i@                           �?�����|@U           �@                           @��k~@�           ��@                            @A��;	/@�           ��@������������������������       ��*���@�            �v@������������������������       ���j��@�            �p@                           �?Ύ��@            |@������������������������       ����u��@Q            @_@������������������������       ����}-@�            Pt@                          �;@��j@�           $�@                           �?�74�?@M           �@������������������������       �il�W�6@$           }@������������������������       ��!�ҟ@)           }@                            �?o�����@e            �d@������������������������       ����
@<            �X@������������������������       ���0W:�@)            @Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@     @b@     @V@      s@      C@     P~@      $@     �l@     �B@     pz@     �W@     �H@      ?@      S@     �o@      P@     �w@     �r@     �}@     @S@     �a@     �A@     �C@     �`@      &@     �n@       @     �W@      (@     �k@     �@@      4@      @      "@     �\@      0@     �d@      _@     @q@     �C@     @Q@      .@       @     �N@       @     �`@              H@             @[@      $@      @       @      @      D@      @     @R@      N@     �b@      1@      @              @      @      �?       @              @               @      @                       @      "@      �?      @      @      ;@      @      @              @      �?      �?      @              �?              @      @                       @       @      �?      �?      @      &@              @              �?      @              @              @              @      @                              @              @      �?      0@      @      O@      .@       @     �K@      �?      _@              F@             @Y@      @      @       @      �?      ?@      @     �P@     �J@      _@      *@     �A@      &@      �?     �B@              Y@              >@              S@      �?      @       @      �?      :@      @     �K@     �D@     �Y@      @      ;@      @      �?      2@      �?      8@              ,@              9@      @       @                      @              &@      (@      6@      @     @R@      4@      ?@     �R@      "@     �\@       @      G@      (@     @\@      7@      ,@      �?      @     �R@      (@     �V@      P@     @_@      6@     �H@      $@      :@     �L@      "@      I@       @      5@      $@      Q@      7@      $@              @     �H@      $@     �M@      F@     �S@      1@      >@      @      5@      :@       @      6@       @      ,@      $@     �B@      "@      @              @     �@@      @      4@      :@     �H@      ,@      3@      @      @      ?@      �?      <@              @              ?@      ,@      @               @      0@      @     �C@      2@      >@      @      8@      $@      @      1@              P@              9@       @     �F@              @      �?              9@       @      @@      4@      G@      @      *@              @      @              8@              (@       @      1@                                      @              (@      "@      6@              &@      $@       @      ,@              D@              *@              <@              @      �?              5@       @      4@      &@      8@      @     �i@     �[@      I@     `e@      ;@     �m@       @     �`@      9@      i@      O@      =@      <@     �P@     �a@      H@     �j@     `f@     �h@      C@      U@     �P@      ?@     @U@      ,@      W@      @     �S@      ,@      S@      <@      4@      6@      H@     �Q@      ;@      Y@      X@     �Y@      3@     �E@      B@      8@      J@      @      N@      @     �J@      @     �B@      ;@      (@      (@      A@      A@      &@      L@      J@     �J@      .@      ;@      5@      &@      8@      @      H@      @      ?@      �?      <@       @       @      $@      ,@      3@      @      B@      .@     �A@       @      0@      .@      *@      <@      �?      (@      �?      6@      @      "@      3@      @       @      4@      .@      @      4@     �B@      2@      @     �D@      ?@      @     �@@       @      @@              9@      @     �C@      �?       @      $@      ,@     �B@      0@      F@      F@     �H@      @      6@      @      @       @       @      @              @              "@              �?      @      @      ,@      @      *@      3@      $@              3@      <@       @      9@      @      <@              4@      @      >@      �?      @      @      $@      7@      *@      ?@      9@     �C@      @      ^@      F@      3@     �U@      *@     `b@       @     �L@      &@     @_@      A@      "@      @      3@     �Q@      5@     �\@     �T@     @X@      3@     �X@     �C@      &@     �T@      "@     �_@             �K@      &@      Y@      =@      "@      @      1@     �P@      2@     �X@     �R@     �P@      0@      J@      (@      @      B@      "@     @Q@             �@@      &@     �F@      0@       @              @     �A@      $@     �E@      A@     �B@       @      G@      ;@      @     �G@              M@              6@             �K@      *@      @      @      &@      ?@       @      L@      D@      =@       @      6@      @       @      @      @      4@       @       @              9@      @              @       @      @      @      0@      "@      ?@      @      "@      @       @               @      ,@               @              &@      @                       @      �?       @      $@      @      <@      �?      *@      �?      @      @       @      @       @                      ,@                      @              @      �?      @      @      @       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJɅ�chG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����9�@�	           ��@       	                    �?��=+�@           T�@                          �:@�=�T@h            �@                           �?>��_�@1           �|@������������������������       ��ǵ+��@|             h@������������������������       �O]\g@�            �p@                          �?@0N��Y�@7            @U@������������������������       ��C-C�8@)            �P@������������������������       ���p��@             3@
                          �?@��R��@�           Đ@                            @+Y/���@�           �@������������������������       ��;���4@u           �@������������������������       ����iR@           �y@                           �?�c+)�[@0             T@������������������������       �}c���@             :@������������������������       �����	@"             K@                          �6@��H�g@�           �@                           �?sGΔ`|@�           ��@                           @8!T�tM@t           �@������������������������       ������@�            �j@������������������������       ���Z�!
@�            �v@                           @�z���@l           ��@������������������������       �����<@           @z@������������������������       �J�P���@d           ؁@                          �8@2�]��@�           ��@                           @��
ѭ@�            �q@������������������������       �2J � �@�            @j@������������������������       �(#+��j	@1            �R@                            @�|��@           `{@������������������������       �[�7��@�            �v@������������������������       ��E�w@0             S@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@      c@      S@     �u@      :@     @      @     �l@      :@     Pz@     �]@      O@      >@     �T@      m@     @Q@      v@     �r@      }@      S@     �`@     �R@      J@     �c@      1@      b@      @     �[@      2@      b@     �H@      B@      2@      K@      X@      @@      a@      `@     �e@      D@      O@      *@      4@     �A@      @     �G@       @      C@      @     �J@      0@      *@      @      ,@     �@@      @     �G@      L@     �P@      $@      M@      $@      (@      @@      @      G@       @      :@             �I@      (@      *@              "@      ;@      @     �C@      I@      L@      $@      0@      @       @       @              =@              *@              ?@       @      @              @      $@              4@      7@      5@      @      E@      @      $@      8@      @      1@       @      *@              4@      $@      "@              @      1@      @      3@      ;@     �A@      @      @      @       @      @              �?              (@      @       @      @              @      @      @      �?       @      @      &@              @       @      @       @              �?              @      @       @      @               @      @      @               @      @      &@              �?      �?      �?      �?                              @                                      @       @              �?                                     @R@     �N@      @@     �^@      (@     �X@       @      R@      ,@     �V@     �@@      7@      &@      D@     �O@      :@     �V@     @R@     �Z@      >@     �Q@     �F@      ;@     @]@      (@     �U@       @     �P@      ,@     �U@     �@@      5@      $@      B@      O@      9@      V@     �N@      Z@      9@      G@      ;@      &@      T@      @      G@             �@@       @      N@      4@      (@      @      .@      ?@      *@     �F@     �A@     �P@      3@      8@      2@      0@     �B@      @     �D@       @      A@      @      ;@      *@      "@      @      5@      ?@      (@     �E@      :@      C@      @      @      0@      @      @              &@              @              @               @      �?      @      �?      �?       @      (@       @      @      �?      @      �?       @              @              @              �?              �?              @      �?              �?                               @      (@      @      @              @                              @              �?      �?                      �?      �?      (@       @      @      j@     �S@      8@      h@      "@      v@      �?     @^@       @     Pq@     @Q@      :@      (@      =@      a@     �B@      k@     �d@     0r@      B@      \@      E@      (@     @`@      @     �q@             �U@      @     �g@      D@      7@      @      "@      X@      6@     �c@     �Z@     `l@      6@      F@       @      @      D@       @     �_@              >@      �?     �R@      (@      @              @      A@      @     �E@     �B@      X@      .@      $@      @      �?      1@             �D@              "@              7@      @      @               @      ,@      �?      9@      1@      ;@      (@      A@      @      @      7@       @     @U@              5@      �?     �I@      @                      @      4@       @      2@      4@     @Q@      @      Q@      A@      @     �V@      �?     �c@              L@       @      ]@      <@      4@      @      @      O@      3@     �\@     @Q@     ``@      @      7@      3@      @     �C@      �?     �L@              5@              K@      .@       @       @       @      @@      3@     �J@      9@      F@      �?     �F@      .@       @     �I@             �X@             �A@       @      O@      *@      (@      @       @      >@             �N@      F@     �U@      @     @X@      B@      (@      O@      @     �Q@      �?     �A@      @     �U@      =@      @      @      4@     �D@      .@      N@     �N@      P@      ,@      F@      5@       @      4@              8@              2@      �?     �C@      *@                      "@      &@      @      9@      A@      &@      @     �D@      ,@       @      &@              2@              2@      �?      5@      *@                      @      "@      @      2@      5@      "@      @      @      @              "@              @                              2@                              @       @      �?      @      *@       @       @     �J@      .@      $@      E@      @      G@      �?      1@      @      H@      0@      @      @      &@      >@       @     �A@      ;@     �J@       @      F@      &@       @      C@      �?      F@      �?      *@      @      B@      0@              @       @      <@      @      ;@      7@     �F@      @      "@      @       @      @      @       @              @              (@              @      �?      @       @      @       @      @       @       @�t�bub�s     hhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJHN�JhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@����@�	           ��@       	                    @��v�P�@u           8�@                           �?��A8@           ��@                            �?�c�kR@�            �v@������������������������       ��hG��
@w             h@������������������������       ��R�J@p            �e@                           �?]<��d@'           �~@������������������������       �bf�hC@�            �r@������������������������       ��I���@}             h@
                            @|��id@g           ��@                           @xa,�}
@1           0}@������������������������       ��~V�7�@u             g@������������������������       ���b��
@�            �q@                           �?ڪ�d@6            �W@������������������������       ������@            �M@������������������������       �=P�/@             B@                            @)�6rb@           v�@                           �?Hd�f�@V           ��@                           �?;�-BN�@�            �@������������������������       ��� �x@�             o@������������������������       �<�(a�	@*           �|@                           �?�� Q�@�           ��@������������������������       ���zI�1@�            �w@������������������������       �����cZ@�           p�@                           �?�����@�           p�@                           @SP\�� @�             p@������������������������       �� ݣ�@o            �f@������������������������       ��w�PEk
@4             S@                           @��D��@$           �|@������������������������       ������@�            �s@������������������������       ����#4@X            �a@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        t@      ]@     @U@     @v@      H@     �~@       @     �m@      6@     �z@     �[@     �L@      G@      M@     �k@      N@     pw@     �t@     p|@     @U@     @\@      7@      <@      b@      @     �j@             �T@             �e@     �@@      3@       @      .@      O@      *@     �`@     �]@     �j@      6@     �N@      &@      6@     �Y@       @     @[@             �E@             �[@      @@      (@      @      *@     �F@      "@     @V@     @T@     �Y@      ,@      =@      @      @      E@      �?     �H@              9@             �M@      *@      @      @      @      *@              @@      :@      J@      @      &@      @      @      7@              1@              &@              D@      @       @       @              "@              1@      (@     �B@       @      2@      �?       @      3@      �?      @@              ,@              3@      "@       @      �?      @      @              .@      ,@      .@       @      @@      @      1@      N@      �?      N@              2@             �I@      3@       @               @      @@      "@     �L@     �K@      I@      $@      7@      @      ,@     �@@      �?      ?@              *@              6@       @      @              @      4@       @      7@     �G@      D@       @      "@       @      @      ;@              =@              @              =@      &@      �?              @      (@      @      A@       @      $@       @      J@      (@      @      E@       @     �Y@              D@             @P@      �?      @      @       @      1@      @      G@     �B@     @\@       @      C@       @      @      B@      �?      U@              ?@              M@              @      @              *@      @      D@      A@      Y@       @      1@               @      5@              B@              @              1@              @      �?              @      �?      ,@      "@      I@       @      5@       @       @      .@      �?      H@              8@             �D@                      @              $@       @      :@      9@      I@      @      ,@      @       @      @      �?      3@              "@              @      �?      @               @      @      �?      @      @      *@               @              �?      @      �?      2@              @              @                                       @              @      @      "@              @      @      �?      �?              �?              @              @      �?      @               @       @      �?                      @             �i@     @W@     �L@     �j@      F@     �q@       @     `c@      6@     `o@     @S@      C@      C@     �E@      d@     �G@      n@      k@      n@     �O@     `b@      L@     �A@     �d@      8@     @k@      @     @V@      ,@     �h@      J@      8@      ;@      @@      [@     �@@     `f@     `a@     �f@     �G@      F@      :@      .@     �R@      $@      N@      @      J@      @     �T@      5@      ,@      $@      4@     �B@      4@     �P@     �H@     �P@      <@      &@      @      @      4@       @      7@      @      5@      �?     �A@      @      �?      @      @      ,@      @      ?@      5@      5@      1@     �@@      7@      $@      K@       @     �B@      �?      ?@      @     �G@      .@      *@      @      1@      7@      0@     �A@      <@     �F@      &@     �Y@      >@      4@     �V@      ,@     �c@             �B@      @     �\@      ?@      $@      1@      (@     �Q@      *@     @\@     �V@     �\@      3@      @@      (@      &@      A@      �?     �K@              4@              B@      @               @      �?      4@             �I@     �B@      I@      &@     �Q@      2@      "@     �L@      *@     �Y@              1@      @     �S@      9@      $@      .@      &@     �I@      *@      O@     �J@      P@       @      N@     �B@      6@     �G@      4@      O@      �?     �P@       @      K@      9@      ,@      &@      &@      J@      ,@     �N@     @S@      N@      0@      @@      @      (@      0@      @      3@      �?      8@      @      8@      @      @       @      @      .@      @      &@      >@      >@      @      8@      @      &@      ,@      @      &@      �?      5@      @      "@      @      @       @      @      @      @      @      8@      2@               @              �?       @      @       @              @              .@                                       @              @      @      (@      @      <@      ?@      $@      ?@      ,@     �E@              E@      @      >@      2@       @      "@      @     �B@      "@      I@     �G@      >@      &@      .@      3@      "@      ;@      *@      =@              <@       @      .@      ,@      @      @      @      8@       @     �A@      B@      0@      "@      *@      (@      �?      @      �?      ,@              ,@      @      .@      @       @       @      �?      *@      �?      .@      &@      ,@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ 2hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @Nb%|J�@�	           ��@       	                    @� �-@           ��@                          �4@ȑb;�@G           ؚ@                           @��f��C@�           h�@������������������������       ���N/�@f           �@������������������������       ��H��1�@g            `e@                           �?�{P�tK@z           H�@������������������������       �m��rH@           �@������������������������       ���Q�z@�            �x@
                           @�w��@�           �@                          �0@ΰ#�@�           ��@������������������������       ����h�@&            �R@������������������������       �\@�{)@�           X�@                          �6@ Ò8�@�            w@������������������������       �fRn��X@�            `m@������������������������       �����c@]            �`@                           �?�� Xi@�           4�@                          �6@o�:��@�           ��@                           �?��;��i@�             x@������������������������       ���,��,@D            @]@������������������������       ��r\�U5@�            �p@                           @߳��@�            �s@������������������������       ��au8��@�            �k@������������������������       �AYQh�<@?            �V@                           @Z�`�e@           Py@                           @*�ld�@�             o@������������������������       �,�B+�.@u            �e@������������������������       ���T���
@1            �R@                           �?'�W�_w@f            �c@������������������������       � �n���
@5            �T@������������������������       ��%J/�@1            �R@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        s@      `@      X@     `v@     �E@     �@      @     �m@      ;@     �{@     @W@      P@      A@      R@     �o@     �S@     �u@     �t@     pz@      Q@     �j@     �V@      I@     �p@      5@      y@      @     �c@      2@     `u@      M@     �D@      9@     �H@     �g@      K@     �m@      k@     `t@      I@     �_@      O@      >@      f@      1@      j@      @     �X@      @     `i@      E@      =@      (@      D@      `@      F@     �a@     �`@      f@      D@      E@      (@      4@     �T@      @     @X@              <@      �?      W@      .@      &@       @      @     �M@      $@     �N@     �M@     @W@      6@      =@      $@      $@      O@      �?     �R@              2@      �?     @S@      $@      &@       @      @     �H@       @      J@     �A@     �Q@      6@      *@       @      $@      5@       @      6@              $@              .@      @                      @      $@       @      "@      8@      6@             @U@      I@      $@     �W@      ,@     �[@      @     �Q@      @     �[@      ;@      2@      $@     �@@     �Q@      A@      T@     @R@      U@      2@      @@      <@      @      P@      "@     �O@      @     �K@      @     �N@      (@      .@      @      0@     �D@      4@      I@     �F@     �O@      "@     �J@      6@      @      >@      @      H@              .@      �?      I@      .@      @      @      1@      =@      ,@      >@      <@      5@      "@     @U@      <@      4@     @W@      @     @h@             �M@      (@     `a@      0@      (@      *@      "@      N@      $@     @X@      U@     �b@      $@     �L@      .@      0@     �N@             �`@              H@      @     �\@      @      @      &@      @     �A@      �?     �J@     �G@     �Y@      "@      @              @      @              8@              �?               @                                      @              $@              $@             �I@      .@      $@      L@             �[@             �G@      @     �Z@      @      @      &@      @      ?@      �?     �E@     �G@     @W@      "@      <@      *@      @      @@      @      N@              &@      "@      9@      "@      @       @      @      9@      "@      F@     �B@      G@      �?      ,@      "@      @      5@             �I@              @       @      0@      @      @      �?              ,@      @      ?@      ,@      >@      �?      ,@      @      �?      &@      @      "@              @      �?      "@      @              �?      @      &@      @      *@      7@      0@              W@     �C@      G@      V@      6@     �Z@              T@      "@      Y@     �A@      7@      "@      7@     �P@      9@     �Z@     @]@     @X@      2@     �F@      6@      E@      J@      5@     �G@              L@      "@     �F@      8@      0@      @      5@      F@      ,@     �P@      W@     @P@       @      ;@      ,@      3@      :@      .@     �C@              ;@      �?      =@      2@      @              @      ;@      @     �B@     �I@     �B@      �?      &@      @      @      $@      �?       @              @      �?      &@      @                      �?      &@       @      @      1@      0@              0@       @      (@      0@      ,@      ?@              5@              2@      *@      @              @      0@      �?     �@@      A@      5@      �?      2@       @      7@      :@      @       @              =@       @      0@      @      $@      @      ,@      1@      &@      =@     �D@      <@      @       @      @      4@      8@      �?      @              6@       @      @      @      @      @      "@      $@       @      8@     �A@      .@      @      $@      @      @       @      @       @              @              (@              @      @      @      @      @      @      @      *@             �G@      1@      @      B@      �?     �M@              8@             �K@      &@      @       @       @      6@      &@      D@      9@      @@      $@      ?@      @              5@      �?      E@              4@              8@      $@       @               @      *@      @      5@      3@      7@      "@      8@      @              &@      �?      ?@              *@              4@      $@       @                      @      @      2@      *@      *@       @      @      @              $@              &@              @              @                               @      $@              @      @      $@      �?      0@      $@      @      .@              1@              @              ?@      �?      @       @              "@      @      3@      @      "@      �?      &@       @      �?      &@              @               @              1@              @                       @      @      @      @      @              @       @      @      @              &@               @              ,@      �?               @              @      @      (@      @      @      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��OhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�ۗ�@�	           ��@       	                    �?����@=           d�@                            �?�|<��S@�           ��@                           @ỹ`IN@           �y@������������������������       ��O�4�n@�             m@������������������������       ���Yߕ	@q            �f@                           @i�����@�            ps@������������������������       ��?��@^            �b@������������������������       ��rJ �i@i            @d@
                            �?� ��b1@n           (�@                           @/���
�@�            �q@������������������������       ��À�f�@Z            �`@������������������������       �K$�#@`             c@                          �9@���#��@�           @�@������������������������       ��a�p�@\           @�@������������������������       ��D�[�@X             `@                          �6@Mn�I�@c           `�@                            �?-w��2@#           H�@                           �?�R�~@�            �w@������������������������       �H��@/            �Q@������������������������       ����1@�            `s@                           @��uP�@7           ��@������������������������       ��m|��@.           `~@������������������������       ��5-�\@	            {@                           @���uf�@@           ��@                           �?Q�,���@�           ��@������������������������       ���t�;0@�            �y@������������������������       �T��vC@�            �n@                          �:@?ݝd��@�            �p@������������������������       ��!Fq�@W            �b@������������������������       �'P�zX�@I            @]@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     @^@     �U@     �v@      ?@     �~@      @     @m@     �@@     �z@     �[@      L@     �F@     �S@     p@     �O@     �v@     �r@     p{@     �V@      b@     �@@      <@     �a@      1@      n@       @     @X@      $@     �i@     �J@      5@      ,@      6@     �Y@      4@     �a@     �a@     `i@      H@      J@      ,@      ,@     �E@      @     �Z@             �H@       @     @Y@      7@      $@      @      .@     �I@      �?     �H@      O@     @Y@      8@      8@      (@      "@      5@      @     �P@              8@              S@      "@      @      �?      @      8@      �?      >@      >@      O@      "@      0@      @      @      ,@      �?      9@              ,@             �B@      @      @      �?      @      2@      �?      0@      3@     �A@      "@       @      @      @      @       @      E@              $@             �C@      @      �?                      @              ,@      &@      ;@              <@       @      @      6@      �?     �C@              9@       @      9@      ,@      @       @      $@      ;@              3@      @@     �C@      .@      $@       @      @      (@              0@              0@       @      *@      $@       @       @       @      (@              &@      ,@      "@      @      2@                      $@      �?      7@              "@              (@      @       @               @      .@               @      2@      >@      $@     @W@      3@      ,@      Y@      *@     �`@       @      H@       @      Z@      >@      &@      &@      @      J@      3@      W@     @T@     �Y@      8@      8@      $@      @      9@       @     �@@       @      .@             �A@      @      @      @      @      5@      @      :@      ;@      <@       @      $@      @       @      @      �?      9@       @      @              5@      @      �?      @              @      @      ,@      @      1@       @      ,@      @      @      3@      �?       @              &@              ,@               @       @      @      0@      @      (@      8@      &@      @     @Q@      "@      "@     �R@      &@     �Y@             �@@       @     @Q@      9@       @      @      @      ?@      (@     �P@      K@     �R@      0@      G@      @       @     @Q@      @      X@              ;@      @     �M@      0@      @      �?              9@      &@      I@      J@     �K@      (@      7@      @      �?      @      @      @              @       @      $@      "@      �?      @      @      @      �?      0@       @      3@      @     `e@      V@      M@     @k@      ,@     �o@      @      a@      7@     �k@      M@     �A@      ?@     �L@     @c@     �E@     `k@      d@     �m@     �E@      Z@     �C@      =@     �`@      @     �g@       @     �R@      1@     ``@      ;@      ,@      $@      5@     �T@      ;@      `@     �V@     �b@      7@      <@       @      "@     �J@             �L@              0@      $@      =@      "@      @      @       @      7@      @      8@      7@      O@      $@              �?      �?      $@              $@              @      �?       @      �?      �?      @              @      @      @      @      ,@      @      <@      @       @     �E@             �G@              (@      "@      ;@       @      @      @       @      4@      �?      1@      4@      H@      @      S@      ?@      4@     @T@      @     �`@       @     �M@      @     �Y@      2@      $@      @      3@     �M@      5@     @Z@      Q@     �U@      *@     �D@      9@      0@      F@      @     �N@       @      =@      @      C@      *@       @      �?      1@      C@      @      K@      A@      F@      @     �A@      @      @     �B@      �?     �Q@              >@       @      P@      @       @       @       @      5@      0@     �I@      A@     �E@      @     �P@     �H@      =@      U@      "@     @P@       @      O@      @     �V@      ?@      5@      5@      B@      R@      0@     �V@     @Q@     �U@      4@      H@     �B@      5@      Q@       @     �G@       @     �E@      @     �K@      ;@      3@      0@      5@     �J@      @     �P@     �G@      L@      3@      >@      3@      0@      H@       @      ,@       @     �A@      @      <@      8@      0@      ,@      *@      ?@      @      A@      =@      ?@      .@      2@      2@      @      4@             �@@               @              ;@      @      @       @       @      6@      �?      @@      2@      9@      @      3@      (@       @      0@      @      2@              3@             �A@      @       @      @      .@      3@      "@      8@      6@      ?@      �?      .@       @       @      @      @      $@              @              6@      �?              @      (@      @      "@      3@      &@      *@              @      @      @      $@               @              0@              *@      @       @              @      *@              @      &@      2@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ1�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�@�	           ��@       	                   �1@����a@:           ��@                           �?G���	@�            �p@                           �?������	@0             S@������������������������       ���dr˩@            �@@������������������������       � �tHx�@            �E@                            �?��I�\4@y            �g@������������������������       �М�3=@F            @[@������������������������       �-�)��@3            @T@
                           �?2|��@�           h�@                          �:@�HQ��@           �|@������������������������       �����@�            w@������������������������       �
�(�n�@8             V@                           @?���M@u           ��@������������������������       �m�ج�@m            �f@������������������������       ��XKc@           �y@                          �<@���NO�@|           J�@                           @
�#�@�           8�@                          �4@JV��@�           ��@������������������������       �6>M�G�@�           ��@������������������������       �L亡��@�           ̒@                          �5@��� /@$            �P@������������������������       �N�)6�x@             9@������������������������       ��Q��^@            �D@                          �?@�j��@�            �p@                           @���>˥@Z            �a@������������������������       �po��@'            @P@������������������������       ��[��4@3            �S@                           �?ͅ��@H            �^@������������������������       �a���-�@2            @T@������������������������       ��c�n�@            �D@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �a@     �U@     �t@     �@@     @@      @     �l@      =@     �}@     �W@     �H@      7@      U@     �p@      R@      w@     �r@     �z@     @U@      W@      8@     �B@     �[@      @     �i@              V@      @      e@     �@@      (@      @      0@     �Y@      @      `@     �V@     �b@      A@      0@               @      "@      �?      Q@              3@             �F@       @      �?              @      6@              ,@      9@     �@@      @      $@               @      �?      �?      .@               @              @       @                               @              @      @      (@              @                      �?              @              @               @       @                               @               @      @       @              @               @              �?      $@              @              @                                      @              @      @      @              @                       @             �J@              &@              D@              �?              @      ,@              "@      2@      5@      @      @                      @              4@              @              @@                                      ,@              @      $@      (@       @       @                      @             �@@              @               @              �?              @                      @       @      "@      @      S@      8@     �A@     @Y@      @      a@             @Q@      @      _@      ?@      &@      @      *@     @T@      @     �\@     �P@     �\@      <@      7@      .@      :@      K@      @      E@              C@      @     �G@      3@      $@      @       @      5@      @      M@      >@      D@       @      4@      (@      6@     �D@      @      E@              <@      @      F@      0@      @       @       @      ,@       @      G@      5@     �B@      @      @      @      @      *@                              $@      �?      @      @      @      @              @       @      (@      "@      @      @     �J@      "@      "@     �G@       @     �W@              ?@       @     @S@      (@      �?              @      N@      @      L@      B@     �R@      4@      3@       @      �?      0@              6@               @              8@      @                              2@       @      5@      @      5@      .@      A@      @       @      ?@       @     @R@              7@       @     �J@       @      �?              @      E@      �?     �A@      =@      K@      @     �k@     @]@      I@     �k@      ;@     pr@      @     �a@      7@      s@      O@     �B@      0@      Q@     �d@     @P@      n@     `j@     Pq@     �I@      h@     �V@      D@      j@      5@     �q@      �?      a@      3@     �q@      J@     �B@      (@     �K@      c@     �J@     `k@      g@     �n@      G@     �g@     �U@      D@     `i@      0@     �q@      �?     �`@      3@      q@      J@     �B@      &@     �K@     `b@     �G@     �j@      f@     `m@      G@      Q@      @@      5@      X@      @     �a@      �?      P@      @      b@      <@      1@      @       @      P@      3@      [@      U@     @`@      6@      ^@      K@      3@     �Z@      $@      b@             �Q@      ,@     @`@      8@      4@      @     �G@     �T@      <@      Z@     @W@     @Z@      8@      @      @              @      @                       @               @                      �?              @      @      @      @      (@              @       @              @                               @               @                      �?                              @              @              �?       @                      @                                      @                                      @      @      �?      @       @              <@      ;@      $@      .@      @      $@      @      @      @      6@      $@              @      *@      (@      (@      5@      ;@      >@      @      *@      "@      @      (@      @      @       @      @      @      0@      @              @       @      &@       @      "@       @      4@       @      "@       @       @      @               @       @      �?      @      $@       @              @      @      @      �?      @       @      �?              @      �?      @      @      @      @              @              @      @                      @      @      �?      @      @      3@       @      .@      2@      @      @       @      @      �?       @              @      @              �?      @      �?      $@      (@      3@      $@      @      @      .@      @      @      �?      @               @              @      @              �?      @      �?      @      @      2@      @       @      $@      @                      �?      �?      �?                      �?       @                      �?              @      "@      �?      @      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ|�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�����@�	           ��@       	                     @�r@           ��@                          �3@'�5-@t           �@                           �?M�~u@�           (�@������������������������       �,�xʍ@�            p@������������������������       ���8��@�           H�@                           �?YCHS%@�           Ї@������������������������       �
���>�@�            Pu@������������������������       �Ծ�7@           Pz@
                           �?�F�8	z@�           ��@                          �3@+0.���@�            �t@������������������������       �ޔ-z�@x             f@������������������������       ��x&�W@[            @c@                           �?��(��_@�            �r@������������������������       ��K��g@_            �c@������������������������       ��r�q�@[            �a@                            @g�1:w�@�           <�@                           @�F~�+@�           X�@                          �7@t��{�9@U           8�@������������������������       �^yn3�i@r            �g@������������������������       �?
�Kt@�           H�@                          �9@?ԅ�X�@F            �[@������������������������       ��xl��
@             I@������������������������       ��c*\�/	@(            �N@                           @���=@           �{@                           @��E�@@�            �p@������������������������       �X�|�X@�            `k@������������������������       �]�۲7B	@            �G@                          �<@���x]�@q            �e@������������������������       �s�9,�@W             a@������������������������       ������#
@             C@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       @v@     �a@     @Y@     pv@     �H@     P~@      @     �j@      :@     �{@     �X@      M@     �C@      R@     @n@      K@     �v@     t@     �z@      P@     @j@     �P@      N@     @l@      7@     �w@             �`@      2@     `r@     �G@      ?@      ,@      2@     �a@      5@     @m@      h@     �q@      A@     @_@      I@     �D@     @e@       @     �q@             �W@      2@     �l@      ;@      ;@      $@      0@     �Z@      (@     �e@     `a@     `m@      <@     �O@      9@      .@      Y@      @     `e@             �L@      @      c@      0@      (@      @      @     @P@       @      T@      T@     @d@      (@      1@      "@      $@      @@      �?      ;@              (@      @      9@      @       @               @      .@       @      "@      @@      D@      "@      G@      0@      @      Q@       @      b@             �F@       @      `@      (@      @      @       @      I@      @     �Q@      H@     �^@      @      O@      9@      :@     �Q@      @      ]@              C@      *@     @S@      &@      .@      @      (@     �D@      @      W@     �M@     @R@      0@      9@      1@      @     �A@       @     �O@              $@             �B@      "@      �?      @      @      5@      @     �D@      <@      <@      @     �B@       @      3@     �A@      @     �J@              <@      *@      D@       @      ,@      @      @      4@             �I@      ?@     �F@      (@     @U@      0@      3@      L@      .@     @V@              D@              P@      4@      @      @       @      A@      "@      O@      K@     �I@      @     �H@      @      .@      6@      ,@     �D@              1@              :@      .@      �?      @       @      0@      @      C@      ?@      <@      �?      4@      @      "@      2@      �?      6@               @              $@      (@      �?       @              *@      �?      5@      ,@      3@      �?      =@       @      @      @      *@      3@              "@              0@      @               @       @      @      @      1@      1@      "@              B@      $@      @      A@      �?      H@              7@              C@      @      @                      2@      @      8@      7@      7@      @      6@               @      8@      �?      1@              .@              :@       @       @                      "@       @      $@      @      .@      @      ,@      $@       @      $@              ?@               @              (@      @      �?                      "@      @      ,@      0@       @             @b@     �R@     �D@     �`@      :@     @[@      @     @S@       @     �b@     �I@      ;@      9@      K@     �Y@     �@@     �_@      `@     `a@      >@      Z@     �I@      6@     �W@      3@     �V@      @     �H@      �?     @^@      9@      *@      1@      <@      T@      ;@     �V@     �S@     �[@      3@      V@      E@      6@     �W@      ,@      U@      @      D@      �?     �[@      9@      *@      .@      <@     �Q@      8@     @S@      Q@     �W@      2@      9@      @      �?      =@       @      *@               @              2@       @      �?              @      0@      @      9@      1@      1@      $@     �O@     �C@      5@     �P@      (@     �Q@      @      C@      �?     @W@      7@      (@      .@      6@     �K@      5@      J@     �I@     @S@       @      0@      "@                      @      @              "@              $@                       @              "@      @      *@      &@      1@      �?      @      @                      @                      @              @                       @              @       @      @      @      @              *@      @                              @              @              @                                      @      �?      @      @      (@      �?      E@      8@      3@      C@      @      3@       @      <@      @      =@      :@      ,@       @      :@      6@      @      B@     �H@      <@      &@      6@      .@      *@      1@      @      *@       @      2@      @      &@      5@      &@      �?      ,@      .@      @      2@     �B@      *@      @      ,@      &@      *@      ,@      @      *@       @      2@      @      "@      .@      &@      �?      ,@      &@      @      .@      =@      @      @       @      @              @                                               @      @                              @              @       @      @       @      4@      "@      @      5@              @              $@       @      2@      @      @      @      (@      @              2@      (@      .@      @      4@       @      @      (@              @              $@       @      1@              @      @       @      @              0@      @      (@      @              �?       @      "@              �?                              �?      @               @      @      @               @      @      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ/�l3hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?J��́�@�	           ��@       	                     @�QR�@           T�@                          �7@~2)"��@T           �@                           �?*�2��@_           �@������������������������       ���� �@            `j@������������������������       ��\`S�@�            �v@                          �:@�z���@�            Pv@������������������������       ��+ǻ�@p             e@������������������������       ������]@�            �g@
                           �?���@�           ��@                           @ϧ��@�            `o@������������������������       �:�fh��@d            `d@������������������������       �Ε>�)3@6             V@                           �?��9Y3@           �{@������������������������       �c�ܻ�@U             `@������������������������       �;|.z�@�            ps@                           @�B�b�?@�           �@                            @�O�8@z           ��@                            �?!մ���@           �|@������������������������       ���+	��@�            `w@������������������������       ���* e@1             U@                           �?OiK�@\            �`@������������������������       �7�*�B�@/             R@������������������������       �<3'
AR@-            �O@                          �3@�ҁ �@*           ��@                           �?/"A�v�
@�           �@������������������������       �����޾	@�            Ps@������������������������       �V�=��,@           �|@                           @�Lc�@�@M           �@������������������������       ��q��Q�@           �z@������������������������       �&n���@=           @@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@      `@      X@     �u@      C@     �~@      (@     �m@      <@     `}@      [@     �P@      @@      V@     �l@      P@     �w@     �q@     �y@      R@     @_@      R@      O@     �a@      ;@     �b@      &@     @_@      5@     �a@     �J@      B@      4@      L@     @T@      A@     �a@     �`@      c@     �B@     �T@      F@      >@      Y@      ,@     �R@      @     �P@      $@      X@      7@      5@      $@      ?@      I@      5@     �S@      H@     @Y@      6@      M@      1@      &@     @P@      @     �K@              <@      $@      M@      "@      2@       @      6@      ;@      .@     �I@      ?@      S@      ,@      1@      @      @      *@      @      :@              1@              3@      @      "@      �?      @      "@      @      1@      (@     �D@      @     �D@      &@       @      J@      @      =@              &@      $@     �C@      @      "@      �?      1@      2@      &@      A@      3@     �A@      $@      9@      ;@      3@     �A@       @      4@      @      C@              C@      ,@      @       @      "@      7@      @      <@      1@      9@       @      1@      (@      "@      &@      @      0@      @      (@              9@      @      �?              @      *@      �?      *@      @      $@      @       @      .@      $@      8@      �?      @      @      :@              *@      "@       @       @      @      $@      @      .@      &@      .@      @      E@      <@      @@      E@      *@      S@      @     �M@      &@     �F@      >@      .@      $@      9@      ?@      *@      P@      U@     �I@      .@      5@      "@      &@      8@      @      ?@      �?      3@      @      $@      *@       @      @       @       @      @      4@      A@      6@      @      ,@       @      @       @      �?      7@      �?      &@      @      @      @       @      @      @      @      @      2@      4@      3@      @      @      �?      @      0@       @       @               @              @      @                       @      @      �?       @      ,@      @              5@      3@      5@      2@      $@     �F@      @      D@       @     �A@      1@      *@      @      1@      7@      @      F@      I@      =@      (@      &@      @      @      "@      @      $@              *@      @      "@      @       @              @      @      @      &@      @      (@      @      $@      .@      ,@      "@      @     �A@      @      ;@      @      :@      *@      &@      @      *@      1@       @     �@@      F@      1@      @     �i@     �L@      A@     `i@      &@     �u@      �?      \@      @     �t@     �K@      ?@      (@      @@     �b@      >@     �m@     �b@      p@     �A@      P@      3@       @      N@      @      R@              E@      @     �S@      7@      @      @      @      H@      ,@      J@      B@     �D@      (@     �J@      @      @      H@      @     �J@              @@      �?      M@      5@      @      @       @      E@      "@      E@      =@      A@      "@     �E@      @      @     �D@       @      E@              ;@      �?      H@      1@      @      @       @     �@@      @      >@      9@      @@      @      $@              @      @       @      &@              @              $@      @                              "@      @      (@      @       @       @      &@      (@       @      (@      @      3@              $@       @      5@       @      �?               @      @      @      $@      @      @      @      @      @              $@              @               @       @      (@      �?      �?                      @      @      @      @      @      @      @      @       @       @      @      .@               @              "@      �?                       @      @       @      @              @             �a@      C@      :@     �a@      @      q@      �?     �Q@      @     @o@      @@      ;@      @      <@      Y@      0@     @g@     @\@      k@      7@     �L@      $@      "@      M@       @     �c@             �D@             �_@      "@      "@              @      K@      @     �P@     �C@     @\@       @      :@      �?      @      7@       @      T@              1@              C@      @      �?              @      7@      �?      8@      "@      J@       @      ?@      "@      @     �A@             �S@              8@             @V@      @       @                      ?@      @      E@      >@     �N@      @     @U@      <@      1@     @U@       @     @\@      �?      =@      @     �^@      7@      2@      @      9@      G@      $@      ^@     �R@      Z@      .@      >@      (@      &@      I@      �?      L@              2@      @     @P@      $@      @       @      *@      3@      "@     �I@      >@      B@       @     �K@      0@      @     �A@      �?     �L@      �?      &@              M@      *@      ,@      @      (@      ;@      �?     @Q@      F@      Q@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�emhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@X���4�@�	           ��@       	                     @}Jm��@�           Ģ@                           @u}�D�@p           ��@                           @�Z�5�6@�           ��@������������������������       �
I�)�@�           Ї@������������������������       ��Y�5��@           �z@                           @7/�"�Z@w           �@������������������������       �Ao�̩	@�             s@������������������������       �q���RM@�            �p@
                           �?�%o�f�@�           ؃@                           @I�ѼJ@�            �r@������������������������       ��le��g@�             m@������������������������       �G�?�.@*             Q@                          �3@�Jެ,@�            �t@������������������������       ����eH�@x            �g@������������������������       �a
����@U             b@                            @���A@�           ��@                           �?᷷�}@�           ��@                          �<@����'@�             r@������������������������       ��p�4]v@�             l@������������������������       �b��z&@$             P@                           �?R�HP �@�           �@������������������������       �����S@�            �s@������������������������       �>����@           �|@                           @'�;@$           P|@                           �? #M@�            �x@������������������������       ��0�sY@�            �t@������������������������       ���|�HG@$            �M@                           �?�K뜍@'             N@������������������������       �ʣS���@             @@������������������������       ���(+3	@             <@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �a@     @V@     @u@     �A@     �}@      &@     `k@      B@      }@      Y@      L@      F@     @Q@      n@      N@     pw@     `r@     �|@     @V@     �d@     @R@     �B@     `k@      .@     pu@      �?      a@      0@     �s@      H@     �@@      4@      6@      b@     �@@     �m@     �d@     �t@      F@      [@      J@      2@      f@      @     Pp@             @V@      *@     `m@      >@      8@      ,@      &@     �Z@      5@     �e@      _@     `q@      @@      Q@     �B@      &@     @b@       @     �c@              N@      $@     �b@      6@      5@      $@      &@      Q@      4@      ]@     �T@      f@      6@     �L@      4@       @     @W@       @      U@             �C@      @     �V@      4@      &@      @       @     �H@      ,@     �R@     �N@     �Y@      0@      &@      1@      @     �J@              R@              5@      @     �N@       @      $@      @      @      3@      @      E@      5@     �R@      @      D@      .@      @      >@      �?     @Z@              =@      @      U@       @      @      @              C@      �?      L@      E@     @Y@      $@      4@      �?      @      ,@      �?      R@              1@              E@      �?      �?       @              :@              <@      4@     �J@      @      4@      ,@      @      0@             �@@              (@      @      E@      @       @       @              (@      �?      <@      6@      H@      @      M@      5@      3@     �E@      (@     �T@      �?      H@      @     �S@      2@      "@      @      &@     �C@      (@     �P@     �E@     �J@      (@      C@      @      @      <@      @      F@              :@              >@      @      @       @      @      0@      @      2@      7@     �B@      @      >@              @      6@      @     �A@              5@              5@       @      �?       @      @      .@      @      0@      1@      @@      @       @      @      @      @              "@              @              "@      @       @                      �?               @      @      @              4@      .@      (@      .@      "@      C@      �?      6@      @     �H@      &@      @      @      @      7@      "@      H@      4@      0@      @      ,@      @       @      (@       @      :@      �?      *@              7@      @      @               @      2@       @      7@      0@      (@      �?      @      $@      @      @      @      (@              "@      @      :@       @      @      @      @      @      �?      9@      @      @      @     �b@     @Q@      J@     @^@      4@     @`@      $@     �T@      4@     �b@      J@      7@      8@     �G@     �W@      ;@      a@     �_@     @`@     �F@      \@      J@     �B@     �Q@      0@     �Y@       @     �G@      @     �\@      A@      .@      $@      :@     @R@      4@     �Z@     �T@     �X@      ;@      1@      &@      .@      3@      @      6@              $@              H@      (@      �?      @      @      ;@      @      =@      ;@      8@      *@      .@      @       @      3@      @      0@              "@              B@      @              @      �?      9@       @      7@      5@      4@      *@       @      @      @                      @              �?              (@       @      �?      �?       @       @      �?      @      @      @             �W@     �D@      6@      J@      *@     @T@       @     �B@      @     �P@      6@      ,@      @      7@      G@      1@     @S@     �K@     �R@      ,@     �@@      &@      (@      2@       @      E@      @      $@      @      ?@       @      �?      @      @      8@      @     �C@      7@      2@      @      O@      >@      $@      A@      @     �C@      �?      ;@              B@      ,@      *@       @      1@      6@      (@      C@      @@      L@      @      C@      1@      .@      I@      @      ;@       @     �A@      ,@     �A@      2@       @      ,@      5@      6@      @      ?@     �F@      @@      2@      ?@      *@      .@      E@      @      :@       @     �A@      ,@      >@      .@       @      ,@      4@      1@      @      :@     �B@      7@      0@      :@      "@      &@      A@      @      7@       @      >@      (@      3@      ,@       @      *@      4@      0@      @      7@      @@      5@      *@      @      @      @       @              @              @       @      &@      �?              �?              �?      �?      @      @       @      @      @      @               @              �?                              @      @                      �?      @       @      @       @      "@       @      @                      �?                                              @                                      @              @       @      @      �?      @      @              @              �?                              �?      @                      �?               @       @               @      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ7b�1hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�D[n��@�	           ��@       	                     @1�a���@�           ~�@                           �?BBT�@�           �@                           �?ᄠ?$\@k           @�@������������������������       �Ų���C@�             y@������������������������       �Ka7��@o           ��@                            �?m�}��@           �{@������������������������       �A�����@r            �f@������������������������       ���@�            �p@
                           �?GQ��{@           ��@                          �?@�-Ex�@�           ȅ@������������������������       �s�-��@�           ��@������������������������       �EN;~�@             �N@                          �9@(�&�@T            �_@������������������������       �� %X��@?            �V@������������������������       �Dī7@             B@                           @(B��@+           (�@                           �?�K��@�           ��@                            �?}��h��@�            @o@������������������������       �{���g�@             H@������������������������       ��,a��@�            @i@                            �?�v�
t,@            |@������������������������       �w��NCO
@M             \@������������������������       ��h�=�R@�             u@                          �2@p��k�@r           p�@                           @ϓ�?	@�            �u@������������������������       �t�X��@@.            �P@������������������������       �ٔk��r	@�            pq@                          �;@g1�s|�@�           ��@������������������������       �|�a�3a@k           @�@������������������������       ���W��
@/             S@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �r@     @_@     @U@     �v@      F@      ~@      @      m@      =@     P|@     �U@      O@     �G@      O@     �m@      R@     �v@     �s@     @}@     @V@     �d@      U@     �I@     �l@     �B@     �l@      @      b@      4@     �k@     �O@     �F@      D@      F@     �a@      H@     �h@     �f@     �l@      O@     �W@      L@      7@     �d@      6@     `a@       @     �T@      "@      c@      ?@      9@      7@      6@     �Z@      A@     �\@     �Z@      e@     �C@      N@     �G@      5@     �\@      3@     �R@       @      M@       @     �Y@      2@      5@      ,@      1@     @Q@      =@     �R@     �Q@     �^@      9@      :@      *@      @      H@      @     �E@              3@       @     �E@       @      @      @      "@      <@      1@      5@      =@     �P@      $@      A@      A@      0@     �P@      .@      @@       @     �C@      @      N@      $@      ,@      $@       @     �D@      (@      K@      E@      L@      .@      A@      "@       @      I@      @      P@              9@      �?      I@      *@      @      "@      @     �B@      @      D@      B@      G@      ,@      $@      @       @      .@      @      8@               @              1@       @      @      @       @      0@              0@      1@      9@      $@      8@      @             �A@              D@              1@      �?     �@@      &@      �?       @      @      5@      @      8@      3@      5@      @     �Q@      <@      <@     �P@      .@     �V@      @     �N@      &@     �P@      @@      4@      1@      6@     �B@      ,@     @T@     �R@     �N@      7@     �M@      2@      8@     �H@      *@     �Q@      @      H@      &@     �L@      >@      2@      0@      4@      A@      @      S@     �P@     �L@      6@     �L@      &@      1@      E@      *@      Q@      @      H@      &@      I@      9@      2@      &@      4@      A@      @     @R@     �L@     �J@      3@       @      @      @      @               @                              @      @              @                              @      "@      @      @      (@      $@      @      1@       @      5@              *@              $@       @       @      �?       @      @      "@      @      "@      @      �?      $@      $@      @      .@              0@              @              @       @              �?              @      @      @      @       @               @              �?       @       @      @              "@              @               @               @               @              @       @      �?      a@     �D@      A@     @`@      @     @o@             @V@      "@      m@      7@      1@      @      2@     �W@      8@     �d@     ``@     �m@      ;@     �G@      (@      &@     �P@      @      [@              A@      @     �Y@      $@      "@      @      "@      <@      6@     �S@     �L@     @T@      ,@      *@      @       @      2@      �?     �G@              &@              ;@      �?       @              @      1@      @      @@      9@     �@@      @      �?               @       @              (@              @              "@                                      �?              @      @      @      @      (@      @              0@      �?     �A@              @              2@      �?       @              @      0@      @      ;@      5@      >@      @      A@      "@      "@     �H@      @     �N@              7@      @      S@      "@      @      @       @      &@      2@      G@      @@      H@      @      @      @      �?      0@              1@              @              8@                      �?       @      @              &@      "@      *@      @      ?@      @       @     �@@      @      F@              4@      @      J@      "@      @       @              @      2@     �A@      7@     �A@      @     @V@      =@      7@     �O@      @     �a@             �K@      @     @`@      *@       @      @      "@     �P@       @     �U@     �R@     �c@      *@      .@      @      @      .@      �?      Q@              ?@              M@      @                              3@              >@      6@     �R@      �?      @                      @              0@                              @                                      @              @      �?      8@              $@      @      @      &@      �?      J@              ?@              J@      @                              .@              7@      5@      I@      �?     �R@      8@      3@      H@       @     �R@              8@      @      R@      $@       @      @      "@     �G@       @     �L@      J@      U@      (@     �Q@      1@      (@      G@       @     �Q@              8@      @     �P@      @      @      @      @      F@       @      E@     �G@      Q@      (@      @      @      @       @              @                              @      @       @               @      @              .@      @      0@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJC��jhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@K���@�	           ��@       	                    �?ʡ�l�@�           ��@                           �?��H��@           ��@                           @���?@�            �u@������������������������       �X�>{@�            �s@������������������������       ��o�X�@             ?@                           �?�^��@4           �}@������������������������       �g)C�<�@l            �e@������������������������       ���ۓ�4@�            �r@
                            �?6�7�@�           @�@                           @��\+f^@J           ��@������������������������       �؄�8��@�           P�@������������������������       �{���6w@�            �j@                            @Y��o8�@�           ��@������������������������       ���#.@�            �u@������������������������       � 5�5�M@�            �q@                           @1	a��@�           �@                          @A@��ԉK@           x�@                            �?̀_q=@�           ؒ@������������������������       �l����@�            �w@������������������������       ����@           �@                           @{�D4>
@             D@������������������������       �
=��,@             4@������������������������       ��?o��:@             4@                          �9@�ryA^@�            Pr@                            �?a��0�R@o            �e@������������������������       ��:n��	@             E@������������������������       ������B@S            ``@                           @t����@K             ^@������������������������       �e��l�@7             U@������������������������       ��L�a`�@             B@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �r@      b@     �S@     �v@      K@     �|@      @     `m@      @@     �{@     �X@     �K@      E@     �M@     �p@      M@      w@     Pu@     �{@      S@     `c@     �N@      D@     @n@      3@     u@      @     �`@      .@     Pr@     �G@      A@      0@      4@     @b@      >@      m@      i@      s@     �D@      H@      :@      3@     @U@      .@     �R@      @      J@      "@     @V@      3@      (@      @      ,@     �I@      0@      T@     @V@     @Y@      *@      7@       @       @      C@      �?      D@              ,@      @      @@       @      @              @      5@      ,@      5@      A@      Q@      @      6@       @       @      :@      �?      D@              *@      @      >@       @      @              @      3@      (@      4@      ?@     �N@      @      �?                      (@                              �?               @                                       @       @      �?      @      @              9@      2@      &@     �G@      ,@     �A@      @      C@      @     �L@      &@       @      @      $@      >@       @     �M@     �K@     �@@      @      &@      @              4@      @      4@              .@              2@      @      �?      @       @      @      �?      =@      2@      "@       @      ,@      &@      &@      ;@      $@      .@      @      7@      @     �C@      @      @      �?       @      7@      �?      >@     �B@      8@      @     �Z@     �A@      5@     �c@      @     `p@             �T@      @     �i@      <@      6@      &@      @     �W@      ,@      c@      \@     �i@      <@      N@      6@      &@     �V@       @     @c@              G@       @     �`@      3@      @      &@       @      E@      &@      W@     �P@     �`@      7@     �H@      $@      $@     �R@       @     �]@             �C@      �?      ]@      *@      @       @              @@      "@     �O@      B@      \@      0@      &@      (@      �?      0@              B@              @      �?      1@      @              @       @      $@       @      =@      >@      7@      @     �G@      *@      $@     �P@       @      [@             �B@      @     �Q@      "@      0@              @     �J@      @      N@      G@     �Q@      @      0@       @      @     �B@             �L@              6@      @      E@      @      *@              @      ;@              C@      8@      G@      @      ?@      &@      @      >@       @     �I@              .@              =@      @      @              �?      :@      @      6@      6@      8@       @     �a@      U@      C@     �]@     �A@      ^@      @      Y@      1@     `b@      J@      5@      :@     �C@      _@      <@      a@     �a@     �`@     �A@      Y@     �Q@      B@     �Y@      @@     @V@      @     @W@      1@     @^@     �F@      2@      4@      =@     �X@      :@     @Z@      \@      X@     �@@     �X@     �N@      A@     @X@      @@     @V@      @     �V@      1@      ^@     �C@      ,@      4@      =@     �W@      :@     �Y@     �[@     �W@     �@@      >@      :@      @      7@      .@      >@      �?      6@      �?      ;@      $@              @      .@      E@      "@      8@     �H@      A@      $@     @Q@     �A@      ?@     �R@      1@     �M@       @      Q@      0@     @W@      =@      ,@      ,@      ,@     �J@      1@     �S@     �N@     �N@      7@      �?      "@       @      @                              @              �?      @      @                      @               @       @      �?                       @       @      �?                               @                      �?      �?                      @                              �?              �?      �?              @                              �?              �?      @      @                                       @       @                     �D@      ,@       @      1@      @      ?@              @              :@      @      @      @      $@      9@       @      ?@      <@      C@       @      3@       @      �?      (@              2@              @              5@      @                       @      ,@      �?      7@      1@      3@      �?       @      @      �?      @              @                              @      �?                       @      @      �?       @              �?              &@       @              "@              &@              @              0@      @                      @      "@              5@      1@      2@      �?      6@      @      �?      @      @      *@              �?              @       @      @      @       @      &@      �?       @      &@      3@      �?      &@      @      �?       @      @      *@                               @       @      @      @       @       @              @      @      *@      �?      &@                      @                              �?              @                                      @      �?      @      @      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ
1hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?O*���@�	           ��@       	                   �:@ ��v�@�           h�@                           �?�\U�3@;           �@                          �4@E�b���@1           �}@������������������������       �ˌ`���@�            �k@������������������������       �"�'+�@�            �o@                            �?T� �g�@
           ��@������������������������       ��n�l�@|            �h@������������������������       ��\�@�           Ђ@
                          �<@E��s�3@n             d@                          �;@8av�z@8            @W@������������������������       �	�@!            �M@������������������������       ��
û�2@             A@                            @�6sc�@6            �P@������������������������       �s����@&            �G@������������������������       �l�u5x
@             4@                           @.�}�@           ^�@                           �?4�T�>�@v           ��@                           @Ǥ��*@�            �w@������������������������       �&Ox�(t
@            �I@������������������������       ���S�q�@�            �t@                           �?������@�           Ԑ@������������������������       ��1 �@�            �@������������������������       ��?��t@�            w@                           @N]Q��u@�           ��@                           @����@V           `�@������������������������       �R��N��@%           �{@������������������������       �"��f�@1            @S@                           @��e�@<           0@������������������������       �k+�ٹ@�            �s@������������������������       ���@�%@s            �f@�t�b��     h�h5h8K ��h:��R�(KKKK��h��B`       Pu@     �`@     �V@      w@      ?@     p~@      @     �k@      @@     0{@     �Z@      H@     �A@      R@     �n@     �S@     �v@     �t@     0y@     �T@     �\@      B@     �@@      \@      @     �l@       @     �T@      @     @d@     �A@      5@       @      ;@     @X@      2@     `a@     �[@     �c@      C@      [@      ;@      9@      Y@      @     @k@      �?     @R@      @     �b@      @@      1@       @      8@     @T@      @      `@     @W@     �b@      A@     �E@      ,@      .@      <@      @      O@      �?      >@       @     �H@      .@      &@      �?      1@      <@      @     �J@      ;@      J@      2@      7@      $@      @      .@      @      ?@              $@              =@      @      @      �?       @      5@       @      .@      ,@      <@      @      4@      @      "@      *@      �?      ?@      �?      4@       @      4@      (@      @              .@      @      @      C@      *@      8@      ,@     @P@      *@      $@      R@             �c@             �E@      �?      Y@      1@      @      �?      @     �J@       @     �R@     �P@      X@      0@      &@      �?      @      6@             �@@              &@      �?      :@      @      �?      �?              3@       @      0@      1@      7@      @      K@      (@      @      I@             �^@              @@             �R@      *@      @              @      A@             �M@     �H@     @R@      $@      @      "@       @      (@      �?      (@      �?      $@      @      *@      @      @      @      @      0@      &@      &@      1@      "@      @      @      @      �?      &@              @      �?      @      @      @      �?      @      @              "@      @       @      ,@       @      �?      �?                      @              @      �?      @      @      @      �?      @       @              @      @       @      (@      @      �?       @      @      �?      @                              �?               @              �?      �?               @       @      @       @      @              @      @      @      �?      �?       @              @               @       @              @      @      @      @      @      @      �?      @      @      @      @                       @              �?               @       @              @       @      @       @       @      �?      �?                      �?      @      �?      �?                       @                                              �?      @       @      �?       @              @     @l@     �X@      M@      p@      :@     p@      @     @a@      :@     q@     �Q@      ;@      ;@     �F@     �b@      N@      l@     �k@     �n@      F@     �`@     �P@     �G@      d@      4@     �]@       @      X@      4@      a@     �J@      0@      4@     �@@     @W@     �C@     �_@     @`@     @]@      <@      B@      6@      ,@      C@      @      @@      �?      1@              ?@      @      @       @      @      7@      ,@      E@     �@@      J@      @      @       @              @              *@              �?              @      @                              �?      @      @      @      @      �?     �@@      4@      ,@     �A@      @      3@      �?      0@              <@      @      @       @      @      6@      @     �B@      ;@     �H@      @     �X@     �F@     �@@     �^@      1@     �U@      �?     �S@      4@     �Z@      G@      *@      2@      =@     �Q@      9@      U@     @X@     @P@      7@      P@      :@      8@     @V@      ,@      J@      �?     �L@      3@      K@      A@      "@      &@      8@      B@      3@      F@     �P@     �H@      0@      A@      3@      "@     �@@      @      A@              6@      �?      J@      (@      @      @      @      A@      @      D@      ?@      0@      @      W@      @@      &@      X@      @     `a@       @      E@      @      a@      2@      &@      @      (@      L@      5@     �X@     @W@      `@      0@      C@      ,@      @     �O@      @     @S@              2@      @     �R@      &@      @      @      @      0@      *@      L@      C@     �R@      @     �A@      ,@      @     �M@      @     �I@              .@      @     �Q@      &@      @      @      @      *@      *@     �G@      B@     �K@      @      @                      @              :@              @      @      @                                      @              "@       @      4@              K@      2@       @     �@@      @      O@       @      8@             �N@      @      @      @      @      D@       @      E@     �K@      K@      &@      B@      &@      @      1@      @      C@       @      2@             �B@      @      @      @      @      >@              7@      9@      F@      @      2@      @      �?      0@              8@              @              8@      �?      �?      �?      �?      $@       @      3@      >@      $@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJM<�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?6�.�~@�	           ��@       	                     @�#�!ٿ@�           ��@                           �?w�}!~@W           �@                          �5@2�2���@�            t@������������������������       �,Dw��t@q             f@������������������������       ��x�	�@[             b@                           �?F<�)��@�           �@������������������������       �Ef)��`@�            �o@������������������������       �w鋾�@�             x@
                           �?��Z㆜@�            �@                          �5@�[�[��@�             k@������������������������       ��Ow��Y@N            �_@������������������������       ��K:W�_@>            �V@                           �?�A�ÿ@           �|@������������������������       ��t�'�@;             Z@������������������������       �8k*L[�@�            0v@                           @�^�PxB@�           ơ@                           @�u	���@B           ��@                           �?�	�sK$@           0�@������������������������       �L6���@�            �w@������������������������       ������@           �z@                            @/8���O@@           �@������������������������       ��I�ѿW@�            @y@������������������������       ��PREa�@C            �Y@                           @��67@T           �@                            �?L`��@M            �Z@������������������������       �S��=��@"            �F@������������������������       ��s��@+            �N@                           @�B&V�@           Ȋ@������������������������       �k�QH��@`           �@������������������������       �KӢ3�@�            `q@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@      [@      W@     �w@     �H@     @@       @     @h@      @@     P}@     �Y@     �L@      =@     �P@     @j@      R@     �u@     Pt@     �{@     @S@     �a@     �K@      N@     �b@      >@     �b@       @     �Y@      5@     �f@     �I@      A@      0@      D@     @U@      E@     �a@      a@     @d@      ?@     �P@      C@     �A@     �\@      4@     @W@      @      K@      &@     @^@      <@      0@      "@      3@      F@      <@     �P@     �R@     �X@      5@      .@      "@      (@      >@       @      G@              .@      �?      K@      0@      "@      @      @      (@      @      :@      9@      @@      @      .@      @      @      7@              3@              "@      �?      =@       @      @              @      @              .@      (@      7@      �?              @      @      @       @      ;@              @              9@      ,@      @      @      �?      @      @      &@      *@      "@      @     �I@      =@      7@     @U@      2@     �G@      @     �C@      $@     �P@      (@      @      @      ,@      @@      9@     �D@     �H@     �P@      0@      2@      *@      &@     �@@              7@      �?      (@       @      6@      @       @              @      (@      $@      0@      5@     �C@      @     �@@      0@      (@      J@      2@      8@      @      ;@       @     �F@      @      @      @       @      4@      .@      9@      <@      ;@      "@      S@      1@      9@     �A@      $@     �K@      @     �H@      $@      N@      7@      2@      @      5@     �D@      ,@      S@      O@      P@      $@     �C@      @      "@      3@       @      "@              (@       @      9@       @       @      @      @      "@      @      2@      7@      3@              ?@      �?      @      $@              @              @              (@      @      �?      @      �?       @              (@      ,@      &@               @      @      @      "@       @       @              @       @      *@       @      �?              @      �?      @      @      "@       @             �B@      (@      0@      0@       @      G@      @     �B@       @     �A@      .@      0@      @      ,@      @@       @      M@     �C@     �F@      $@      @      @       @      @      �?      0@      �?      @      @       @      @       @                      @       @      3@       @      (@      @      >@       @      ,@      &@      @      >@       @     �@@      @      ;@      &@      ,@      @      ,@      =@      @     �C@      ?@     �@@      @     �i@     �J@      @@      m@      3@      v@             �V@      &@      r@      J@      7@      *@      ;@     @_@      >@      j@     �g@     pq@      G@     �\@      B@      3@     �a@      $@      j@             �O@      $@     �b@      A@      0@      $@      ,@      Q@      :@     �^@     @W@     �a@     �@@     @Q@      3@      @     @S@      @     �b@              E@      @     �W@      1@      "@      @      @     �F@      &@     @U@      J@     �S@      ;@     �@@      &@       @      ?@      @      K@              =@      @     �F@      @      @      @      @      3@      @      A@      ;@      G@      ,@      B@       @      @      G@      @     @X@              *@              I@      $@      @      �?      @      :@      @     �I@      9@      @@      *@      G@      1@      *@     @P@      @      M@              5@      @      L@      1@      @      @       @      7@      .@      C@     �D@      O@      @     �@@      (@      $@      N@      @      F@              *@      @      E@      .@      @      @       @      5@      $@      8@      B@     �I@      @      *@      @      @      @              ,@               @              ,@       @              �?               @      @      ,@      @      &@             @V@      1@      *@     �V@      "@     �a@              <@      �?      a@      2@      @      @      *@     �L@      @     @U@      X@     `a@      *@      @                      "@              ?@              �?              @                                      @              @      @      ?@      �?      @                      @               @              �?              @                                                      @       @      &@      �?       @                      @              7@                              �?                                      @              �?      @      4@             �T@      1@      *@     �T@      "@      \@              ;@      �?     @`@      2@      @      @      *@     �I@      @     �S@     @V@      [@      (@      P@      $@       @     �H@      @     �T@              9@      �?      X@      &@      �?       @      @      =@       @     �F@      I@     �U@      $@      2@      @      @     �@@      @      >@               @              A@      @      @      �?      "@      6@       @      A@     �C@      6@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��"ghG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �6@s�|==r@�	           ��@       	                     @�]h|@�            �@                          �5@�R~�@k           �@                            �?��̫�@�           �@������������������������       �\��7^@�           �@������������������������       ������
@�            �w@                           @:�
�@|            �g@������������������������       �E|�w�@S             `@������������������������       ���<o�	@)             O@
                          �5@���~�@�           x�@                           �?"����@[           ��@������������������������       ���3�_�@�            �o@������������������������       ��1F׀@�            0s@                           �?2;<��@9            �W@������������������������       �#_�dyY@             I@������������������������       ����=e|@            �F@                           �?��g�r@�           �@                           @�	���@�           (�@                           �?�����@�           ��@������������������������       ���*a�@�            �i@������������������������       �4�e���@a           �@������������������������       ���Dh�@             4@                            @R��&l@�           ��@                          �7@Mf�l��@m           ��@������������������������       �
}k�7�	@H            �X@������������������������       ��|D�� @%           `}@                          �8@��B��@M             _@������������������������       �4~U�̸@             F@������������������������       �b�K��@2             T@�t�bh�h5h8K ��h:��R�(KKKK��h��B        v@      `@     �U@     �t@      C@     P@      @     �m@      ;@     �|@     @U@     �P@      @@      O@      m@      Q@     `x@      s@     �z@     �R@     �g@      N@     �H@     �j@      ,@     px@       @      a@      3@     �r@     �E@      H@      ,@      :@     �a@      7@     Pp@      h@     �q@      D@     @]@      I@      6@     @e@      @     pr@      �?     @X@      0@      k@      3@     �B@      ,@      2@     �Y@      .@      h@     �a@     @m@      =@     �Z@     �H@      .@     �c@       @      o@              U@      $@     �h@      .@      A@      *@      ,@      W@      ,@     �e@     @a@     �j@      8@      T@     �F@      ,@     @`@       @     `d@              M@      $@     �b@      (@      :@      *@      @     �Q@      ,@     �`@     �]@      d@      4@      ;@      @      �?      =@             @U@              :@              H@      @       @              "@      6@              D@      4@      K@      @      $@      �?      @      &@      @     �G@      �?      *@      @      4@      @      @      �?      @      &@      �?      3@       @      4@      @       @              @      @      @      <@      �?      @      @      ,@      @      @      �?      @      &@      �?      ,@      �?      0@      �?       @      �?      @       @              3@              @      @      @                                                      @      �?      @      @     �R@      $@      ;@     �E@       @      X@      �?     �C@      @     �T@      8@      &@               @      C@       @      Q@     �J@     �I@      &@     @Q@      @      8@     �D@      @     �S@      �?      A@      @     �P@      3@      @              @      >@      @     �J@     �G@      I@      &@     �D@      �?      @      9@      @     �C@              "@              A@       @      �?              �?      $@       @      6@      0@      ;@       @      <@      @      2@      0@      @     �C@      �?      9@      @     �@@      &@      @              @      4@      @      ?@      ?@      7@      @      @      @      @       @      �?      2@              @              .@      @      @               @       @      �?      .@      @      �?              @               @       @      �?      "@              �?               @      �?      @                      @      �?      @      @      �?              �?      @      �?                      "@              @              @      @                       @       @              $@      �?                     @d@      Q@     �B@     @]@      8@     �[@      @     �Y@       @     `d@      E@      2@      2@      B@     �V@     �F@      `@     @\@     �a@      A@     �P@      D@      8@     �N@      .@      H@      @     �N@      @     @T@      3@      .@      .@      5@     �I@      3@      Q@     �N@     @S@      4@     �P@      A@      8@     �N@      *@      H@      @     �N@      @      T@      1@      .@      .@      5@     �G@      3@     @P@      N@      S@      4@      0@       @      @      3@              7@       @      .@      @      7@      @      @      @       @      2@       @      5@       @      4@       @     �I@      :@      1@      E@      *@      9@       @      G@      @     �L@      (@      (@      &@      3@      =@      1@      F@      J@      L@      (@              @                       @                                      �?       @                              @              @      �?      �?             �W@      <@      *@      L@      "@      O@              E@       @     �T@      7@      @      @      .@      D@      :@     �N@      J@     �P@      ,@     @T@      2@      $@      G@      @      K@              @@       @     �P@      1@               @      *@      C@      8@     �I@     �E@      N@       @      ;@       @      @      .@              @                              &@      �?                      �?      @      @      *@      @       @       @      K@      0@      @      ?@      @      H@              @@       @     �K@      0@               @      (@     �@@      5@      C@      B@      M@      @      ,@      $@      @      $@      @       @              $@              0@      @      @      �?       @       @       @      $@      "@      @      @      @      @       @      @              �?              �?              *@      @                              �?                      @      �?       @      &@      @      �?      @      @      @              "@              @      @      @      �?       @      �?       @      $@      @      @      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�*�ChG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?Ed��%�@�	           ��@       	                    �?X��@�           x�@                           �?!z���k@[           ��@                           @;�̦��@�            �k@������������������������       �F:�Bb�@R            �`@������������������������       ��4cV�@7            @U@                            �?h�[�w�@�            �u@������������������������       �0���?�@�            @l@������������������������       �!6i,��@O            @^@
                          �:@%%9�{@�           ��@                            @s~���@           ��@������������������������       ���i 0@           �y@������������������������       � ���Y[@�            �y@                          @@@� +�@�             n@������������������������       �\�}�c@{             i@������������������������       ���j�~r
@            �C@                            @���&Q@�           ֡@                          �6@�����@�           ��@                           @j�=�3@           `�@������������������������       �DJ���H@N           H�@������������������������       �|[d�W�@�           x�@                          �7@�?�r�@i           ��@������������������������       �
5h�*+
@F            �^@������������������������       ��=3���@#           `}@                           @+�Ї@           0|@                           @�8�1^@�            @l@������������������������       �sj-��@-             U@������������������������       ��FM^I@]            �a@                           @� ٝZ@�             l@������������������������       ��d�И	@*            @P@������������������������       ���ůA'@f             d@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �v@      `@     �W@     @t@     �B@     �~@      @      k@      <@     �{@     @Z@      K@      :@      T@     p@     �N@     0w@     �q@     `|@      W@     @c@     �Q@     @P@     @^@      >@      b@      @     �[@      5@      b@     �L@      =@      ,@     �F@     �V@      A@      a@     �_@     `h@     �B@      N@      .@      >@      F@       @     �P@       @      :@      @     �J@      3@      @       @      @      C@      .@      D@     �D@      U@      *@      5@       @      ,@      2@      �?      <@      �?      "@      @      7@      @                      @      *@      @      &@      3@     �E@      @      $@      �?      @      .@              5@      �?       @      @      1@      @                      @      @       @      @      @      <@              &@      �?       @      @      �?      @              �?              @                              �?      @       @       @      (@      .@      @     �C@      *@      0@      :@      �?      C@      �?      1@       @      >@      0@      @       @      @      9@      &@      =@      6@     �D@      $@      6@       @      $@      8@              6@              "@      �?      2@      ,@      @       @      @      3@      &@      $@      (@      =@       @      1@      @      @       @      �?      0@      �?       @      �?      (@       @      �?                      @              3@      $@      (@       @     �W@      L@     �A@     @S@      <@     �S@      �?      U@      0@      W@      C@      8@      (@      C@     �J@      3@      X@     �U@     �[@      8@     �S@      C@      2@      J@      5@     @S@      �?     �I@      ,@     @U@      =@      4@       @      >@      D@      "@      V@     �N@     �T@      4@      @@      ;@      @     �@@      $@      ?@      �?      8@      "@      I@      @      *@      �?      $@      <@      @      D@      :@      J@      "@      G@      &@      &@      3@      &@      G@              ;@      @     �A@      8@      @      @      4@      (@      @      H@     �A@      ?@      &@      0@      2@      1@      9@      @       @             �@@       @      @      "@      @      @       @      *@      $@       @      9@      <@      @      0@      &@       @      3@      @      �?              @@       @      @      @      @      @      @      *@      "@      @      8@      ;@      @              @      "@      @      �?      �?              �?               @      @              �?       @              �?      @      �?      �?             @j@      M@      >@     `i@      @     �u@       @     �Z@      @     pr@      H@      9@      (@     �A@     �d@      ;@     `m@     �c@     0p@     �K@     �c@     �F@      8@     @e@      @     �q@       @     @R@      @     �n@      B@      2@      $@      =@     �`@      1@     �h@     �`@     �j@     �@@     �R@      7@      3@     �^@       @     @k@             �J@       @     �g@      3@      .@      @      &@      U@      &@      a@     �T@     �b@      5@      <@      @      $@     �L@             �R@              2@              V@      @      @      �?      &@     �C@      $@     �P@      A@     �J@      &@      G@      1@      "@     @P@       @     �a@             �A@       @     �Y@      (@      "@      @             �F@      �?     �Q@     �H@     �W@      $@     �T@      6@      @      H@      @     @Q@       @      4@      @     �K@      1@      @      @      2@      H@      @     �M@      I@     �P@      (@      >@      @       @      ,@              *@                      �?      @      �?                       @      &@      �?      ,@      1@      @      @      J@      0@      @      A@      @      L@       @      4@      @     �I@      0@      @      @      0@     �B@      @     �F@     �@@     �O@      "@      K@      *@      @     �@@       @      M@              A@      �?     �H@      (@      @       @      @      A@      $@     �C@      8@     �F@      6@      9@      @       @      .@       @      ;@              7@              4@      $@      @               @      1@              1@      $@      9@      5@      &@      �?       @      @      �?       @              "@              @      @      @                      @              @      @      @      *@      ,@      @              (@      �?      3@              ,@              *@      @                       @      ,@              $@      @      4@       @      =@      @      @      2@              ?@              &@      �?      =@       @      @       @      @      1@      $@      6@      ,@      4@      �?      $@      @                              3@              @      �?       @                      �?      @      @      @      @       @      @              3@              @      2@              (@               @              ;@       @      @      �?      �?      &@      @      3@      (@      1@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ+l�.hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��@�	           ��@       	                    �?�Gũ�@           ̙@                           �?�s���@d           ��@                           @�����@�            �m@������������������������       ��X/���@             k@������������������������       ��(9�"@             6@                            @�'�>�z@�            �t@������������������������       ��.��@�            `n@������������������������       ����"o@:            �V@
                          �:@}8���@�           ܐ@                           �?�Y��@�           (�@������������������������       �)����L@�            �p@������������������������       ��{�I��@R           ��@                          �@@~$O�ra@�             q@������������������������       ��J&�0@�             n@������������������������       �)��
�e	@             A@                            �?Ѷ�� �@�           ��@                           @�D1���@|           ��@                           �?@:=�@�            Pp@������������������������       �7���`�
@w            �g@������������������������       �Ӭ~�q,
@)            @R@                           �?bdL~�@�            �v@������������������������       �,1�M&�@l            �e@������������������������       �P�'�I@p            �g@                           @��d"l�@           ��@                           @|��2�@�           �@������������������������       �4fnT@�            �w@������������������������       ��X�R8�@�           0�@                           @kk�T�@|           �@������������������������       �|p�RDb@�            `m@������������������������       �.0 �6@�            pw@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       t@     ``@     @V@     `u@      A@     �|@       @     `n@     �@@     �}@     �V@      L@     �B@      S@     �i@     @Q@     x@     pr@     @~@     �S@     �_@      S@      L@      b@      2@     @a@       @     �^@      5@     �c@      G@      =@      1@     �I@     @R@      ?@     �e@     �_@      i@      A@     �E@      5@      8@     @P@      @     �I@              >@      @     �K@      ,@      @       @      *@      9@      &@     �I@      F@     @V@      ,@      2@      @      0@      4@       @      3@              &@              :@      @      �?      @      $@      "@      @      (@      7@      G@      @      (@      @      &@      2@       @      3@              &@              5@      @      �?      @      $@      "@      @      (@      4@     �F@      @      @              @       @                                              @                                                              @      �?              9@      ,@       @     �F@      @      @@              3@      @      =@      $@      @      @      @      0@      @     �C@      5@     �E@       @      6@      *@       @     �A@              :@              (@              4@      @       @      @      @      "@      @      :@      *@     �@@      @      @      �?              $@      @      @              @      @      "@      @       @                      @              *@       @      $@      @     �T@     �K@      @@      T@      (@     �U@       @      W@      2@      Z@      @@      8@      "@      C@      H@      4@     �^@     �T@     �[@      4@     �Q@      >@      1@      J@      &@      U@      @      K@      .@     @W@      5@      ,@      @      =@      C@      @     @Z@     �I@     �V@      0@      B@      @      @      *@      @      A@              1@              @@      @       @      �?      @      &@      @      H@      .@      @@      @      A@      7@      ,@     �C@       @      I@      @     �B@      .@     �N@      .@      (@      @      :@      ;@       @     �L@      B@      M@      (@      *@      9@      .@      <@      �?      @      @      C@      @      &@      &@      $@      @      "@      $@      .@      2@      @@      5@      @      *@      2@      $@      9@      �?      @      @      A@      @      &@       @      @      �?      @      $@      (@      2@      @@      4@      @              @      @      @                              @                      @      @      @       @              @                      �?             `h@     �K@     �@@     �h@      0@     �s@             @^@      (@     �s@      F@      ;@      4@      9@     �`@      C@     `j@      e@     �q@     �F@      Q@      3@      .@      P@       @     �U@              6@      �?      V@      (@       @       @       @      C@      "@     �Q@      :@     @S@      $@      9@              @      5@       @     �G@              *@      �?     �D@      @       @      @              .@      @      9@      "@      C@       @      3@              @      .@       @      @@              &@      �?     �@@      @                              $@      �?      1@      "@      =@       @      @                      @              .@               @               @               @      @              @      @       @              "@             �E@      3@      (@     �E@              D@              "@             �G@       @              �?       @      7@      @     �F@      1@     �C@       @      1@      &@      �?      5@              9@               @              :@       @                      @      (@       @      7@      ,@      "@      @      :@       @      &@      6@              .@              @              5@      @              �?      @      &@      �?      6@      @      >@       @     �_@      B@      2@     �`@      ,@      m@             �X@      &@     �l@      @@      9@      (@      1@     �W@      =@     �a@     �a@     �i@     �A@      S@      7@      .@      X@      &@      c@             �I@      $@     �a@      2@      1@      @      @      J@      =@      U@     �S@     `a@      7@      B@      0@      @     �D@      @      F@              6@              F@      &@      @      @              :@      &@      =@     �B@      >@      .@      D@      @       @     �K@      @     @[@              =@      $@     @X@      @      ,@      @      @      :@      2@     �K@      E@     @[@       @     �I@      *@      @     �B@      @     �S@              H@      �?     �V@      ,@       @      @      ,@     �E@             �L@     �O@      Q@      (@      4@       @      �?      *@      �?     �D@              <@              >@       @      @       @              0@              ,@      @@      7@      @      ?@      &@       @      8@       @      C@              4@      �?      N@      (@      @      @      ,@      ;@             �E@      ?@     �F@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�IhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@��L5�@�	           ��@       	                    @��=N�@�           ¢@                           �?�l҆�@@�           p�@                          �5@:G�_�@�           ��@������������������������       �8It�K�@P           Ȁ@������������������������       �t��fO�@>            �W@                          �1@�����%@�           ��@������������������������       ��1�_N�	@�            Pt@������������������������       �$�~@$           ��@
                          �3@�� o�@j           (�@                          �2@��fk�>@�            0r@������������������������       �5��S	@�            @k@������������������������       ��F=�� 	@,            @R@                           �?wƄ d@�             r@������������������������       ���T�@A            @Z@������������������������       �X�t)@q             g@                           �?���A�@�           ��@                          @A@��.�8@�           (�@                          �:@��b�L@�           (�@������������������������       �ԙxM��@)           `}@������������������������       ��YAj�@�            �r@                           �?p)	{@             @@������������������������       �+�%W�@             0@������������������������       �>��_�@
             0@                           @F�n�@�           �@                           @�5ؗ)@	           �z@������������������������       �Y28`.�@�            �t@������������������������       ����Q�G@B             X@                           @����@�            �q@������������������������       �I���"@4             T@������������������������       ��UU��\@�             i@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@      b@      U@     Pv@      A@     �~@       @     @o@      <@     �|@     @^@      M@      B@     �N@     �n@     �M@     Pv@     �r@     �y@     �V@     �g@     �R@      E@      m@      *@     �v@      �?     �a@      (@      r@      N@     �E@      *@      5@      b@      7@      k@      f@     �r@      H@     @a@      C@      <@     �f@      (@     pq@      �?     �\@      @     �n@      E@      ?@      $@      0@     @[@      2@     �c@      \@      n@     �E@      L@      4@      $@     @R@      "@     @R@      �?      E@      @     �N@      7@      ,@       @      ,@      B@      @      M@      B@     �R@      2@     �K@      (@       @     @Q@      @      K@      �?      @@      @     �G@      2@      *@       @      $@      B@      @      H@      @@     @P@      1@      �?       @       @      @       @      3@              $@              ,@      @      �?              @                      $@      @      $@      �?     �T@      2@      2@     �[@      @     �i@              R@      �?     �f@      3@      1@       @       @     @R@      &@     �X@      S@     �d@      9@      $@       @       @      2@       @     �R@              3@              N@      @              �?      �?      (@      @     �A@      ,@      J@      ,@      R@      0@      0@      W@      �?     ``@             �J@      �?     �^@      .@      1@      @      �?     �N@      @     �O@      O@     �\@      &@      J@     �B@      ,@      I@      �?      U@              :@      @      G@      2@      (@      @      @     �A@      @     �N@      P@      L@      @      =@      (@      (@      A@              I@              "@              3@      "@      �?              �?      4@      @      <@      7@      C@       @      ;@      &@      "@      @@             �B@              @              0@      @      �?              �?      *@      @      $@      3@      :@       @       @      �?      @       @              *@              @              @      @                              @              2@      @      (@              7@      9@       @      0@      �?      A@              1@      @      ;@      "@      &@      @      @      .@      �?     �@@     �D@      2@      @      ,@      @      �?      $@              2@               @      �?      @       @      @                      @              "@      3@      @              "@      4@      �?      @      �?      0@              .@      @      4@      �?       @      @      @      (@      �?      8@      6@      *@      @     @a@     @Q@      E@      _@      5@     �_@      @     �[@      0@      e@     �N@      .@      7@      D@      Y@      B@     �a@      ^@      \@     �E@      M@      F@     �@@      P@      (@      K@      @     �R@      $@      Q@      @@      $@      0@      8@     �L@      7@     @R@     @P@      N@      6@     �L@     �A@      =@      O@      (@      K@      @     �R@      $@     �P@      ;@      "@      $@      8@      L@      7@     @R@      P@      N@      6@      A@      2@      2@     �B@      @     �D@       @      D@      "@     �A@      *@      @      @      2@      D@      @     �K@     �C@      ?@      1@      7@      1@      &@      9@      @      *@      @      A@      �?      ?@      ,@       @      @      @      0@      3@      2@      9@      =@      @      �?      "@      @       @                                               @      @      �?      @              �?                      �?                              @      @       @                                                       @               @              �?                      �?                      �?      @      �?                                                       @      @      �?      @                                                              T@      9@      "@      N@      "@     @R@      �?      B@      @      Y@      =@      @      @      0@     �E@      *@     �P@     �K@      J@      5@     �L@      .@      @      A@      @     �K@              6@      @     @R@      ,@       @      @      �?      7@       @      C@      =@      >@      0@      E@       @       @      >@      @      J@              5@      @     �K@      $@       @       @              3@       @      8@      6@      2@      .@      .@      @      @      @              @              �?              2@      @               @      �?      @              ,@      @      (@      �?      7@      $@      @      :@      @      2@      �?      ,@      @      ;@      .@      @      @      .@      4@      &@      =@      :@      6@      @       @      �?      @      @      �?      (@      �?       @      @      $@      @       @       @      "@      �?       @      "@      @      @       @      5@      "@      �?      5@      @      @              (@              1@      (@      �?      �?      @      3@      "@      4@      5@      1@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�
�[hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?������@�	           ��@       	                    �?��-s��@           ��@                           �?l����E@}           �@                           �?&����@�             j@������������������������       ��G����@o            �e@������������������������       �����.e@             B@                           �?��%eK�@�            0y@������������������������       ��d�t^�@�             v@������������������������       ����V��@$            �I@
                           �?W~x�@�           �@                           @}h��P�@�             u@������������������������       �����@�            �j@������������������������       �
�9��[@S             _@                           @/2���>@�           ��@������������������������       ���m @x           8�@������������������������       ��Mß@A            �[@                           @�42D��@�           ¡@                           @50*�@�           |�@                           @�3㶌@�           �@������������������������       ��|j�'@{            �@������������������������       �d�ئ�4@@           �@                           @����@�            �u@������������������������       ����)-�@7            �U@������������������������       ���Y@�            �p@                          �6@��0.�?@            �@                           @��4�U@J           ��@������������������������       �N�El<*@<           0@������������������������       ����T�@             =@                          �<@�QB���@�             s@������������������������       �/�K��@�             o@������������������������       �3fR3v@%            �L@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       @t@      a@     �U@     @u@      D@     �z@      @     �m@     �A@     0z@     @Z@      Q@      >@      U@     �p@     �O@     py@      s@      |@     �S@     @^@     �R@      J@      a@      9@     �`@      @     @]@      8@     �`@      I@      B@      0@     �J@     �[@     �A@     �b@     @b@     �f@     �C@      D@      2@      6@      K@       @     �R@      �?     �C@      "@     �K@      *@      3@      @      8@     �F@      @      J@     �L@      N@      $@      6@      @      $@      5@              >@      �?      *@      @      $@      $@      @       @      @      $@      �?      (@      2@      7@      @      1@      @      @      0@              9@              (@      @       @      "@      @       @      �?      $@              (@      2@      4@      @      @       @      @      @              @      �?      �?      �?       @      �?       @              @              �?                      @              2@      (@      (@     �@@       @     �F@              :@      @     �F@      @      *@      @      4@     �A@      @      D@     �C@     �B@      @      1@      "@      "@      =@      @      C@              6@      @      E@      @      $@      @      3@      <@      @      C@      =@     �B@      @      �?      @      @      @      �?      @              @              @              @              �?      @               @      $@               @     @T@     �L@      >@     �T@      1@      M@      @     �S@      .@      T@     �B@      1@      &@      =@     @P@      >@     @X@     @V@     @^@      =@      @@      0@      (@      5@       @      7@      �?      0@      �?     �E@       @       @              @      9@      .@      B@      7@     �I@      @      3@      "@       @      3@              "@      �?      (@      �?      =@      @       @                      2@      (@      6@       @      B@      @      *@      @      @       @       @      ,@              @              ,@      @                      @      @      @      ,@      .@      .@       @     �H@     �D@      2@      O@      .@     �A@      @      O@      ,@     �B@      =@      .@      &@      9@      D@      .@     �N@     �P@     �Q@      8@      C@      =@      0@     �L@      ,@      <@      @      I@      ,@      A@      7@      ,@      @      2@     �A@      $@     �J@      M@      P@      3@      &@      (@       @      @      �?      @              (@              @      @      �?      @      @      @      @       @       @      @      @     `i@      O@      A@     `i@      .@     �r@             �^@      &@     �q@     �K@      @@      ,@      ?@     @c@      <@      p@      d@     �p@      D@      a@     �C@      5@      \@       @     @i@             �U@      @     �i@      7@      *@      @      *@     @V@      *@     `c@     �X@     @f@      B@      X@      :@      (@     @W@       @      b@             @R@      @     �`@      6@      $@      @      @     �S@       @     �_@     �R@      b@      ;@      L@      "@       @     �G@      @     �U@             �E@      �?      O@      &@      $@       @      @     �F@      @     @R@      ;@     �O@      4@      D@      1@      $@      G@      �?      M@              >@      @     �Q@      &@              �?       @     �@@      �?      K@     �G@     �T@      @      D@      *@      "@      3@              M@              *@      �?     �R@      �?      @       @      @      &@      @      <@      9@     �@@      "@      $@      @      @      �?              4@              @      �?       @      �?              �?      @      @              @      &@      "@      @      >@      $@      @      2@              C@              $@             �P@              @      �?      @       @      @      8@      ,@      8@      @     �P@      7@      *@     �V@      @      X@              B@      @     �S@      @@      3@      "@      2@     @P@      .@     �Y@     �N@     �V@      @     �B@      .@      $@      K@      �?     @R@              9@      @      L@      1@      3@      @      @     �G@      @      P@      B@     �L@             �A@      .@      $@     �I@      �?     �Q@              4@      @      K@      1@      3@              @     �G@      @      M@      B@     �I@               @                      @               @              @               @                      @                              @              @              >@       @      @     �B@      @      7@              &@      @      6@      .@              @      ,@      2@       @     �C@      9@      A@      @      9@       @             �B@       @      4@              "@      @      4@      "@              @      $@      1@       @      @@      3@      6@       @      @              @              @      @               @               @      @                      @      �?              @      @      (@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ~N�mhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�	���@�	           ��@       	                     @�&�n@           �@                            �?8k�v�@j           ��@                           �?u`?�@            ��@������������������������       �x(j@�             u@������������������������       ���<)�!@K           P�@                           �?3�%�@J            @]@������������������������       ����;f
@             I@������������������������       �.�<�Vj
@+            �P@
                          �:@�L�@�@�           ��@                           �?@�^�@S           ��@������������������������       ���u-9�@]             b@������������������������       ��(�-�@�            �x@                           �?��u�>6@b            `c@������������������������       ����Al�
@             :@������������������������       ��^�=i�@P             `@                          �4@�B�L#�@�           ��@                          �1@ġ\
?@�           |�@                           @��fZ�i@*           �}@������������������������       ����ҷ
@�            �m@������������������������       �L�I@G�
@�             m@                          �3@7/�#<@�           8�@������������������������       ����"0@)           �}@������������������������       ����@�            @m@                          �7@=���@�           ��@                           @���AR@;           �@������������������������       ��\2�>�@�             w@������������������������       ���D��Y@Y            �a@                           �?/4��W@]           H�@������������������������       ��� @�            @m@������������������������       �[䬱�@�            �s@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     �\@     �X@     Pu@      I@      |@      "@     �o@      <@     �z@      ]@     @P@      B@     �Q@     q@     �Q@     0v@     Pt@     P{@     �S@     �a@     �M@     �L@      c@      A@      _@      @     �`@      2@      a@      N@      C@      2@      G@     �_@      @@      a@     �b@     �b@      G@     @S@      C@      9@     @Y@      ,@      R@      @      R@      &@     �X@      8@      6@      &@      3@     �S@      8@     @R@     �R@     @Z@      @@      R@      @@      8@     @V@      &@     �M@      @     @P@      &@     @S@      8@      2@      &@      0@      P@      8@      Q@     �Q@     �W@      9@      =@      (@      (@      B@              :@      @      .@      @      A@      @      �?       @      @      :@       @      9@      >@     �I@      &@     �E@      4@      (@     �J@      &@     �@@      @      I@       @     �E@      1@      1@      "@      "@      C@      0@     �E@      D@     �E@      ,@      @      @      �?      (@      @      *@              @              5@              @              @      ,@              @      @      &@      @       @      �?              @              "@              �?               @              @               @                      @      @      @      @      @      @      �?      @      @      @              @              *@                              �?      ,@               @       @      @             �P@      5@      @@      J@      4@      J@      �?     �N@      @     �C@      B@      0@      @      ;@     �H@       @      P@     @R@      G@      ,@      I@      $@      9@     �C@      ,@     �I@      �?      I@      @      =@      <@      &@      @      7@      E@      @      M@      K@      9@      *@      1@      @      @      *@      �?      &@              2@       @      @      @      @                      .@              *@      3@      "@             �@@      @      2@      :@      *@      D@      �?      @@      @      8@      6@       @      @      7@      ;@      @     �F@     �A@      0@      *@      0@      &@      @      *@      @      �?              &@       @      $@       @      @      @      @      @      @      @      3@      5@      �?      @       @      �?                      �?              �?      �?      @      �?                       @                      �?      �?      @      �?      (@      "@      @      *@      @                      $@      �?      @      @      @      @       @      @      @      @      2@      .@             @e@      L@     �D@     �g@      0@     `t@       @     �^@      $@      r@      L@      ;@      2@      8@     @b@     �C@     @k@      f@     �q@     �@@     �O@      4@      2@     �[@      @     @h@              O@             @f@      5@      ,@      $@      @      K@      4@     @_@      Y@      e@      *@      8@      "@       @      <@      @      V@              5@              W@      @      @      @      @      4@      �?     �E@      E@     �P@      @      $@               @      @      @      K@              &@             �D@      �?      @      @      @      $@              6@      >@      =@      @      ,@      "@      @      6@              A@              $@             �I@       @                      @      $@      �?      5@      (@     �B@      �?     �C@      &@      $@     �T@             �Z@             �D@             �U@      2@      "@      @              A@      3@     �T@      M@     �Y@      @      ;@      @      @      N@              R@              <@             �P@      *@      @      �?              8@      ,@     @P@      ;@     �P@              (@      @      @      6@              A@              *@              4@      @      @      @              $@      @      1@      ?@     �B@      @     �Z@      B@      7@     �S@      &@     �`@       @      N@      $@      \@     �A@      *@       @      1@      W@      3@     @W@     @S@     @]@      4@     �J@      ,@      2@     �D@             �R@              :@       @     �G@      &@      "@      @      @     �G@      "@      I@     �D@     �B@      (@      D@      @      2@     �B@             �I@              3@      @      D@      @      "@      @      @     �@@       @      ?@      7@      =@      (@      *@      @              @              8@              @      @      @      @                      @      ,@      @      3@      2@       @              K@      6@      @     �B@      &@     �L@       @      A@       @     @P@      8@      @      @      $@     �F@      $@     �E@      B@      T@       @      9@      @      �?      2@      "@      :@       @      1@       @     �C@      @      �?      �?       @      *@      @      &@      0@      ;@      @      =@      0@      @      3@       @      ?@              1@              :@      2@      @      @       @      @@      @      @@      4@     �J@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��PhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @י4� @�	           ��@       	                    �?��n�@
           �@                           @���
�@�           ��@                          �:@8��U�@H           8�@������������������������       �2q���@!           �|@������������������������       �ɗ��6@'             N@                           �?S�� �@~           8�@������������������������       �3ݢ*�@�            �v@������������������������       ���+�uD@�            `o@
                           @f�43��@D           t�@                            @��6>�s@r           ��@������������������������       �3[H�c@�           8�@������������������������       �G���~@�            �q@                           @F@��q@�            �s@������������������������       ����?Q@�            �i@������������������������       �vp���
@M            �[@                           �?����6l@�           ��@                          �6@)ڨNІ@i           ��@                           @ 2~�}@@�            0v@������������������������       �U�� ��@D            @\@������������������������       ���O�@�            @n@                           @�rsn��@�            �m@������������������������       �s׾\��@y             j@������������������������       �p�)fQs@             <@                            �?�ݏ^1�@/           p�@                          �6@�����@�            @q@������������������������       ����&�@`            �c@������������������������       �B�s�ں@I             ^@                           @��"%�Y@�           Ђ@������������������������       ���n�K@"           �{@������������������������       ��*M��@d             d@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �b@      X@     �u@      B@     �z@      @     �l@     �D@     �{@     �Z@     �P@      D@     @U@     @o@     �P@     Pw@      t@     py@     �T@     `i@     �S@     �N@     �h@      ,@     ps@      @     �c@      8@     �s@     �Q@      A@      ;@     �F@     �c@      ;@     @l@     �f@      p@     �K@     @X@      @@      4@     �R@      "@     �d@      @     �S@      @     @b@      A@      &@      *@      (@      O@      "@      Y@      W@     @a@      =@     �E@      $@      ,@      <@      @      O@      @      B@      @      K@      8@       @      @      @      =@       @      M@      E@      O@      0@      E@       @       @      ;@      @     �N@      �?      ;@      @      G@      5@      @      �?      @      ;@       @     �K@      C@      O@      (@      �?       @      @      �?              �?       @      "@      @       @      @      �?      @               @      @      @      @              @      K@      6@      @     �G@      @     @Z@              E@      �?      W@      $@      @       @      @     �@@      �?      E@      I@      S@      *@     �B@      &@      @      :@      @     �Q@              8@             �E@      @      �?              @      8@              7@      ?@     �G@      *@      1@      &@      �?      5@             �A@              2@      �?     �H@      @       @       @      @      "@      �?      3@      3@      =@             �Z@      G@     �D@     �^@      @      b@       @     �S@      1@     �d@      B@      7@      ,@     �@@      X@      2@     �_@     �V@     �]@      :@      S@     �A@      ;@     �Y@       @     @\@             @P@      (@     �]@      6@      4@      $@      3@      T@      0@     �X@     @Q@     �W@      &@      J@      6@      0@     @T@             �T@              B@      @     @X@      ,@      $@      $@      @      P@      $@     �R@     �F@     @T@      @      8@      *@      &@      6@       @      >@              =@      @      5@       @      $@              .@      0@      @      9@      8@      *@      @      >@      &@      ,@      4@      @      ?@       @      *@      @      H@      ,@      @      @      ,@      0@       @      ;@      6@      8@      .@      *@      @      ,@      &@      @      ,@       @      &@      @      :@      (@       @      �?      ,@      &@       @      0@      2@      ,@      &@      1@      @              "@              1@               @              6@       @      �?      @              @              &@      @      $@      @     @`@      R@     �A@     `b@      6@      ^@      �?     �R@      1@     �`@      B@     �@@      *@      D@      W@      D@     `b@     `a@     �b@      ;@     @S@      6@      ,@     �R@      ,@     �F@      �?      9@      @      D@      3@      &@      @      @     �C@      ,@     �M@     �J@      P@      "@      C@      1@      @     �H@       @     �D@              ,@              6@      .@       @               @      2@      @     �A@      A@      F@      @      @      @      @      3@       @      "@              @               @              @                      @      @      $@       @      :@      �?     �@@      &@      @      >@              @@              $@              ,@      .@      @               @      .@              9@      :@      2@       @     �C@      @      @      :@      (@      @      �?      &@      @      2@      @      @      @      �?      5@       @      8@      3@      4@      @     �A@       @      @      7@      (@      @              $@      @      .@      @              @      �?      4@      @      6@      0@      4@      @      @      @              @                      �?      �?              @      �?      @                      �?      @       @      @                     �J@      I@      5@      R@       @     �R@              I@      (@     @W@      1@      6@      $@     �B@     �J@      :@      V@     �U@     �U@      2@      "@      <@      @      2@      @      ;@              2@      @      2@      @      @       @      $@      0@      @      8@      7@     �G@       @      @      $@      @      @              5@              "@      @      0@      @      @       @               @      �?      0@      "@     �A@      @      @      2@      �?      (@      @      @              "@               @       @                      $@       @      @       @      ,@      (@      @      F@      6@      .@      K@      @      H@              @@       @     �R@      (@      3@       @      ;@     �B@      5@      P@     �O@      D@      $@      B@      0@      ,@      F@      �?      ;@              6@       @     �N@      $@      3@      @      :@      <@      &@      G@      A@      <@       @       @      @      �?      $@       @      5@              $@              ,@       @              @      �?      "@      $@      2@      =@      (@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�o�shG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @Z#�X�@�	           ��@       	                   �6@�(Գ0@�           ��@                           @Ar���?@i           ԛ@                           �?1,�w��@{           ȕ@������������������������       ��_`�T@�           ��@������������������������       �l�ى�7@�           �@                           @Y��X��@�            0x@������������������������       �6Y�P@�            pt@������������������������       �J���l@'             N@
                           @�yc�@�           X�@                           �?�$��ڴ@C           �@������������������������       ���Q��@�            �x@������������������������       ����%�@I           `@                           �?c�r�@A            �Z@������������������������       �l�N�@            �A@������������������������       �������@-            �Q@                          �6@�~�#�@�           ��@                           @�/��@�           ��@                           �?ʿ��@@T           `�@������������������������       ���ޏc@�            �n@������������������������       �ڃEqE@�            �q@                           @�iX�1@A            �Z@������������������������       ���9��@             8@������������������������       ����1�@1            �T@                           @`��,TS@-            @                           @��
&@@�             v@������������������������       ����I@�            `k@������������������������       ��=fK	�@Q            �`@                           @Ԋ��`Z@T            @b@������������������������       �_i�S�@G            �^@������������������������       �����j@@             8@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        u@     `c@      \@     pu@      :@      ~@      @     `h@      8@     0~@     �Z@      O@      G@      N@     �p@      O@     �t@     t@     z@     @T@      l@     @Z@     �P@     0q@      .@     �v@      �?      ^@      .@     �v@     �O@     �I@      ;@      >@      g@      @@     @n@     `l@     0t@      L@     �]@     �J@     �C@     �g@      @     @q@             �T@      ,@      n@      @@      C@      $@      *@     @Z@      $@     �c@     ``@      l@     �C@     �U@      :@      =@     @c@      @      k@             @Q@      &@     �i@      :@      <@      @      "@     @U@      @     @^@     �U@     @g@      B@      C@      1@      @     �O@      @     @_@              B@             @[@      "@      ,@      @      @      F@      @     �M@      A@     �Z@      0@     �H@      "@      6@     �V@              W@             �@@      &@     @X@      1@      ,@      �?      @     �D@      @      O@     �J@      T@      4@      @@      ;@      $@     �A@      �?     �M@              ,@      @     �A@      @      $@      @      @      4@      @      C@      F@      C@      @      <@      7@      $@      A@      �?     �B@              ,@       @      A@      @      $@      @      @      3@      @      8@     �C@      A@       @      @      @              �?              6@                      �?      �?       @                              �?              ,@      @      @      �?     �Z@      J@      ;@     �U@      "@     �U@      �?     �B@      �?     �^@      ?@      *@      1@      1@      T@      6@     �T@      X@     �X@      1@      W@      F@      ;@     @U@       @      S@      �?      ?@      �?      ]@      ?@      *@      ,@      ,@     �Q@      1@     @R@      T@     �U@      1@      7@      ;@      2@      C@      @      6@      �?      4@             �H@      .@      $@      (@       @      @@      "@      >@      =@      B@      $@     @Q@      1@      "@     �G@       @      K@              &@      �?     �P@      0@      @       @      @     �C@       @     �E@     �I@      I@      @      ,@       @              �?      �?      $@              @              @                      @      @      "@      @      $@      0@      *@              "@       @                      �?       @                               @                                       @               @      @      @              @      @              �?               @              @              @                      @      @      �?      @       @      &@      "@             �[@      I@      G@      Q@      &@      ^@      @     �R@      "@     �]@     �E@      &@      3@      >@     �T@      >@     @V@     �W@     �W@      9@     �Q@      8@      6@     �D@      @     �W@       @      E@      �?      R@      6@      @      @      @      D@      "@      K@     �I@     �K@      &@     �O@      4@      2@     �@@      @     �Q@       @     �@@      �?      L@      6@      @      @      @      @@      "@      J@      E@      G@      "@      C@      @      "@      4@      @     �A@              ,@              1@      *@      �?       @      �?      &@      @      0@      6@      <@      @      9@      *@      "@      *@       @     �A@       @      3@      �?     �C@      "@      @      �?       @      5@      @      B@      4@      2@      @       @      @      @       @              8@              "@              0@                              @       @               @      "@      "@       @      �?              @      �?               @                              "@                                                              �?      �?              @      @      �?      @              0@              "@              @                              @       @               @       @       @       @      D@      :@      8@      ;@      @      :@      �?     �@@       @     �G@      5@      @      0@      7@      E@      5@     �A@     �E@     �C@      ,@      >@      *@      3@      4@      @      *@      �?      =@      @      8@      0@      @      &@      0@      ;@      $@      =@      E@      7@      *@      ,@      "@      $@      $@      @      "@      �?      3@      @      0@      &@      @              &@      7@      $@      ,@      =@      *@       @      0@      @      "@      $@      �?      @              $@      @       @      @              &@      @      @              .@      *@      $@      @      $@      *@      @      @       @      *@              @       @      7@      @              @      @      .@      &@      @      �?      0@      �?      "@      *@      @      @       @      *@              @       @      ,@      @              @      @      ,@      @      @      �?      (@              �?                      @                                              "@                                      �?      @      �?              @      �?�t�bub�s     hhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJUtGhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�Iԍd�@�	           ��@       	                     �?TO��K�@           ��@                           @«Q_�@C           p�@                          �;@�@�            �m@������������������������       �����<@}            �h@������������������������       ����o�@            �C@                           �?�Г	@�             r@������������������������       ��z:`�@7            �W@������������������������       �A=�UR@y            �h@
                          �?@P���w�@�           ��@                            �?)��/�@�           L�@������������������������       ������@�            �s@������������������������       ��u�A�U@�           ؆@                           @B!��@6            �U@������������������������       ��T��e�@             F@������������������������       �b�e}-@            �E@                          �6@���q"Z@�           ��@                           @F��u@�           ��@                           @DJڟ @,           ��@������������������������       ����4�{@`           ��@������������������������       ���jzO�@�            t@                           �?یr�N@�           ��@������������������������       �z3H
@�            @n@������������������������       ��7����
@�            Px@                           �?�ra5�M@�           �@                            @���0@�            @m@������������������������       ��a~%o	@~             h@������������������������       ��`�>�@            �D@                          �:@�v���@8           �@������������������������       ����o@�            @t@������������������������       ����4@j            �f@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     @^@     �R@     @w@     �B@     @}@      "@     @l@      ;@     p}@      \@     �P@     �C@      Q@     @m@     �O@     v@      s@     P|@     @T@     �a@      Q@     �G@      c@      =@     �`@      @     @_@      0@      d@     �I@     �@@      6@     �F@      Y@      =@      `@     �b@      f@      E@     �A@      4@       @     �P@      @      G@      @     �A@      @     @P@      @      &@      &@      (@      C@      @      6@      I@     �N@      2@      4@      (@      @      ;@       @      :@       @      1@       @      E@      @       @      @      @      "@      @      $@      *@      4@      @      4@      @      @      :@      �?      5@       @      .@       @     �B@      �?       @      �?      @       @      @      @      (@      4@      �?               @      �?      �?      �?      @               @              @      @               @       @      �?              @      �?               @      .@       @      �?      D@      @      4@      �?      2@      @      7@       @      @       @      @      =@      @      (@     �B@     �D@      .@      @              �?      (@      �?       @              @      �?      "@              @      @      �?      *@       @      @      (@      @      @       @       @              <@       @      (@      �?      ,@      @      ,@       @              @      @      0@      �?       @      9@      A@      $@      [@      H@     �C@     @U@      8@     @V@      @     �V@      "@      X@     �F@      6@      &@     �@@      O@      7@     �Z@     �X@     �\@      8@     �Y@     �@@      <@     �S@      8@     �U@      @     @V@      "@     @W@     �D@      4@       @      ?@      O@      4@     �Y@     �T@      [@      4@      >@      ,@      *@      @@      �?      =@      �?      2@       @      ?@      .@      @       @      @      2@      ,@      B@      &@      =@      @      R@      3@      .@     �G@      7@      M@       @     �Q@      @      O@      :@      0@      @      9@      F@      @     �P@      R@     �S@      ,@      @      .@      &@      @               @              �?              @      @       @      @       @              @      @      .@      @      @      �?      *@      "@       @                                                       @      �?      �?      �?              @      @      @      �?              @       @       @      @               @              �?              @       @      �?       @      �?                               @      @      @     �g@     �J@      <@     �k@       @     �t@      @     @Y@      &@     `s@     �N@     �@@      1@      7@     �`@      A@      l@     �c@     Pq@     �C@     �X@      @@      7@     @b@      @     �p@              S@       @     @j@      @@      :@      &@      @     @U@      3@     `c@     @Y@     �i@      4@     �K@      5@      ,@      X@      @     ``@              C@       @     @`@      :@      1@      @      @     �K@      2@     �W@     �N@     �Y@      ,@      C@      "@      @     �L@      �?     @W@              :@             �V@      2@      "@      @       @      A@      @      L@      B@     �P@      ,@      1@      (@       @     �C@       @      C@              (@       @     �C@       @       @      �?       @      5@      (@      C@      9@     �B@             �E@      &@      "@      I@      �?      a@              C@              T@      @      "@      @       @      >@      �?     �N@      D@     �Y@      @      8@      @      @      0@             �M@              2@              0@       @                       @       @      �?      5@      1@      F@      @      3@      @      @      A@      �?     @S@              4@              P@      @      "@      @              6@              D@      7@     �M@      �?     @W@      5@      @     �R@      @     �P@      @      9@      "@      Y@      =@      @      @      1@     �H@      .@     �Q@     �K@     �Q@      3@      6@       @      @      *@      �?      @@               @              B@      @                      @      6@      @      B@      *@      6@      "@      4@       @      @      *@              ;@              @              :@      @                      @      .@      @      @@      (@      3@      @       @                              �?      @              @              $@      �?                              @              @      �?      @      @     �Q@      3@       @     �N@      @      A@      @      1@      "@      P@      8@      @      @      &@      ;@      &@      A@      E@     �H@      $@     �I@      2@              I@              8@              @      @     �C@      $@      @      @      &@      1@      "@      2@      8@      <@      @      4@      �?       @      &@      @      $@      @      (@      @      9@      ,@      @      �?              $@       @      0@      2@      5@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��EBhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�ڧ��@�	           ��@       	                    @;�C@           ̙@                          �:@��\w@           �@                            @��;Z�y@p            �@������������������������       ���:CQ@h           �@������������������������       ���4!�@           �y@                            @M��b'@�            �l@������������������������       ��a66:@[            �a@������������������������       ���&B�@:            �U@
                            �?��˺@           �z@                          �3@�w��@�            �k@������������������������       ��>2*@             H@������������������������       ��9;�]n@i            �e@                           @G\^��`@�             j@������������������������       ���a@O            @_@������������������������       �}u�V@4             U@                           @Z�/4�[@�           ��@                          �4@8G{��@5           ��@                           @I���)@�           ��@������������������������       ��i$�N6@&           �|@������������������������       ���X�
@~             f@                          �6@-q�Sf@�           ��@������������������������       �(67{`�@�             k@������������������������       �n|Ë�@	           `z@                          �2@r�ɏ|�@_           Ȏ@                           �?"�&��
@�            �v@������������������������       �T��0`	@y             i@������������������������       �I}3+@d            `d@                          �;@�c6�@�           h�@������������������������       �<�}�@T           p�@������������������������       ��6S�Q@.            �O@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        u@      `@     @W@     �u@      B@     `~@      @     `m@      A@     �x@      X@      S@     �F@     �O@     �n@      M@      x@     �s@      |@     @U@     �^@      P@      L@      c@      :@     @b@      @     �[@      <@     �_@      K@     �G@      >@      C@     �]@      ;@     �c@     �b@     @c@     �C@     @W@      C@      A@      [@      5@     �[@      @     �S@      8@     �V@      H@     �B@      4@      8@     �V@      3@     �_@     @[@     �\@      ?@     �T@      5@      6@      V@      4@     �Z@       @     �K@      4@     �S@      C@      ;@      "@      6@     �R@      &@     �[@     �T@     �W@      ;@      K@      *@       @     �N@      @     �Q@       @      8@      $@      K@      &@      .@      @      @      E@      @     �P@      E@      Q@      ,@      =@       @      ,@      ;@      *@      B@              ?@      $@      9@      ;@      (@      @      1@      @@      @     �E@     �D@      :@      *@      $@      1@      (@      4@      �?      @      @      7@      @      (@      $@      $@      &@       @      0@       @      1@      :@      4@      @      @      "@      @      &@              @       @      3@              &@       @       @      $@      �?      *@      @      (@      *@       @      @      @       @      "@      "@      �?               @      @      @      �?       @       @      �?      �?      @      @      @      *@      (@              >@      :@      6@      F@      @      B@              @@      @      B@      @      $@      $@      ,@      <@       @      ?@     �C@      D@       @      ,@      1@      ,@      ;@      @      ,@              5@       @      .@              @      @      @      *@      @      "@      2@      :@      @      @              @      "@               @              @              �?               @                                      �?      @      $@              "@      1@      "@      2@      @      @              1@       @      ,@              @      @      @      *@      @       @      .@      0@      @      0@      "@       @      1@       @      6@              &@       @      5@      @      @      @      @      .@       @      6@      5@      ,@       @      &@      @      @      &@              0@              $@              2@       @       @       @       @      @              @      1@      $@      �?      @      @       @      @       @      @              �?       @      @      @      @      @      @      "@       @      0@      @      @      �?     �j@     @P@     �B@     �h@      $@     @u@      �?     @_@      @     �p@      E@      =@      .@      9@     �_@      ?@     @l@     �d@     `r@      G@     @\@      @@      3@     �]@      @     �h@              Q@      @      d@      ;@      2@      $@      ,@     �Q@      =@     �^@     @X@     �a@      >@     �B@      .@      "@      N@      �?      Y@             �@@             �S@      &@      @       @      @      A@      &@     �Q@     �J@     @Z@      &@      8@      @      "@     �E@      �?     �N@              6@             �K@      "@       @       @      @      6@      "@      O@      C@     @T@      &@      *@       @              1@             �C@              &@              7@       @      @                      (@       @       @      .@      8@              S@      1@      $@     �M@      @      X@             �A@      @     �T@      0@      *@       @      &@      B@      2@     �J@      F@      B@      3@      5@      @      @      (@      �?      J@              $@      @      >@      @      $@      @      �?      ,@      �?      4@      (@      $@      @     �K@      &@      @     �G@      @      F@              9@      �?      J@      *@      @      @      $@      6@      1@     �@@      @@      :@      ,@      Y@     �@@      2@     �S@      @      b@      �?     �L@       @      [@      .@      &@      @      &@      L@       @     �Y@      Q@      c@      0@      4@      &@      @      5@       @     �K@             �A@             �J@      �?      �?              @      2@       @     �C@      8@     �Q@       @       @               @      "@       @      <@              6@              >@              �?                      .@              9@      1@     �D@      �?      (@      &@      @      (@              ;@              *@              7@      �?                      @      @       @      ,@      @      >@      �?      T@      6@      (@      M@      �?     @V@      �?      6@       @     �K@      ,@      $@      @       @      C@              P@      F@     �T@      ,@     �R@      4@      @     �K@      �?     �T@              6@       @      K@      &@      "@      @      @      A@             �K@      E@     �P@      ,@      @       @      @      @              @      �?                      �?      @      �?      �?      @      @              "@       @      0@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�є0hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @=%<�B�@�	           ��@       	                    @�Y%k�@�           $�@                           �?e��UѰ@`           ��@                            �?��옖%@g           x�@������������������������       �ٮp�$�@�            �u@������������������������       �$���$Q@�           ��@                          �5@��|N�@�           ��@������������������������       ����m@           �z@������������������������       �)�S��@�            �v@
                           �?��o��@�           ��@                          �2@:0I7�y@�            �x@������������������������       ��ׯw%*@            �H@������������������������       �7�NNi@�            �u@                           @Z��;]@�           (�@������������������������       ���M�!�@9           0@������������������������       ��]1M�@g            @f@                           �?V���a}@�           ܐ@                           @�硜��@           |@                          �7@j��GT�@�            Pr@������������������������       �����	�@|            �g@������������������������       ��S,�@=            �Y@                           �?�a���8@[            �c@������������������������       �mv���	@             G@������������������������       ���	D��	@<            �[@                           @ػ��@�           ��@                           @Z�^�'�@P           �@������������������������       �_OXf��@'           �}@������������������������       ��զ$|@)            �Q@                          �4@���I�
@4            �T@������������������������       ��U�y�@             D@������������������������       ��uiR@            �E@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �a@      U@      w@     �I@     �}@      @     �n@     �@@     �|@     �X@      J@      ?@     @P@      n@      S@     Pv@     pr@     @{@     �Q@      m@      W@     �H@     0q@      9@     �w@      �?      d@      8@      u@     �N@     �C@      5@      C@      f@      I@     �p@      i@     �u@     �L@     �c@      E@     �A@     �c@      .@     `o@      �?     �X@      .@     `m@      @@      5@      1@      0@      ]@      ;@     `e@     @Y@     �k@     �@@     �S@      7@      6@     �W@      @     @a@             �J@      @     @]@      0@      *@      "@      $@     @Q@      @     @X@     �K@     �b@      .@      ?@      @      .@     �D@      @      ?@              <@      �?      F@      @      @      @      @      A@       @      5@      3@      F@      $@     �G@      1@      @     �J@      @     �Z@              9@       @     @R@      (@      "@      @      @     �A@      @      S@      B@     @Z@      @     �S@      3@      *@     @P@       @     @\@      �?      G@      (@     �]@      0@       @       @      @     �G@      4@     �R@      G@      R@      2@      <@      @       @     �C@       @      N@              4@      @     �R@      @      @       @              8@       @      K@     �A@     �F@      "@      I@      .@      &@      :@      @     �J@      �?      :@      @     �E@      (@      @              @      7@      (@      4@      &@      ;@      "@      S@      I@      ,@      ]@      $@      `@             �N@      "@     @Y@      =@      2@      @      6@     �N@      7@     �X@     �X@      `@      8@      >@      3@      $@     �D@      @     �@@              @@       @     �C@       @       @      �?      &@      5@      $@      9@     �C@     �K@      (@       @              @      @              "@              @               @      �?                      @              @                      &@              6@      3@      @     �A@      @      8@              =@       @     �B@      �?       @      �?       @      5@      @      9@     �C@      F@      (@      G@      ?@      @     �R@      @     �W@              =@      @      O@      ;@      $@      @      &@      D@      *@     @R@      N@     @R@      (@      ?@      4@      @     �P@      @      Q@              .@      @      F@      1@      @              &@      7@      $@     �K@     �F@      N@      (@      .@      &@              "@       @      ;@              ,@              2@      $@      @      @              1@      @      2@      .@      *@              X@     �H@     �A@     @W@      :@     �X@       @     �U@      "@     �^@      C@      *@      $@      ;@      P@      :@      V@     �W@     �U@      ,@     �E@      *@      .@     �C@      "@     �E@      �?     �E@      @     �H@      1@      @      @      @      3@      @      B@      E@     �G@      @      :@      $@      .@      :@      @      ;@      �?     �@@      @      9@      0@      @      @      @      $@      @      4@      :@      7@      @      1@      @      @      2@      @      ;@              .@              2@      @      �?      �?       @      @      @      2@      3@      1@      �?      "@      @       @       @      �?              �?      2@      @      @      "@      @      @      �?      @       @       @      @      @      @      1@      @              *@      @      0@              $@              8@      �?                              "@      �?      0@      0@      8@      @       @                      �?      @      @              @               @                                      @              @      @       @      @      "@      @              (@              &@              @              6@      �?                               @      �?      *@      *@      0@             �J@      B@      4@      K@      1@     �K@      �?     �E@      @     �R@      5@       @      @      8@     �F@      3@      J@     �J@      D@      @      D@     �A@      4@     �J@      1@      H@      �?      C@      @     �L@      5@       @      @      6@      @@      2@      G@     �E@     �A@      @     �A@      <@      4@      J@      (@     �A@      �?      B@      @      L@      3@      @      �?      3@      6@      (@      D@      D@      @@      @      @      @              �?      @      *@               @              �?       @      �?      @      @      $@      @      @      @      @              *@      �?              �?              @              @              1@                      �?       @      *@      �?      @      $@      @      �?      $@                                      @              @               @                              �?       @              �?      @      @              @      �?              �?                              �?              "@                      �?      �?      &@      �?      @      @      �?      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ_ɻhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���@�	           ��@       	                    @��-A@�           �@                           �?�j�@�           x�@                            @�V��h@>           @@������������������������       ��e�x@�            �s@������������������������       �m��B��@w             g@                          �;@j�4r7@�           P�@������������������������       ���si&�@n           h�@������������������������       ��uY�6�@M            @_@
                          �2@�5֯j@           0z@                          �1@��N�QJ@%            �N@������������������������       ��	��.@             E@������������������������       ��>:�[@             3@                           @�E�A@�@�            `v@������������������������       ���!�s@�             k@������������������������       �P8bwfT@Z            �a@                           �?�Oz�@�           �@                           �?_cP�e�@           �@                            @׌Cc2@            �|@������������������������       ���@�            �w@������������������������       �rW�m@1            �S@                          �8@"t{9�+@�             u@������������������������       ���@�            �q@������������������������       ���1Ld@$            �J@                            @8$8r^I@�           ��@                          �6@&�T�M@�           X�@������������������������       �ߪ!Ή0@�           �@������������������������       ���:��O@           P{@                           �?2,��O@�            Pq@������������������������       �.�B���
@[            �a@������������������������       �"Ca��@W            �`@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        v@      `@      W@      v@      D@     �}@      @     @m@      9@     @|@      [@      Q@      B@     �P@     @l@     �O@     �w@     �q@     �{@      T@     �_@     @P@     �M@      c@      ?@     �b@      @     �]@      1@      b@     �H@      F@      ;@     �F@      W@     �A@     �`@     @^@     �a@     �E@     @U@     �D@     �C@     @_@      :@     �\@      @     �T@      &@     @Z@      H@      >@      4@      ?@     �P@      :@      [@     �V@     �V@     �A@      =@      0@      *@      F@      @     �M@       @     �F@      @      M@      6@      (@      $@      $@      B@      @      F@      >@     �D@      .@      3@      *@      @      @@      @      C@              1@              D@      *@      &@      @      @      =@              9@      .@      ?@      (@      $@      @      @      (@              5@       @      <@      @      2@      "@      �?      @      @      @      @      3@      .@      $@      @      L@      9@      :@     @T@      5@      L@      @     �B@      @     �G@      :@      2@      $@      5@      ?@      5@      P@      N@      I@      4@      G@      .@      4@     @Q@      4@     �J@      @      9@      @     �E@      5@      2@      @      *@      :@      *@      J@     �G@      G@      3@      $@      $@      @      (@      �?      @       @      (@       @      @      @              @       @      @       @      (@      *@      @      �?      E@      8@      4@      <@      @     �@@              B@      @     �C@      �?      ,@      @      ,@      9@      "@      9@      ?@      J@       @      (@       @      @      $@              @              @              �?              �?                                              @      (@      �?      &@               @      @              @              @              �?              �?                                               @       @      �?      �?       @       @      @              �?               @                                                                               @      @              >@      6@      0@      2@      @      :@              =@      @      C@      �?      *@      @      ,@      9@      "@      9@      ;@      D@      @      ,@       @      ,@      0@              $@              6@      @      >@              @      @      @      ,@      @      (@      1@      >@      @      0@      ,@       @       @      @      0@              @      �?       @      �?       @      @       @      &@      @      *@      $@      $@       @      l@     �O@     �@@     �h@      "@     �t@              ]@       @     @s@     �M@      8@      "@      5@     �`@      <@     �n@     `d@     �r@     �B@      O@      (@      ,@     �O@             �_@             �I@      �?      W@      .@      @              @     �I@      @     �T@     �O@      `@      6@      @@       @      $@      ?@             @Q@              ?@              P@      $@      @              @      ;@       @     �A@      D@     �R@      2@      :@       @       @      :@             �N@              :@             �N@      "@                      @      1@      �?      A@      A@      M@      @      @               @      @               @              @              @      �?      @                      $@      �?      �?      @      1@      &@      >@      @      @      @@              M@              4@      �?      <@      @      �?               @      8@      �?     �G@      7@      K@      @      6@      @      @      =@             �H@              4@      �?      8@      @      �?                      8@              A@      6@      F@      @       @              �?      @              "@                              @                               @              �?      *@      �?      $@      �?     `d@     �I@      3@      a@      "@     �i@             @P@      @      k@      F@      4@      "@      .@     �T@      9@     @d@      Y@     �e@      .@     �`@      B@      .@     @Z@       @      f@              E@      @     �e@     �C@      3@      @      ,@      Q@      *@     �a@     �S@     �b@      &@      M@      5@      &@     @R@      �?      a@             �A@      �?     �\@      :@      .@      @       @      D@      @     @X@     �F@     �Z@      @     @S@      .@      @      @@      @      D@              @      @      M@      *@      @              (@      <@      @      F@      A@     �E@      @      <@      .@      @      ?@      �?      <@              7@             �E@      @      �?       @      �?      .@      (@      5@      5@      6@      @      &@      $@      �?      3@              *@              .@              <@      �?      �?                       @      @       @      &@      0@              1@      @      @      (@      �?      .@               @              .@      @               @      �?      *@      @      *@      $@      @      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJz��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�-����@�	           ��@       	                    �?Oi�Fi@�           ��@                          �8@��5�F�@l            �@                            �?����@�           �@������������������������       �HC�WN@�            �p@������������������������       ��??lۺ
@J           P@                           �?�d�h-e@w            �g@������������������������       ��`�@9             T@������������������������       �k0Q��@>            @[@
                           @��B|��@|           0�@                            �?L����@^           ��@������������������������       ���Z@e           x�@������������������������       �*��Q#@�           ��@                          �6@dT}M�@           ~@������������������������       ���U�[@�            `s@������������������������       ������L@c            `e@                           @��$k��@�           ��@                           �?� YE�@           ��@                           @��R6� @A           �@������������������������       �~u�Z*@            {@������������������������       ���g��F@6            �S@                          �4@��RxcH@�            �s@������������������������       �znн�@j             c@������������������������       ���p�y@d            �d@                          �3@���ې�@�            �s@                           @=�bv�@5             U@������������������������       ���� Ge @             &@������������������������       ���v�@.            @R@                           �?�#(�l<@�            @m@������������������������       �Im��@5            �S@������������������������       ������@g            `c@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       0s@      a@     @W@      v@      C@     p@       @      l@      :@     P}@     @W@     �Q@      G@     �S@     �o@     �O@     �w@     @q@     `y@     �V@     `i@     @V@     �J@     @p@      5@     @y@      @     @`@      ,@     @v@      J@      E@      @@     �I@      i@     �F@     Pp@      f@     �s@     �M@     �P@      6@      ,@      T@      @     �e@             �F@      �?     �`@      4@      (@      @      ,@     @P@      @     @X@     �N@     �^@      4@     �K@      1@      @      R@       @     �c@             �D@      �?     �Z@      *@       @              &@     �E@      �?      R@     �H@     @Z@      ,@      ;@      �?      @      :@             �H@              1@      �?     �B@      @      @              @      3@      �?      4@      2@      ;@      @      <@      0@      �?      G@       @     �Z@              8@             @Q@      @      @              @      8@              J@      ?@     �S@      $@      &@      @      "@       @       @      1@              @              <@      @      @      @      @      6@      @      9@      (@      1@      @       @      @      @      @      �?      @               @              &@      @      @       @               @       @      $@      @      @      @      "@              @      @      �?      ,@               @              1@                      @      @      ,@      �?      .@      @      *@       @      a@     �P@     �C@     �f@      1@     �l@      @     @U@      *@     �k@      @@      >@      :@     �B@     �`@     �D@     �d@      ]@     �g@     �C@     �V@      I@      ?@      b@      "@     `d@      @     @R@      *@     �a@      4@      8@      ,@      >@      Z@      B@     �[@     �S@     �c@      @@      >@      6@      0@     �N@      @      I@       @      9@      @      M@      @      &@      *@      4@      J@      &@      @@     �D@     �T@      .@     �N@      <@      .@      U@      @     @\@      �?      H@      @     �T@      ,@      *@      �?      $@      J@      9@     �S@     �B@     @R@      1@      G@      1@       @     �A@       @      Q@              (@             @T@      (@      @      (@      @      ?@      @      K@      C@      A@      @      0@      @      @      <@      �?     �K@              &@             @P@      @      @       @              4@             �@@      5@      <@      @      >@      $@      @      @      @      *@              �?              0@      @       @      @      @      &@      @      5@      1@      @      @      Z@      H@      D@     �W@      1@     �X@      @     �W@      (@     @\@     �D@      <@      ,@      ;@      K@      2@      ]@     �X@     �W@      ?@      Q@      <@      =@     �R@      0@      Q@      @     @R@      $@     �Q@      @@      5@      (@      6@     �C@      ,@      V@     @Q@      R@      4@      B@      0@      8@     �E@      *@      9@      @      F@      "@     �A@      0@      4@       @      2@      5@      "@      Q@      G@     �G@      $@      :@      ,@      5@      >@      @      6@      @     �B@       @      A@      .@      2@      @      0@      2@      "@      L@     �D@     �D@      $@      $@       @      @      *@      @      @              @      �?      �?      �?       @       @       @      @              (@      @      @              @@      (@      @      ?@      @     �E@              =@      �?      B@      0@      �?      @      @      2@      @      4@      7@      9@      $@      2@      �?              2@       @      <@              $@              2@      "@                      @       @      @      $@      (@      *@      @      ,@      &@      @      *@      �?      .@              3@      �?      2@      @      �?      @      �?      0@              $@      &@      (@      @      B@      4@      &@      4@      �?      ?@              6@       @      E@      "@      @       @      @      .@      @      <@      >@      6@      &@      @      @      "@      @              ,@              @              @      @                               @      @      @      (@      @      @              �?                              �?                              �?                                      �?                      @      �?              @       @      "@      @              *@              @              @      @                              �?      @      @      @      @      @      =@      1@       @      0@      �?      1@              3@       @     �A@      @      @       @      @      *@      �?      5@      2@      1@      @      $@      @              @              �?               @              1@      @      @      �?      @      �?      �?      @      @      @              3@      (@       @      "@      �?      0@              &@       @      2@       @      �?      �?       @      (@              0@      &@      ,@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�C7hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�����@�	           ��@       	                    �?��'a_�@�           x�@                            @4�H��@n           �@                          �7@��м@           Py@������������������������       �|T]�@�            Pq@������������������������       �MW��V@P             `@                           �?Aj�t�@j            �e@������������������������       �Bg����@,            @U@������������������������       ��|ik@>            @V@
                            �?���@�           l�@                           @���
@�            0r@������������������������       �w&�a�@�             p@������������������������       ��֤T�j@            �@@                            @��J�@�           ��@������������������������       �cu1yz@�            �l@������������������������       �#�uy^@B           ��@                          �5@�xf<�@�           ֡@                            �?i��u[�@f           p�@                           @rg#j��@            ��@������������������������       �'�uj�>@           �{@������������������������       �
�8s2@�            pw@                          �4@�bU�p�@f           X�@������������������������       �)tn�@2           P}@������������������������       ��~���G@4            �U@                          �9@1�6���@A           x�@                           @�&S�f@i           ��@������������������������       �@-�&��@           �z@������������������������       �;�HI�Z
@X            �`@                          �?@@+�P^b@�            �u@������������������������       �h'��n@�             s@������������������������       ���4L��@             F@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �r@      a@     �S@     Pv@      F@     @|@      "@     @o@     �E@     �|@     @`@     �P@     �B@     �J@     @m@      L@     0w@     `r@     �|@     @T@     @a@     �P@     �H@     `b@      ;@     �b@      "@     @`@      >@     �a@     �I@     �C@      *@     �@@     �W@      8@     �b@      `@     �d@     �F@     �F@      7@      5@     �L@      @      Q@      @      @@      @      F@      1@      "@      �?      @      C@      "@     �I@      H@     �T@      .@      <@      1@      $@     �C@      �?     �J@      �?      7@      �?      ?@      "@      @      �?      @      ?@       @      <@      ;@     �R@      &@      6@      @      @      >@      �?     �C@      �?      $@      �?      5@      @      @              @      ,@       @      4@      2@     �M@      "@      @      (@      @      "@              ,@              *@              $@      @      �?      �?       @      1@               @      "@      .@       @      1@      @      &@      2@      @      .@       @      "@      @      *@       @      @                      @      �?      7@      5@       @      @      "@              @      *@              @       @      @      @      @      @       @                      @      �?      @      $@       @       @       @      @      @      @      @       @              @      �?       @       @       @                       @              0@      &@      @       @     @W@      F@      <@     �V@      7@      T@      @     �X@      9@     @X@      A@      >@      (@      :@     �L@      .@     �X@     @T@     �T@      >@      6@      .@      @      >@       @      .@      @      B@      "@      9@      �?      &@      @      "@      1@      @      .@      8@      6@      .@      5@      $@      @      >@      @      .@      @      ?@      "@      0@      �?      "@      @       @      1@      @      *@      8@      5@      &@      �?      @      �?               @                      @              "@               @              �?                       @              �?      @     �Q@      =@      8@      N@      .@     @P@      @      O@      0@      R@     �@@      3@      @      1@      D@      &@      U@     �L@     �N@      .@      3@       @       @      4@      �?      4@      �?      2@      @      A@      @      &@              @      (@      @      =@      0@      *@      @      J@      5@      6@      D@      ,@     �F@       @      F@      *@      C@      :@       @      @      *@      <@      @     �K@     �D@      H@      $@     �d@     @Q@      >@     @j@      1@      s@              ^@      *@     �s@     �S@      <@      8@      4@     `a@      @@     �k@     �d@     �r@      B@     �T@      A@      0@      _@      @     @j@             �R@      @     �g@      B@      5@      *@       @      O@      *@     @a@     �[@     �j@      4@     �D@      :@      "@     �P@      �?     �Z@              A@      @     �[@      ;@      &@      *@      @     �D@       @     �X@     �P@     �a@      $@      (@      ,@       @      I@             �O@              $@             �M@      .@      @      @      @      6@       @      M@      @@     �Q@      @      =@      (@      �?      0@      �?     �E@              8@      @     �I@      (@      @       @              3@             �D@     �A@     �Q@      @     �D@       @      @      M@      @      Z@              D@             �S@      "@      $@              @      5@      @     �C@      F@     �R@      $@      B@       @      @     �H@      @     @V@              >@             �P@      "@       @                      1@      @      @@     �B@     @Q@      @      @                      "@              .@              $@              (@               @              @      @              @      @      @      @     �T@     �A@      ,@     �U@      *@     �W@              G@      $@      `@     �E@      @      &@      (@     @S@      3@     �T@      K@     @T@      0@     �G@      9@       @      M@       @      M@              <@      "@     �X@      5@       @      �?      @      J@      @      O@      @@     �B@      $@     �E@      ,@      @     �D@      �?      F@              :@      "@     �O@      3@       @      �?      @      G@      @      H@      <@      4@      "@      @      &@      @      1@      �?      ,@               @             �A@       @                       @      @      �?      ,@      @      1@      �?     �A@      $@      @      <@      &@      B@              2@      �?      >@      6@      @      $@      @      9@      (@      5@      6@      F@      @      4@       @      @      <@      "@      ?@              2@      �?      9@      4@      @      $@      @      7@      (@      *@      5@     �E@      @      .@       @                       @      @                              @       @                      �?       @               @      �?      �?        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ5R6EhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @)��x6�@�	           ��@       	                     �?��Tf�@�           ��@                           �?v�tgt@_           ��@                           �?�Z�Ƨ@�           0�@������������������������       �-W��� @�            �m@������������������������       �,�ᶲ(@           �{@                           �?�'�G��@�           Ė@������������������������       ��d���@x           ��@������������������������       ���E:�@0            �@
                           �?��@��U@}           p�@                          �6@!t���@�             q@������������������������       ��s#�	@r            �h@������������������������       ���S�5@2            �S@                           @�h�Ѩ�@�            �u@������������������������       ��}�A@�            pr@������������������������       �բGBP@!            �J@                           �?�$�oE�@�           �@                          �:@���|V"@�           p�@                          �3@Bf��ʓ@\           ��@������������������������       �����x@            �k@������������������������       ���B �@�            �u@                           �?ɳ�?�@\             c@������������������������       �r]�T&@             ;@������������������������       ���D��@L            @_@                           �?�mQo�d@           `{@                           @�5�]ă@�             m@������������������������       �rw�[1}
@+            �S@������������������������       ���֚6
@\            `c@                           @U��ufN@�            �i@������������������������       �`�� I�@b            `a@������������������������       �����p@,            �P@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       `s@     �`@     �V@     �u@      D@     @}@      @     `m@      9@     ~@     @W@     �M@      E@     �T@      l@     �R@     �v@     0t@      |@      Q@     �i@     �T@     �J@     �o@      8@     v@      @      d@      .@     �u@      J@      E@      9@      G@      e@      F@     @o@     �j@     �v@     �H@      d@     @S@      E@      h@      5@     �n@      @     @^@      $@     �p@      G@      >@      8@     �D@     �`@      D@     @h@     �e@     �p@      C@     �D@      (@      5@     �P@       @     @X@             �F@      �?      Z@      &@      @      @      @     �G@      @     �M@     �F@     �W@       @      (@      @      "@      9@      @      .@              5@      �?      =@       @      @      @       @      2@      �?      :@      8@      <@      @      =@       @      (@      E@      @     �T@              8@             �R@      @                      @      =@       @     �@@      5@     �P@      @      ^@     @P@      5@     @_@      *@     �b@      @      S@      "@     �d@     �A@      ;@      4@      A@     �U@     �B@     �`@     @`@     �e@      >@      I@      ,@      &@     �G@       @     @Q@      @      ?@      @      S@      0@      @      @      $@     �E@      .@     @P@      G@     �O@      $@     �Q@     �I@      $@     �S@      @     @T@      �?     �F@      @     �V@      3@      5@      .@      8@     �E@      6@     �Q@      U@     �[@      4@     �F@      @      &@     �N@      @     �Z@             �C@      @     @T@      @      (@      �?      @     �A@      @      L@      D@     �W@      &@      :@      �?      �?      3@       @      I@              ;@      @      :@      @       @      �?      �?      ,@              .@      5@     �G@      @      *@                      &@       @      H@              7@      �?      5@       @       @              �?      @              $@      (@     �B@       @      *@      �?      �?       @               @              @      @      @      �?              �?              "@              @      "@      $@      @      3@      @      $@      E@      �?      L@              (@             �K@      @      @              @      5@      @     �D@      3@      H@      @      .@      @      @     �D@      �?     �E@              (@             �G@              @              �?      5@      @      B@      0@     �C@      @      @              @      �?              *@                               @      @                      @                      @      @      "@              Z@     �H@      C@     @W@      0@     �\@      �?     �R@      $@     @`@     �D@      1@      1@      B@     �L@      ?@      \@      [@     �U@      3@     �O@     �@@      :@     �I@      ,@     �P@      �?     �C@      $@     �M@     �@@      ,@      *@      >@      B@      5@      S@     �Q@      G@      0@     �F@      8@      3@      C@      "@      P@              =@      "@     �J@      9@      @      "@      7@      :@      &@      R@      L@     �@@      .@      4@      @      "@      0@              ?@              $@              3@      $@              @      �?      .@      @      =@      7@      2@      @      9@      2@      $@      6@      "@     �@@              3@      "@      A@      .@      @      @      6@      &@      @     �E@     �@@      .@      $@      2@      "@      @      *@      @       @      �?      $@      �?      @       @       @      @      @      $@      $@      @      .@      *@      �?       @      �?       @      �?               @      �?      �?      �?      @       @                       @                      �?              �?      �?      $@       @      @      (@      @                      "@              @      @       @      @      @      $@      $@      @      .@      (@             �D@      0@      (@      E@       @     �H@              B@             �Q@       @      @      @      @      5@      $@      B@     �B@     �D@      @      1@       @      @      9@      �?      8@              :@             �E@      �?       @                      "@      @      1@      5@      >@      �?       @      @      �?      *@              �?              (@              .@      �?       @                       @      @      @       @       @              "@      @      @      (@      �?      7@              ,@              <@                                      @              &@      *@      <@      �?      8@       @      @      1@      �?      9@              $@              <@      @      �?      @      @      (@      @      3@      0@      &@       @      0@       @              0@      �?      1@              @              3@      @              @      @      @      �?      *@      ,@      @      �?       @              @      �?               @              @              "@      �?      �?      �?              @      @      @       @      @      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ>�7mhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?ǡ��	�@�	           ��@       	                    �?ơYV@           �@                           @�z�L��@l           0�@                          �9@eO8��@           `z@������������������������       ��r	Y@�            @u@������������������������       ���8n�@4            �T@                           �?�<���@_             d@������������������������       �n`�p�@             �K@������������������������       ��>�v$@?            @Z@
                           �?v4��9@�           ؐ@                           �?���X��@�            @x@������������������������       ����nI�@�             u@������������������������       ����h�@!             I@                          �;@}WmBe@�           ��@������������������������       �,��@@L           H�@������������������������       ��}E[�@d             e@                           �?,���@�           ��@                           �?��	��@�           X�@                            @v�I�@           �y@������������������������       ��m���
@�            `t@������������������������       ��}��h@7            �T@                           @�SqF�}@�             w@������������������������       ��(C��
@�            �l@������������������������       �1�v[�
@U            `a@                           @-�՘�V@�           �@                           @�|��X@�           Ȅ@������������������������       ��/;��S@�            �q@������������������������       ��{p�˰@�            �w@                            �?/"7���@           H�@������������������������       ��u'��@-           �}@������������������������       ��R��@�            u@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       `t@     �`@     �X@     �u@     �F@     0|@      2@     �m@      6@     �|@     �W@     �R@     �G@     �P@     �p@      Q@     `v@     �r@     �y@      V@      c@     �R@     �N@     �`@     �@@     �`@      .@     @`@      1@      f@     �E@     �E@      6@     �C@     @Z@     �A@     @^@      a@      b@     �E@      K@      :@      ?@      G@      @      K@      @      B@      �?     �O@      &@      *@       @      "@      D@      ,@     �C@     �F@     @S@      &@     �G@      $@      6@     �C@       @      E@      @      ;@      �?      B@      "@      *@       @      @      8@      &@      ;@      =@      N@      "@     �D@      @      1@      ?@       @     �C@      @      0@              <@      @      &@              @      1@      $@      6@      8@      K@      "@      @      @      @       @              @      @      &@      �?       @      @       @       @              @      �?      @      @      @              @      0@      "@      @      �?      (@              "@              ;@       @                      @      0@      @      (@      0@      1@       @      @      @      @      @              �?                               @       @                       @      @              @       @      @      �?      @      *@      @      @      �?      &@              "@              3@                               @      $@      @      @       @      (@      �?     �X@     �H@      >@     @V@      >@      T@       @     �W@      0@     @\@      @@      >@      4@      >@     @P@      5@     �T@      W@     �P@      @@      8@      (@      &@      7@      @     �A@              F@      @     �K@      .@      &@       @      (@      9@      @      @@     �D@      6@      &@      8@      (@      $@      2@      @      <@             �D@      @     �J@      .@      @       @      @      7@      @      ?@      8@      6@       @                      �?      @              @              @               @              @              @       @              �?      1@              @     �R@     �B@      3@     �P@      :@     �F@       @      I@      &@      M@      1@      3@      2@      2@      D@      1@      I@     �I@     �F@      5@     �L@      2@      $@      G@      7@     �F@      @     �B@      &@     �F@      ,@      .@       @      (@      <@      "@     �D@     �A@     �D@      3@      1@      3@      "@      4@      @              �?      *@              *@      @      @      $@      @      (@       @      "@      0@      @       @     �e@     �M@      C@      k@      (@     �s@      @      [@      @     �q@      J@      ?@      9@      ;@     �d@     �@@     �m@      d@     �p@     �F@      J@      ,@      .@     �R@      @      a@              C@      �?     �\@      1@       @              @      G@       @      T@      K@     �Y@      4@      :@      @      &@     �A@      @      S@              5@             �L@      @      �?              @      4@       @      >@      ?@     @P@      .@      7@      @      "@      <@             @P@              (@             �H@      @                      @      .@              <@      9@     �H@      "@      @               @      @      @      &@              "@               @       @      �?                      @       @       @      @      0@      @      :@      @      @     �C@              N@              1@      �?      M@      &@      �?              @      :@              I@      7@      C@      @      (@      @      @      9@             �F@              @             �D@      $@      �?              �?      $@              B@      .@      1@      @      ,@       @              ,@              .@              *@      �?      1@      �?                      @      0@              ,@       @      5@             �^@     �F@      7@     �a@      "@     �f@      @     �Q@      @     �d@     �A@      =@      9@      4@     �]@      ?@     �c@     �Z@      d@      9@     �L@      6@      @      M@       @     @T@             �@@      �?     �X@      1@      ,@      0@      @     �K@      @     @Q@      E@      S@      "@      9@      .@      �?      A@       @      @@              ,@      �?     �A@      @      �?      @      @      ;@      @      @@      1@      <@      @      @@      @      @      8@             �H@              3@              P@      (@      *@      &@              <@      �?     �B@      9@      H@      @     @P@      7@      2@      U@      @      Y@      @     �B@      @      Q@      2@      .@      "@      1@     �O@      9@      V@     @P@     @U@      0@     �B@      2@      &@      J@      @     �C@              ,@              A@      1@      @      @      (@      A@      1@     �K@     �H@     �L@       @      <@      @      @      @@             �N@      @      7@      @      A@      �?       @      @      @      =@       @     �@@      0@      <@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�2oyhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @���k��@�	           ��@       	                    �?��?	�#@�           �@                           �?�=9�Q@M           ��@                          �7@���	W@�            Pu@������������������������       �G�!�}9@�            �l@������������������������       ����"k�@C            �[@                          �:@�6�d@}           ؂@������������������������       ��(J8k@5           �~@������������������������       �ǴY�cM@H            �\@
                           @߄7�9@�           p�@                           �?-\��_@�           l�@������������������������       �0~���@�            w@������������������������       �d��@�           P�@                           @��!��r@           �@������������������������       ����)?�@�           �@������������������������       ��k��Y
@|            �g@                           �?��$�E�@�           ��@                          �3@���+�@�            �u@                           �?&u���
@]             b@������������������������       ����2*
@.            �P@������������������������       ��+���@/            �S@                          �4@�'�lt@�            �i@������������������������       �ˤ��/
@             9@������������������������       ����N�@{            �f@                          �6@B!�/��@�           ��@                          �1@/����^@�            �x@������������������������       ������@8            �V@������������������������       �O�*�$�@�             s@                           �?�ޥ!X[@�            @u@������������������������       ��n�e^@�            �o@������������������������       ��eO11@9             V@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       pv@     `a@     @U@     Pu@      B@      }@      @     `k@     �A@     �|@     @Z@      K@      @@     @U@     �n@     �N@     `u@      s@     �|@      V@     �p@      W@     �M@     �p@      7@     0u@      @     `a@      4@     �u@      P@     �@@      3@      I@      f@     �G@     �o@     `i@     `w@      L@     @S@      J@      >@      U@      *@     @Q@       @     �M@      *@     @W@      5@      (@      &@      9@      O@      4@     �Q@     �P@     �a@      5@      4@      *@      &@      =@      @     �@@              9@      �?     �F@      .@      @      @      @      2@       @      ;@      4@      K@       @      ,@      @      �?      6@       @      ;@              0@      �?      :@      @      �?              @      *@              7@      0@      G@      @      @      @      $@      @      �?      @              "@              3@      $@      @      @              @       @      @      @       @      @     �L@     �C@      3@     �K@      $@      B@       @      A@      (@      H@      @      @      @      3@      F@      2@      F@     �G@      V@      *@      J@      @@      $@     �E@      $@      B@      �?      9@      &@      E@      @      @      �?      0@      @@      *@     �D@     �C@      P@      *@      @      @      "@      (@                      �?      "@      �?      @      @      �?      @      @      (@      @      @       @      8@             �g@      D@      =@     �f@      $@     �p@      �?      T@      @     �o@     �E@      5@       @      9@     �\@      ;@     �f@      a@      m@     �A@     �V@      :@       @     �]@       @     ``@             �H@      @      d@      ;@      4@      @      0@      O@      9@     �W@     �Q@     @^@      4@     �A@       @      @      9@             �N@              5@             �K@       @       @              @      5@       @      C@      :@      H@      (@     �K@      2@      @     �W@       @     �Q@              <@      @     �Z@      3@      2@      @      (@     �D@      7@      L@     �F@     @R@       @     �X@      ,@      5@     �N@       @     `a@      �?      ?@      @     �W@      0@      �?       @      "@     �J@       @     �U@     @P@     �[@      .@     �R@      $@      5@     �E@       @     @Z@      �?      <@      @     �S@      ,@      �?       @       @      >@      �?      P@     �E@     �W@      ,@      8@      @              2@              A@              @      �?      0@       @                      �?      7@      �?      7@      6@      1@      �?     @W@     �G@      :@     @S@      *@     @_@      �?      T@      .@     �[@     �D@      5@      *@     �A@     �P@      ,@     �V@     @Y@      U@      @@      B@       @      "@      3@      �?      G@              C@      @      :@      ,@       @              @      =@      @      >@      ?@      ;@      (@      1@       @      @       @              A@              1@              @       @                      �?       @      �?      ,@      ,@      (@               @       @      @      @              (@              $@              @      @                              @              "@              @              "@                      @              6@              @               @      @                      �?       @      �?      @      ,@      @              3@      @      @      &@      �?      (@              5@      @      4@      @       @              @      5@      @      0@      1@      .@      (@      @      �?                      �?       @                      �?                      @                      @      @               @      @      �?      0@      @      @      &@              $@              5@      @      4@      @      @              @      2@       @      0@      .@      &@      &@     �L@     �C@      1@      M@      (@     �S@      �?      E@      "@      U@      ;@      *@      *@      >@      C@       @      N@     �Q@     �L@      4@      A@      0@       @      =@      @      O@              8@             �K@      &@      @      �?       @      8@       @     �C@      A@      @@      $@       @      @              $@      �?      @              @              1@      @      @              �?       @              .@      �?      @       @      :@      $@       @      3@      @     �L@              5@              C@      @      @      �?      �?      0@       @      8@     �@@      ;@       @      7@      7@      "@      =@      @      1@      �?      2@      "@      =@      0@      @      (@      <@      ,@      @      5@      B@      9@      $@      *@      .@      "@      5@      @      $@      �?      .@       @      *@      "@      @      "@      <@      &@      @      .@      >@      3@      "@      $@       @               @       @      @              @      �?      0@      @              @              @      �?      @      @      @      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJnnwhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?T��J�~@�	           ��@       	                     �?��62�@9           l�@                          �3@[�L@B           �@                           @�p�]R@~            `i@������������������������       ��Y^N��
@d            �c@������������������������       �����Q�@             F@                          �=@6�RD��@�             s@������������������������       ��S*�=@�            @q@������������������������       ��q�.Zw
@             <@
                           �?T���o@�           ��@                            @���;��@=           �~@������������������������       �+�$�	@�            u@������������������������       �t�e+�@k            �c@                           �?��ӂ@�           ��@������������������������       �xa�@�            �k@������������������������       �L��:M�@&           P}@                           �?� >���@|           \�@                           @%@x��@�           ��@                           �?Y�i�@S           P�@������������������������       �`-V8��@�            �r@������������������������       �_�[*(�@�           ��@                           �?囒��@Q            �`@������������������������       �ݑ�V�
@             D@������������������������       ��2eN�R@7            @W@                          �6@�¾g�&@�           ��@                          �2@��,Μ;@�           p�@������������������������       ��j\LR�@�            �w@������������������������       ��E��@
           Py@                            �?8�k?>@�            w@������������������������       �n�%z0s@A             Y@������������������������       ��q��:@�            �p@�t�b�/     h�h5h8K ��h:��R�(KKKK��h��B`        t@     �b@     @W@     pw@      =@     P}@      *@      m@      >@     �{@     �T@     �O@      >@     �R@     @m@      I@     �y@     �q@     `|@     �R@      d@      J@     �E@     �d@      .@     �l@      @     @Y@      ,@     �f@      ?@      4@      ,@       @     �Z@      0@      c@      ^@     �k@      >@     �H@      ;@      0@      K@      @      M@      @      B@      �?     �R@      @      @      $@      @      ?@      @      D@      >@      G@      &@      $@      (@      @      9@              <@              &@              >@      �?       @                      &@              4@      *@      @@      @      "@      "@       @      .@              9@              $@              >@      �?       @                      "@              0@      @      6@       @      �?      @       @      $@              @              �?                                                       @              @      @      $@       @     �C@      .@      (@      =@      @      >@      @      9@      �?      F@       @      @      $@      @      4@      @      4@      1@      ,@      @     �B@      $@      @      =@      @      =@      @      7@             �D@       @      @      "@      @      0@       @      4@      .@      ,@      @       @      @      @                      �?               @      �?      @                      �?      �?      @      �?               @                     �[@      9@      ;@     @\@      (@     �e@       @     @P@      *@     @[@      <@      *@      @      @     �R@      *@     @\@     �V@      f@      3@     �D@      @       @      @@      �?     �T@      �?      @@      �?      I@       @      @       @      @      >@      �?     �H@     �C@     �W@      $@      8@       @       @      5@             �O@              1@              D@      @      �?              �?      0@      �?      A@      =@     �R@       @      1@      @      @      &@      �?      4@      �?      .@      �?      $@      @       @       @       @      ,@              .@      $@      4@       @     �Q@      3@      3@     @T@      &@     @V@      �?     �@@      (@     �M@      4@      $@       @      �?     �F@      (@      P@     �I@     �T@      "@      <@      @      2@      1@      @      5@              "@      @      .@      "@      @              �?       @      @      5@      4@      6@      @      E@      ,@      �?      P@      @      Q@      �?      8@      @      F@      &@      @       @             �B@      @     �E@      ?@      N@      @      d@      X@      I@      j@      ,@     �m@      @     �`@      0@     @p@      J@     �E@      0@     �P@      `@      A@     p@     �d@      m@     �F@     �R@     �L@      ?@     �]@      *@     �T@      @     @S@      .@     �Y@      7@      ?@      $@     �C@      K@      2@      Y@     �U@     @Y@      ?@     @Q@      B@      =@     �[@       @      O@      @      Q@      .@     @V@      7@      7@       @     �A@      I@      .@     @V@     �T@     @V@      ?@      >@      @      @     �A@       @      6@              >@      �?      :@      "@      @      @      $@      1@      @     �@@      6@      <@      @     �C@      ?@      7@     �R@      @      D@      @      C@      ,@     �O@      ,@      1@      �?      9@     �@@       @      L@      N@     �N@      9@      @      5@       @       @      @      4@              "@              *@               @       @      @      @      @      &@      @      (@               @      @              @       @      @              �?              @                                       @      �?      @      @      @              @      .@       @      @      @      *@               @              "@               @       @      @       @       @       @      �?      @             @U@     �C@      3@     �V@      �?     �c@             �K@      �?     �c@      =@      (@      @      ;@     �R@      0@     �c@      T@     ``@      ,@      H@      5@      (@     @P@      �?     �]@             �C@      �?      ]@      0@      "@      �?      @      I@      @      \@      N@     �V@       @      9@      $@      @      ;@             �O@              8@             @R@      "@      @              @      2@      @     �C@      5@      F@      @      7@      &@      @      C@      �?      L@              .@      �?     �E@      @      @      �?              @@       @     @R@     �C@      G@      @     �B@      2@      @      9@              C@              0@              E@      *@      @      @      4@      8@      "@     �F@      4@     �D@      @       @      @      @      @              &@              @              @      @              �?      "@       @      @      2@       @      0@              =@      .@      @      4@              ;@              (@              C@      "@      @      @      &@      0@      @      ;@      2@      9@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ%�4hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����@�	           ��@       	                    �?��G#�@�           P�@                            �?64B�@�@d           Ȁ@                           �?�"t l/@�            @t@������������������������       �������@L            �^@������������������������       ���q��@�            @i@                           �?�ר�9�@�            �j@������������������������       �کi��y@?            @X@������������������������       �؆/�d@M             ]@
                           @���o�@�           �@                          �:@];�J�@O           ��@������������������������       ��mtd�@�           P�@������������������������       �u����h@�            �p@                            �?��t	�z@E            �Y@������������������������       �����'
@             ?@������������������������       �S�Q̊$@2             R@                          �5@�6�4f�@�           �@                          �3@��Ŀ�@�           H�@                            @$Ԓ�@u           X�@������������������������       ���X��^@           �@������������������������       ���Ñ_@r            �e@                           �?D�٣į@-           p~@������������������������       �Ř�h�@}            �h@������������������������       ��9j�@�            r@                           @�g3P�@$           �@                          �9@|Y9YO�@A           �@������������������������       �'�v`�@�            �s@������������������������       ��f�!s@y            �h@                          �6@���2��@�            v@������������������������       �-x�%��
@/             U@������������������������       �T8�B��@�            �p@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       x@      a@     �U@     �u@     �B@     @}@      $@     �l@      ?@     0{@     �^@      J@      B@      Q@      o@      N@     �u@     �r@     `{@     @R@     @b@     �P@     �K@     `b@      5@     �a@      "@      ]@      6@     �_@     �I@      <@      9@      E@     @[@      ;@     `a@     @a@      f@      B@     �K@      3@      1@     �K@      @     �N@      @      9@      @     �E@      2@      "@      @      @     �B@      @     �H@     �G@      N@      ,@      ;@      "@      (@      B@             �C@              (@      @      >@      $@      @      @       @      8@      @      ;@      <@      E@      @      (@      �?      @      $@              0@              @              (@       @       @       @              (@      �?      @      .@      4@              .@       @      @      :@              7@               @      @      2@       @      @      @       @      (@      @      4@      *@      6@      @      <@      $@      @      3@      @      6@      @      *@      �?      *@       @      @              �?      *@       @      6@      3@      2@      @      0@      @      @      @       @       @              "@              @      @                      �?      @       @       @      &@      $@      �?      (@      @      �?      *@      @      ,@      @      @      �?       @      @      @                      @              ,@       @       @      @     �V@     �G@      C@      W@      0@     �S@      @     �V@      1@     �T@     �@@      3@      4@     �C@      R@      4@     �V@     �V@     @]@      6@     �R@      C@     �B@      V@      .@     �Q@      @     �T@      1@      S@      @@      0@      0@      =@     �P@      ,@     �S@     �U@     �\@      4@     �M@      0@      9@      L@      ,@     �Q@      @     �E@      ,@     @P@      9@      (@       @      4@      H@      @     �N@      N@      V@      2@      0@      6@      (@      @@      �?               @      D@      @      &@      @      @       @      "@      3@      @      1@      ;@      ;@       @      0@      "@      �?      @      �?       @               @              @      �?      @      @      $@      @      @      (@      @       @       @      @      @      �?              �?       @              @              @              �?       @      @                      �?              �?              *@      @              @              @              @               @      �?       @       @      @      @      @      &@      @      �?       @     �m@     �Q@      @@      i@      0@     �t@      �?     �\@      "@     Ps@      R@      8@      &@      :@     �a@     �@@      j@      d@     Pp@     �B@      [@      D@      1@     �_@      @     �j@              S@       @     `j@      B@      2@      @      (@     �Q@      7@     @b@      Y@      h@      5@     @R@      2@      .@     �U@       @     �c@              K@             �b@      4@       @      �?      @      L@      ,@     @V@      H@     @`@      (@     �C@      .@       @     @R@             ``@             �F@             @`@      *@      @      �?      @      H@      @     �R@      C@     �]@      (@      A@      @      @      *@       @      ;@              "@              3@      @      �?              �?       @      @      ,@      $@      (@             �A@      6@       @     �D@      @     �K@              6@       @      O@      0@      $@      @      @      .@      "@     �L@      J@     �O@      "@      *@      "@      �?      8@              1@              $@              8@      $@      �?               @      @              6@      3@      B@      @      6@      *@      �?      1@      @      C@              (@       @      C@      @      "@      @      @      &@      "@     �A@     �@@      ;@      @     ``@      ?@      .@     �R@      &@     �\@      �?      C@      @     �X@      B@      @      @      ,@     @Q@      $@     �O@      N@      Q@      0@      U@      2@      @     �A@       @     �R@              >@      @      O@      3@      @               @      F@       @     �@@      ?@      H@      (@     �N@      (@      @      4@       @      E@              2@      �?     �D@      (@                      �?      ?@              9@      8@      3@      @      7@      @      �?      .@      @      @@              (@       @      5@      @      @              �?      *@       @       @      @      =@      "@     �G@      *@      $@     �C@      @     �D@      �?       @      @      B@      1@       @      @      (@      9@       @      >@      =@      4@      @      (@              �?      @      �?      2@              @       @      (@      @                              $@      �?      @       @      @             �A@      *@      "@     �@@       @      7@      �?      @       @      8@      &@       @      @      (@      .@      @      9@      ;@      1@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�JhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?m��p5�@�	           ��@       	                   �:@�7X��@           P�@                           @G�9�V5@(           |�@                            @j}�g8@           �@������������������������       �B��\.�@�           ȅ@������������������������       �n��޶z@P           `�@                             @3��0�@             :@������������������������       ��QUL>. @             .@������������������������       ��}�F��?             &@
                            �?���q��@�            Pw@                          �=@��4d˱@F            �]@������������������������       �c��+7�@%             P@������������������������       �M�����@!             K@                           @����@�            �o@������������������������       ����9j@I             [@������������������������       ��6�|n@`            `b@                          �6@��E��H@�           �@                           @�X<��@�           ��@                            �?��ʢ4M@p           ��@������������������������       � ;��ќ
@�            �p@������������������������       �6�TFy@�           @�@                           @��d��@g           �@������������������������       �9�񗠁@           �{@������������������������       �Hߗ챕
@T            �`@                           �?���@@�           �@                            �?C�r@�            �n@������������������������       �k!_�
@\            �a@������������������������       ���w�^@B            @Z@                           @�l}w�@#           p|@������������������������       �#"K�z@�            p@������������������������       ����8(@�            �h@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     `a@     �S@     �u@      ?@     �|@      @     `n@      ,@     0z@      [@     �K@      A@     @R@     �k@     �R@     �x@      t@     �}@      V@     @a@     @Q@     �K@      `@      6@      a@      @     �]@      &@      b@     �H@      >@      7@     �G@     �W@     �B@      e@     �`@      e@     �C@      ]@     �A@      ?@     �Y@      3@      `@      @     �U@      &@      ^@     �@@      6@       @      @@      Q@      ;@     `a@     @Y@     �`@      @@     �\@      ?@      ?@     �Y@      2@      `@      @     �T@      &@      ]@     �@@      6@       @      @@      Q@      :@      `@     @Y@     ``@      @@     @P@      5@      *@      P@      @      R@      @      C@      @     �S@      "@      .@      @      .@     �D@      ,@     �R@      J@     �U@      3@      I@      $@      2@      C@      &@      L@             �F@      @      C@      8@      @      @      1@      ;@      (@      K@     �H@      F@      *@      �?      @                      �?                      @              @                                              �?      &@              �?                      @                                                              @                                              �?      @              �?              �?      �?                      �?                      @                                                                      @                              6@      A@      8@      ;@      @      "@      �?      @@              9@      0@       @      .@      .@      ;@      $@      =@      @@     �B@      @       @      ,@      @      @              @              *@               @      @              "@      "@      @      @       @      $@      &@      @              �?       @      @                              @              @       @              @      @      @      @      @       @      "@      �?       @      *@      �?      �?              @               @              @      @              @       @              �?      @       @       @      @      4@      4@      5@      4@      @      @      �?      3@              1@      &@       @      @      @      4@      @      5@      6@      :@      @      @      "@      $@      *@      �?      �?      �?      @                      "@      @      �?      @       @      @      (@      "@      $@      �?      ,@      &@      &@      @       @      @              .@              1@       @      @      @      @      (@              "@      *@      0@       @      h@     �Q@      8@     �k@      "@     �s@             @_@      @      q@     �M@      9@      &@      :@     �_@     �B@     �l@     �g@     �r@     �H@     �Y@      C@      2@     `c@      @     `p@              W@      �?      i@      <@      5@       @      "@     @U@      :@      e@     �]@      l@      ?@      K@      6@       @     �Z@             @e@             �I@      �?      `@      1@      1@      @      @     �F@      8@     �[@      T@     �b@      7@      @       @      �?      A@             �I@              (@              C@      @      �?      @      �?      1@      �?      8@      &@      I@      (@     �G@      4@      @      R@             �]@             �C@      �?     �V@      (@      0@      �?      @      <@      7@     �U@     @Q@     �X@      &@     �H@      0@      $@     �H@      @      W@             �D@              R@      &@      @      @      @      D@       @      M@      C@      S@       @      E@      @      $@      D@      @     �O@              A@              M@      $@      @       @      @      ;@       @     �B@      :@     @Q@      @      @      "@              "@              =@              @              ,@      �?              �?              *@              5@      (@      @      @     @V@      @@      @     @P@      @     �L@             �@@       @     �R@      ?@      @      @      1@      E@      &@      O@     �Q@     �S@      2@      =@      �?      @      1@       @      @@              &@              >@      (@      @                      6@              9@      2@      ;@      *@      3@      �?       @      @              4@               @              .@              �?                      $@              5@      *@      4@      @      $@               @      $@       @      (@              @              .@      (@       @                      (@              @      @      @      "@      N@      ?@       @      H@      @      9@              6@       @      F@      3@      �?      @      1@      4@      &@     �B@     �J@     �I@      @      9@      4@      �?      B@      �?      ,@              2@      �?      :@      (@      �?              @       @      "@      8@      >@      6@      @     �A@      &@      �?      (@      @      &@              @      �?      2@      @              @      &@      (@       @      *@      7@      =@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�>hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��%���@�	           ��@       	                   �5@���!@�            �@                            @�zG�t@�           �@                          �4@��W�8�@           �z@������������������������       �a�:�@�            �t@������������������������       �����-�@A            �W@                           �?D�WA$V@�            �q@������������������������       ��ӟ�z@:            �U@������������������������       �H	v���@w            @h@
                           @CW��y|@.           (�@                           �?�["�@�           Ѓ@������������������������       �����u@p             g@������������������������       ��8,\�@            |@                          �;@���=�@�            �p@������������������������       �������@l            �e@������������������������       ��̷1�@8             W@                          �3@�"o#�@�           �@                           @��Nl�@v           Ў@                            @���P^D@�           ��@������������������������       �L71�5�
@�           �@������������������������       ��x��@b             c@                           �?J^��@�            �l@������������������������       �Q��4�@<            �W@������������������������       ��̍Tm@P            �`@                           �?���Oa@>           ��@                            @w=L6-�@�           p�@������������������������       ����f�@=           @������������������������       �zi$�i4@S            @_@                           @=�E�@�           ȅ@������������������������       ���ŧ�x@           �|@������������������������       ���2��@�            `m@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       Ps@     �]@     @W@     �v@     �I@     p|@      &@     �j@     �@@      |@     �V@     �Q@     �B@     @T@     @p@      Q@     �x@     �q@     @{@     @W@     @[@     �N@      M@     `a@     �@@     @`@      &@      ]@      :@     `b@      E@      D@      1@     �H@     �[@      C@     �c@     @`@     �b@      F@      M@      &@      .@     @U@      0@      R@              C@      @     �Q@      ,@      2@      �?      ,@      H@       @      R@     @P@     �R@      4@     �@@      @      @      O@      @      D@              3@      @      I@      @      ,@              @      ?@      @      B@      A@     �I@      2@      =@      @      @      H@      @     �@@              .@      @     �D@      @       @               @      7@      @      1@      :@     �F@      1@      @      @              ,@              @              @      �?      "@              @              @       @              3@       @      @      �?      9@      @      "@      7@      *@      @@              3@       @      4@      "@      @      �?      "@      1@      �?      B@      ?@      8@       @      @      @      @      &@              @               @      �?      &@      @      �?                      @      �?      $@      &@      &@              3@              @      (@      *@      ;@              1@      �?      "@      @      @      �?      "@      &@              :@      4@      *@       @     �I@      I@     �E@      K@      1@      M@      &@     �S@      3@     @S@      <@      6@      0@     �A@      O@      >@     @U@     @P@      S@      8@     �@@      A@      ?@     �F@      &@     �E@      &@      K@      0@      F@      ;@      4@       @      ;@     �E@      6@      K@     �H@      E@      4@      2@      "@      .@      (@              :@      �?      .@      @      *@      @      @      �?      @      .@      @      (@      @      &@      @      .@      9@      0@     �@@      &@      1@      $@     �C@      (@      ?@      5@      1@      @      7@      <@      .@      E@     �E@      ?@      ,@      2@      0@      (@      "@      @      .@              8@      @     �@@      �?       @       @       @      3@       @      ?@      0@      A@      @      .@       @      @       @      @      *@              *@      @      <@              �?      @      @      .@      @      3@      @      5@              @       @      @      �?               @              &@              @      �?      �?      @      @      @       @      (@      &@      *@      @      i@      M@     �A@      l@      2@     Pt@             �X@      @     �r@      H@      ?@      4@      @@     �b@      >@     �m@     `c@     �q@     �H@     �J@      6@      *@      W@      @     @e@              H@             @d@      &@      "@      @      "@      O@      (@     @\@      I@     �a@      *@      C@      @      @      S@      @     @a@             �E@             �^@      $@       @      @      @     �G@      @     �T@      D@     �[@      (@      7@      @      @     �L@      �?     �[@             �@@              Y@      @       @      @       @      D@      @      Q@     �A@     �X@       @      .@      �?      �?      3@      @      <@              $@              7@      @                      @      @       @      .@      @      (@      @      .@      .@      "@      0@              @@              @             �C@      �?      �?              @      .@      @      >@      $@      =@      �?      @       @      @      @              (@               @              ,@                                      "@      �?      &@      "@      $@      �?      "@      @      @      "@              4@              @              9@      �?      �?              @      @      @      3@      �?      3@             `b@      B@      6@     �`@      ,@     `c@             �I@      @     `a@     �B@      6@      1@      7@      V@      2@     @_@     @Z@      b@      B@     �R@      *@      "@      O@      "@     @S@              :@      @     �Q@      :@      @      &@      "@     �E@      (@      D@      J@      L@      4@      O@      $@      @      F@       @     �R@              0@      @     �E@      8@       @      &@      "@     �B@      &@      @@      D@      G@      0@      *@      @       @      2@      �?      @              $@      �?      ;@       @      @                      @      �?       @      (@      $@      @      R@      7@      *@     �Q@      @     �S@              9@      �?     @Q@      &@      0@      @      ,@     �F@      @     @U@     �J@     @V@      0@     �D@      0@      @     �M@      @      O@              8@      �?      F@      @       @      @      @      :@      @      K@      C@      I@      "@      ?@      @      @      &@              0@              �?              9@      @       @       @      $@      3@              ?@      .@     �C@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�G-hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B                              @�e���@�	           ��@                           �?�
r�Le@            0�@                          �@@�\���@^           x�@                            �?f�U9�@O           ��@������������������������       �yZ��@!           �{@������������������������       ����5�@.           �}@������������������������       �(����@             ;@                          �4@d� 'w@�           ��@	       
                    @�1�@y           ��@������������������������       ��c�Uv@�           �@������������������������       �~��ΎB@�            �s@                          �=@׻LV@)           P�@������������������������       �A\Y��@�           ��@������������������������       ��V*�@�@4            �V@                          @@@�bP��@�           Đ@                           @d�M��@�           P�@                           @`^+��@U           P�@������������������������       ��� �@�           ��@������������������������       �%Z�}@k            `e@                           @�rZm�@A            �Z@������������������������       ���@
@             �I@������������������������       ���#M@!            �K@������������������������       ��f�p̔@             =@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       0u@     �_@      Z@     �t@     �I@     �}@      &@     `j@      C@     �{@      \@     @P@      A@      K@      n@     @P@     �v@     �r@     `{@      [@     �m@     @V@      L@     0p@     �A@     0x@      @     �`@      :@     �t@      Q@      D@      4@      @@     �f@     �H@     @p@     @j@     0u@     �R@     @S@     �E@      =@      W@      2@      V@      @      L@      0@     �W@      :@      1@      @      ,@      O@      ;@     @R@     �O@     �Z@      >@     @S@      D@      :@     �V@      2@      V@      @     �H@      0@     �W@      :@      ,@      @      ,@      N@      8@     @R@     �M@     �Z@      >@      C@      5@      @      I@      (@      C@      @      <@      *@      A@      "@      @      @      &@     �B@      $@      ;@      6@     �J@      3@     �C@      3@      3@      D@      @      I@      �?      5@      @     �N@      1@       @      @      @      7@      ,@      G@     �B@     �J@      &@              @      @       @                              @                              @                       @      @              @                     @d@      G@      ;@     �d@      1@     �r@      @     �S@      $@     �m@      E@      7@      *@      2@     �]@      6@     `g@     `b@      m@     �F@      L@      1@      $@      Z@      @     �c@             �I@      @     @b@      ,@      .@      @       @     �I@      "@     @Y@     �S@     �b@      *@     �F@      "@      @     �M@      @     �Z@             �C@       @     @^@      @      @      @       @      A@      @      P@      H@     @Z@       @      &@       @      @     �F@       @     �J@              (@       @      9@      "@      &@                      1@      @     �B@      >@     �F@      @     �Z@      =@      1@     �O@      (@     �a@      @      <@      @     @W@      <@       @      @      0@     �P@      *@     �U@     @Q@     �T@      @@     �X@      =@      &@     �N@      @     �`@              <@      @      V@      6@       @      @      (@     �O@      (@     �R@     �M@     �Q@      ;@       @              @       @      @      @      @                      @      @                      @      @      �?      &@      $@      *@      @      Y@      C@      H@     @Q@      0@      W@      @      S@      (@     �[@      F@      9@      ,@      6@      N@      0@     �Y@      W@     �X@     �@@     �X@      A@      E@     @Q@      *@      W@      @      S@      (@     �[@      C@      9@      $@      5@      N@      0@     @Y@     �V@     �X@     �@@     @W@      ;@      D@     �K@      *@     �U@      @     �P@      (@     �X@     �B@      5@      @      1@      J@      0@     �X@     @T@     �U@      9@     �P@      :@     �C@     �D@      &@      Q@      @      M@      (@     �Q@      >@      4@      @      1@     �F@      ,@     �S@     �P@     �Q@      7@      ;@      �?      �?      ,@       @      3@               @              <@      @      �?                      @       @      4@      .@      1@       @      @      @       @      ,@              @              $@              &@      �?      @      @      @       @               @      $@      &@       @              @              @              @              @              @      �?                      �?       @                      @      @      @      @               @      $@                              @              @              @      @      @      @               @      @      @      �?      �?      @      @              @                                      �?      @              @      �?                      �?      �?      �?        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ���8hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?t��5�@�	           ��@       	                   �<@��e��@/           ��@                          �3@�؛�x^@�           ȗ@                           @�k�i�@1           �~@������������������������       �����@�            �x@������������������������       �=�Q~�
@9             W@                          �:@�앲�@�            �@������������������������       ��)�C,�@           ��@������������������������       �[���8�@f            @e@
                           �?��&�9h@y            �e@                          @@@���T\@             E@������������������������       �k^{Q�	@             =@������������������������       �XL��J@             *@                           @4��Q��@^            �`@������������������������       �	��F�@2            �R@������������������������       ��e��@,            �L@                           �?)!�B�L@|           R�@                          �7@S��Ŝ+@           ��@                           @l,��@�           �@������������������������       �+}�+F@�             p@������������������������       �I�Y*@�            x@                           @a��߉@x            `g@������������������������       �}�U˹@8             W@������������������������       ��z�E	@@            �W@                           �?�*�8ݱ@d           ��@                           @��\%I2@{           �@������������������������       �^u&�@�             w@������������������������       �W��I�@�            `n@                           @��#5S�@�           P�@������������������������       ��M:�<@�             s@������������������������       � &����@-           �}@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �`@      [@      x@      D@      }@      @      o@      B@     p}@      W@     �O@      8@     @Q@      m@      N@     0v@     �q@     �{@      P@     @`@     @R@     @Q@     �e@      :@     `b@      @     �a@      6@      d@      I@     �A@      .@      E@     �[@     �A@     @^@      `@     �f@      >@      ]@      J@      K@     @d@      9@     �a@      @      `@      4@     �b@     �C@     �A@       @     �A@     �X@      ;@     @\@     �\@     @e@      =@     �A@      "@      6@     �M@      @     �K@       @      :@      @     �D@      1@       @      �?      @     �A@      @     �A@     �G@      S@      @      :@      @      (@      H@      @      E@       @      .@      @      D@      (@       @      �?      @     �@@      @      >@      B@     �P@      @      "@      @      $@      &@              *@              &@              �?      @                               @              @      &@      $@             @T@     �E@      @@     �Y@      6@     �U@       @     �Y@      0@     @[@      6@      ;@      @      ?@     �O@      6@     �S@     �P@     �W@      7@     �R@     �B@      @@      S@      2@     �T@      �?     @R@      .@      X@      1@      4@      @      =@      K@      0@     @P@      L@     �R@      4@      @      @              ;@      @      @      �?      >@      �?      *@      @      @      �?       @      "@      @      *@      &@      3@      @      ,@      5@      .@      &@      �?      @              (@       @      &@      &@              @      @      (@       @       @      .@      *@      �?      �?      @       @                      @                              @      @               @      @      @       @      �?      @      @              �?       @       @                      @                              @      �?               @      @      @                              @                       @                                                                      @                                       @      �?      @      �?              *@      1@      *@      &@      �?      �?              (@       @      @      @              @       @      "@      @      @      &@       @      �?      @      (@      &@       @      �?      �?              "@       @       @      @              �?              @      @      @      @      �?              @      @       @      "@                              @              @      �?              @       @      @      �?       @      @      @      �?      i@      O@     �C@     �j@      ,@     �s@      �?      [@      ,@     `s@      E@      <@      "@      ;@     �^@      9@     @m@     �c@     0p@      A@      S@      @      0@     �P@      @     @_@              F@      @      ^@      ,@       @               @      H@      @     �U@      L@      _@      2@      J@      @      0@     �N@       @     @Y@              ?@      @     �V@      $@      @              @      A@      �?     �R@      B@      Z@      *@      ,@      @       @      ;@             �E@              @              C@       @      @              @      &@      �?      A@      (@      D@      &@      C@       @       @      A@       @      M@              9@      @     �J@       @                      �?      7@              D@      8@      P@       @      8@      �?              @      @      8@              *@              =@      @      @              @      ,@       @      *@      4@      4@      @      *@      �?              @      @      &@              "@              @       @      @                      (@      �?      @      "@      $@      @      &@                      �?              *@              @              9@       @                      @       @      �?      "@      &@      $@       @     @_@      L@      7@     `b@       @      h@      �?      P@      &@     �g@      <@      4@      "@      3@     �R@      6@     `b@     �Y@     �`@      0@     �N@      :@      @     @R@      @     �T@      �?      @@       @     �S@      @      @      @      @      D@      @     �M@     �G@      O@      @      ?@      .@      @      D@      @      I@              7@       @      F@      @      @       @      @      3@      @      B@      8@      G@      @      >@      &@      �?     �@@      @      @@      �?      "@              A@      @      �?      �?              5@              7@      7@      0@      �?      P@      >@      1@     �R@       @     �[@              @@      @      \@      5@      0@      @      *@      A@      3@      V@     �K@     @R@      "@     �@@      .@      @      7@       @      D@              ,@             �I@       @      @      �?       @      &@      @      9@      9@      ?@      "@      ?@      .@      *@     �I@             �Q@              2@      @     �N@      *@      $@      @      &@      7@      .@     �O@      >@      E@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                              @�Ob�t@�	           ��@       	                   �4@HP��W@�           إ@                           �?��wzn@2           H�@                            �?BQ��c�@�            pt@������������������������       ��\B8@k            @e@������������������������       �gMC2\�@c            �c@                           �?�j_h7�@d           X�@������������������������       �$u�z�
@-            ~@������������������������       �)�~#�@7           �~@
                           �?Yڟ��@�           h�@                          �?@7ҡ�v@�           ��@������������������������       �8&��@q           ��@������������������������       ���U��5@#            �L@                            �?e훼��@"           (�@������������������������       ��挥��@�           ��@������������������������       �8"6�@�            @n@                          �5@z�b)�@�           t�@                           �?�Zl^�@R           p�@                           @H.,�؁@�            0q@������������������������       ����,�@�            �k@������������������������       �V�ّ�@             K@                           @IoI�@�            �q@������������������������       ��qHן@�            pp@������������������������       ��|J��@             4@                          �@@�8	�H�@_           x�@                          �:@|�+x@P           ؀@������������������������       ��c�R�4@�            Pw@������������������������       �SX��k@a            �d@������������������������       �+�\;� @             4@�t�bh�h5h8K ��h:��R�(KKKK��h��B        Pv@     �_@     �U@     �u@     �G@     `}@      &@     `m@      7@     �|@     @X@     @R@      <@     �K@     @l@     �G@     �x@     �s@     @{@     @S@     �n@     �V@     �L@     �o@      4@     @w@       @     �`@      0@      v@     @Q@     �G@      3@      @@     `d@     �A@     �q@     @h@      v@     �L@     �U@      8@      :@     �\@      �?     `j@              M@      @      g@      5@      8@      "@              R@      $@     �a@     �Y@     �e@      ?@      >@       @      .@      >@             �@@              *@      @      H@      @      $@      @              7@      @      1@      8@      G@      .@      "@      @      @      2@              6@               @              9@       @      @      @              3@      �?      @      *@      2@      "@      5@      @      $@      (@              &@              @      @      7@      �?      @                      @       @      $@      &@      <@      @      L@      0@      &@      U@      �?     @f@             �F@      �?      a@      2@      ,@      @             �H@      @     �_@     �S@      `@      0@     �@@      (@      @      F@              W@              ,@             @P@      @      @      @              4@             �J@     �H@     @Q@      &@      7@      @      @      D@      �?     �U@              ?@      �?     �Q@      (@      $@       @              =@      @     @R@      >@      N@      @     �c@     �P@      ?@     `a@      3@      d@       @     @S@      $@      e@      H@      7@      $@      @@     �V@      9@      a@     �V@      f@      :@     �A@     �@@      3@     �K@      $@     �H@      @     �D@      @     �P@      (@      .@      @      3@     �A@      &@     �P@      G@     @U@      (@      A@      9@      @      I@      $@     �F@      @      ?@      @     �P@      (@      *@      @      2@      A@       @     @P@      G@     @T@      $@      �?       @      (@      @              @              $@              �?               @      �?      �?      �?      @       @              @       @     �^@      A@      (@      U@      "@      \@       @      B@      @     @Y@      B@       @      @      *@      L@      ,@     �Q@     �F@      W@      ,@      Y@      >@      @     �F@      "@      R@              =@       @     @Q@      ?@      @      @      $@     �B@      $@     �G@     �@@     @S@      "@      7@      @      @     �C@              D@       @      @       @      @@      @      �?              @      3@      @      7@      (@      .@      @     @\@      B@      =@     �W@      ;@     �X@      @      Y@      @     �[@      <@      :@      "@      7@     �O@      (@     �\@     @^@      U@      4@     �K@      ,@      ,@     �G@      (@     @R@      �?      J@      �?      O@       @      (@      �?      @      A@      @      I@     �M@     �H@      @     �@@      @      @      @@      @     �A@              @@              7@      @      @      �?              (@      �?      7@      :@      ?@      @      =@      @      @      7@      @      :@              9@              2@      @      @      �?              $@      �?      7@      8@      3@      �?      @      �?      �?      "@              "@              @              @                                       @                       @      (@       @      6@      "@      "@      .@       @      C@      �?      4@      �?     �C@      @       @              @      6@      @      ;@     �@@      2@       @      6@      @      "@      .@       @     �A@      �?      4@      �?      C@      @       @              @      2@       @      6@     �@@      2@      �?              @                              @                              �?                                      @      @      @                      �?      M@      6@      .@     �G@      .@      9@       @      H@      @      H@      4@      ,@       @      4@      =@      @      P@      O@     �A@      .@     �L@      1@      *@      G@      ,@      9@       @      H@      @     �G@      ,@      ,@      @      3@      =@      @      P@      O@     �A@      .@     �C@      (@      &@      ;@      "@      5@              8@      @      B@      (@       @      @      0@      1@      �?      J@     �E@      5@      ,@      2@      @       @      3@      @      @       @      8@      �?      &@       @      @      �?      @      (@      @      (@      3@      ,@      �?      �?      @       @      �?      �?                                      �?      @               @      �?                                                �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ<�^>hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?5�f���@�	           ��@       	                    �?g��O9@'           �@                           @�;�;l@n           ��@                          �<@���I�@�            `v@������������������������       �`��% @�            0t@������������������������       �@4oG]
@            �A@                           @w"G�(@�            �i@������������������������       ��x�k>�
@,            �R@������������������������       �T`�I�@X            @`@
                           �?<n��&@�            �@                           @�3'Y�@            |@������������������������       �j��q��@m            �e@������������������������       ���؆l
@�            0q@                          �5@����@�           0�@������������������������       �w�54�@�            �w@������������������������       ���ى�u@�            �p@                           �?P>��^1@�           ��@                            @�Y?[@�           �@                          �;@E�Y8@�           8�@������������������������       �g��h:@H           P�@������������������������       �Y���r@F            @_@                          �3@^ gCF@           �{@������������������������       �V���g@:             V@������������������������       �2�'�u@�            0v@                          �1@8}��@�           0�@                           @*��m`�	@�            �k@������������������������       ���]��@:            �U@������������������������       ��e��	@R             a@                          �>@��5.K@T           h�@������������������������       ���e�mG@?           X�@������������������������       �;�5�;@             A@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@     ``@     �Y@     �t@      D@     �}@      @      l@     �A@     �{@     �\@     @Q@     �E@     @U@     �p@     �N@     Pw@      r@     {@     @R@     �b@     �E@     �D@     �`@      .@      n@      @      X@      .@     �j@      J@      7@      1@      5@     �Y@      4@     �_@      `@      h@      =@      L@      ,@      9@      D@      @     �P@      @      A@      @      F@      7@      1@      $@      .@      =@      @      I@     �G@      P@      (@      @@      $@      .@      .@             �L@      @      2@      @     �A@      4@      *@      $@      @      1@      �?     �B@      9@     �@@      "@      @@      @       @      .@              L@       @      (@       @      A@      ,@      *@      "@      @      .@      �?      A@      7@     �@@      "@              @      @                      �?      �?      @      �?      �?      @              �?      �?       @              @       @                      8@      @      $@      9@      @      "@              0@       @      "@      @      @              $@      (@       @      *@      6@      ?@      @      .@       @       @      &@      @       @              @              @                                      @      �?      �?       @      @              "@       @       @      ,@       @      @              $@       @      @      @      @              $@      @      �?      (@      ,@      8@      @      W@      =@      0@      W@      "@     �e@              O@      $@     `e@      =@      @      @      @     �R@      1@      S@     @T@      `@      1@      B@       @      @      ?@      @     @P@              9@             �S@      &@      �?              @      A@       @     �B@      ?@     �P@      &@      $@      �?      @      $@      @      7@              @              ?@      @      �?              @      .@      �?      2@      2@      ,@      $@      :@      @      �?      5@              E@              3@             �G@      @                              3@      �?      3@      *@     �J@      �?      L@      5@      &@     �N@      @     @[@             �B@      $@     @W@      2@      @      @      �?      D@      .@     �C@      I@     �N@      @      .@      (@      @     �A@             @P@             �@@              O@      @      @      @              5@       @      ;@      <@     �I@      @     �D@      "@      @      :@      @      F@              @      $@      ?@      .@              @      �?      3@      @      (@      6@      $@       @      e@      V@      O@      i@      9@      m@      �?      `@      4@      m@      O@      G@      :@      P@     �d@     �D@     �n@      d@      n@      F@      T@      F@      C@     �\@      3@     �T@      �?      Q@      1@     �V@      =@      @@      1@      I@      P@      7@     �\@     �R@     �Z@      :@     �K@      ?@      2@     �V@      @      G@              B@      @      M@      (@      .@      $@      6@     �C@      .@      P@     �A@     �Q@      3@     �G@      :@      2@     @Q@      @      F@              <@      @     �H@      &@      "@      @      0@     �A@      .@     �F@      5@     �L@      1@       @      @              5@               @               @              "@      �?      @      @      @      @              3@      ,@      ,@       @      9@      *@      4@      8@      *@      B@      �?      @@      (@      @@      1@      1@      @      <@      9@       @      I@      D@      B@      @      @       @      @      @      �?      "@              @              @      @                      �?      @              $@      (@      3@              2@      &@      .@      5@      (@      ;@      �?      ;@      (@      :@      ,@      1@      @      ;@      4@       @      D@      <@      1@      @      V@      F@      8@     �U@      @     �b@              N@      @     �a@     �@@      ,@      "@      ,@     �Y@      2@     �`@     @U@     �`@      2@      *@      @      @      0@              K@              .@             �D@              �?      �?      �?      "@       @      5@      .@      :@       @      @      �?              $@              4@               @              .@                              �?      @              ,@       @      (@      �?      "@       @      @      @              A@              *@              :@              �?      �?              @       @      @      *@      ,@      �?     �R@     �D@      5@     �Q@      @      X@             �F@      @     @Y@     �@@      *@       @      *@     �W@      0@      \@     �Q@      [@      0@     @R@      D@      .@     @Q@      @      W@             �F@      @     @Y@     �@@      *@       @      *@     �W@      0@      Z@     @Q@     �X@      0@       @      �?      @      �?      �?      @                                                                                       @      �?      $@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJɇ}hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?i���C�@�	           ��@       	                    @����@$           ��@                          �5@�ɛW/�@3           ��@                          �3@�U� @�           ��@������������������������       ��t�0@V           p�@������������������������       �"զmsp@�            �l@                           �?���u�@I           ��@������������������������       ��F�4�d@            �i@������������������������       �[�ɚe�@�            pt@
                           @���K~@�            �w@                          �6@��L�# @�             n@������������������������       �5d�Fy@S            `a@������������������������       �Q݈%`@A            @Y@                          �6@��ݭU
@]            `a@������������������������       ��k���@B            �W@������������������������       ��g��@             F@                          �6@��ȁ@�           J�@                           �?�5N��Y@@           0�@                          �3@x:,'y�@T           (�@������������������������       �$���@�            �p@������������������������       �)�ܮ��@�             o@                            �?�,�w��@�           8�@������������������������       �G�s�n
@�            `o@������������������������       ���X�J[@X           `�@                          @A@��zs@S           Ȍ@                          �9@�!l E^@A           �@������������������������       ��nO�o@           @|@������������������������       ��j����@#           �{@                            @j�ޔ:6	@             <@������������������������       �����@             0@������������������������       ��[���@             (@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       pt@      `@      ]@     �s@      =@      }@      @      m@      6@     �}@     �\@      N@      ?@      T@     @l@     @Q@      w@     0r@      ~@     @S@     �a@     �A@      E@      a@      ,@     �m@      @      X@      @      n@      I@      3@      0@      7@     �X@      .@     �c@     �_@      j@      B@      Y@      6@      @@     �Z@      &@     �g@      @     �T@       @     �g@      C@      1@      .@      2@     �Q@       @     �]@     �T@     @f@     �@@     �M@      &@      $@      R@       @     ``@             �E@              [@      *@       @      *@      @     �C@      �?     �Q@      H@     �`@      3@      A@      @      $@      H@              X@             �@@             @V@      @      @       @      @      ?@              L@      A@      W@      $@      9@      @              8@       @     �A@              $@              3@      @      �?      &@      �?       @      �?      .@      ,@     �E@      "@     �D@      &@      6@     �A@      "@      M@      @      D@       @     �T@      9@      "@       @      (@      @@      @      H@     �A@     �E@      ,@      $@      @      $@      "@      @      4@      @      3@      �?      3@      .@      @              @      *@      �?      6@      3@      1@       @      ?@      @      (@      :@      @      C@              5@      �?     �O@      $@      @       @      @      3@      @      :@      0@      :@      (@      E@      *@      $@      =@      @     �G@              *@       @      I@      (@       @      �?      @      <@      @      C@      F@      >@      @      =@      $@      "@      7@       @      0@              "@       @      D@      @      �?      �?      @      2@      @      3@      4@      4@       @      .@       @      @      ,@              0@              @              3@      @      �?                      @      @      $@      3@      $@              ,@       @      @      "@       @                      @       @      5@      �?              �?      @      &@      @      "@      �?      $@       @      *@      @      �?      @      �?      ?@              @              $@      @      �?                      $@              3@      8@      $@      �?      @       @      �?      @              =@              @              @       @      �?                      @              2@      "@      "@      �?      $@      �?              @      �?       @                              @      @                              @              �?      .@      �?              g@     @W@     �R@     �f@      .@     �l@      �?      a@      2@      m@      P@     �D@      .@     �L@     �_@      K@     `j@     �d@      q@     �D@      X@      E@      >@     �[@      *@      d@              R@      ,@     �c@      C@      9@      @      4@      R@      7@     ``@     @U@     �e@      6@     �C@      ;@      1@      J@      &@     �K@              =@      $@      O@      0@      (@      @      0@      6@       @     �D@      D@     �E@      (@      2@      @      (@      @@      @      :@              ,@      @      =@      @      @              @      .@      @      1@      @@      >@      @      5@      4@      @      4@      @      =@              .@      @     �@@      "@      @      @      $@      @      @      8@       @      *@      @     �L@      .@      *@     �M@       @     @Z@             �E@      @     �W@      6@      *@       @      @      I@      .@     �V@     �F@     ``@      $@      $@      @      @      :@             �B@              @      �?      <@      @      @               @      @      @      <@      0@     �P@       @     �G@      $@      @     �@@       @      Q@             �B@      @     �P@      3@      "@       @       @      F@      (@      O@      =@      P@       @     @V@     �I@      F@     �Q@       @      Q@      �?     @P@      @      S@      :@      0@       @     �B@     �K@      ?@      T@     �S@      Y@      3@      U@     �E@     �E@     �P@       @      Q@      �?     @P@      @     �R@      8@      .@      @      B@      K@      ?@     �S@     �S@     �X@      3@      J@      9@      4@      C@       @      @@      �?      3@      @      G@      *@      @      @      5@      4@      0@     �E@      C@     �D@      (@      @@      2@      7@      =@              B@              G@      �?      =@      &@       @      @      .@      A@      .@      B@     �D@     �L@      @      @       @      �?      @                                              �?       @      �?       @      �?      �?              �?               @              @      @                                                                              �?       @              �?              �?               @               @       @      �?      @                                              �?       @                      �?                                                �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJj��hhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�T5���@�	           ��@       	                   �3@@
�^@�           ��@                            @8�y��w@           �@                          �1@1m�@�           d�@������������������������       �ޡ�Կ~
@@           p�@������������������������       �!��o]�@S           X�@                          �2@�7��\}@�            �v@������������������������       ���K�@�             q@������������������������       ��jXx��
@?            �W@
                           �?=z5�3@c           ��@                           �?�sd'7@�            �w@������������������������       ��E/��@T            �a@������������������������       ���#8�:@�            @n@                           �?b�O���@l           ��@������������������������       ��}���@�             r@������������������������       ��5�#@�            s@                          �7@�����@�           ė@                           @�N�u�@�            0r@                           �?4�Y�F@�            �o@������������������������       �6u[��I
@;             Z@������������������������       ����E[�@\            �b@                           @;��I
�	@             B@������������������������       �RM棿@	             ,@������������������������       ��
�)�@             6@                          �<@q�q��@           8�@                           @T��@6           x�@������������������������       ��w���@�            �x@������������������������       �Ur�5�]@=           �@                            �?��n@�            �s@������������������������       ��Il.@@             X@������������������������       ��-���P@�            �k@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �s@      b@     @V@      w@      A@     �}@      @      o@      <@     �|@     �Y@     @Q@     �A@      L@     �k@     �P@     �v@     �q@     p|@     �U@     `e@      J@     �C@     @l@      .@     �w@       @     �a@      $@     `s@     �J@     �D@      *@      4@     �a@      ?@     `n@     `d@     �r@      I@     �S@      4@      6@      a@       @      l@      �?      U@      @     @i@     �@@      .@      @       @     @V@      4@     `a@      V@      k@      7@     �H@      *@      (@     �Z@      �?     �d@             �N@      @     �b@      0@      ,@      @      @     �P@      .@     �Z@     �P@     `f@      *@      5@      @      "@     �G@      �?     �U@              =@             �U@      @       @      �?              D@      @     �H@     �E@     @W@      @      <@      $@      @      N@              T@              @@      @      P@      "@      (@       @      @      ;@      &@     �L@      7@     �U@      $@      =@      @      $@      >@      @     �L@      �?      7@             �I@      1@      �?              @      6@      @     �@@      6@      C@      $@      7@      @      �?      8@      @      B@      �?      2@             �F@      @      �?              �?      1@      @      =@      0@      :@      $@      @              "@      @              5@              @              @      (@                       @      @              @      @      (@             @W@      @@      1@     @V@      @      c@      �?      L@      @      [@      4@      :@      $@      (@      J@      &@      Z@     �R@     �S@      ;@      F@      1@      &@      B@      @     �B@      �?      A@      @     �G@      @      (@      @      @      2@      @      A@      <@      3@      $@      9@      @      @      @       @      .@      �?      7@              "@      �?      @              �?      @      �?      ,@      &@      &@      �?      3@      *@       @      ?@      @      6@              &@      @      C@      @      @      @      @      (@      @      4@      1@       @      "@     �H@      .@      @     �J@      �?     �\@              6@             �N@      .@      ,@      @      @      A@      @     �Q@     �G@      N@      1@      9@      "@      @      7@             �H@              $@              A@      (@      @      @      @      2@       @      6@      <@     �A@      "@      8@      @      @      >@      �?     �P@              (@              ;@      @      "@      @       @      0@      @      H@      3@      9@       @     @b@      W@      I@      b@      3@     �Y@      @     @[@      2@     �b@     �H@      <@      6@      B@     �S@     �A@     �]@     �^@     �c@      B@     �F@      @      @      D@      �?      0@              $@      @      9@      @       @      �?      @      3@      &@     �@@     �@@      4@       @     �E@      @      �?      B@      �?      (@              $@      @      4@      @       @      �?      @      .@      "@      ?@      :@      4@       @      8@      @              0@      �?      @               @      @      $@       @                              @              $@      0@      @       @      3@      @      �?      4@              @               @      �?      $@      @       @      �?      @      &@      "@      5@      $@      .@      @       @              @      @              @                              @                               @      @       @       @      @                       @              @      �?                                                                                      �?               @      @                                              @              @                              @                               @      @       @              @                     @Y@     @U@     �F@      Z@      2@     �U@      @     �X@      ,@     �_@     �E@      :@      5@      ?@      N@      8@     �U@     �V@     `a@      <@     @S@      K@      :@     �V@      $@     @P@      �?     @S@      $@      Z@      :@      5@      (@      6@      H@      2@     �P@     �K@     �Y@      :@      8@      *@      *@     �D@      @      :@      �?      E@      @     �G@      2@      *@                      2@      (@      B@      :@      G@      *@     �J@     �D@      *@      I@      @     �C@             �A@      @     �L@       @       @      (@      6@      >@      @      >@      =@      L@      *@      8@      ?@      3@      *@       @      5@      @      6@      @      6@      1@      @      "@      "@      (@      @      4@     �A@     �B@       @       @      @      @      �?              $@              $@      @       @       @              @      @      @       @      @      0@      @      �?      6@      8@      ,@      (@       @      &@      @      (@              ,@      .@      @      @      @      @      @      .@      3@      ?@      �?�t�bub��     hhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ#֤hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?A(/�@�	           ��@       	                    �?ٟ��@           ,�@                          �;@	Ľ'{@c            �@                            �?�]��A@<           (�@������������������������       ��kP��@f            �b@������������������������       �d6��a@�            �v@                           �?Kz�)�@'            �O@������������������������       �P,�h��	@             <@������������������������       �~hۻ�
@            �A@
                           �?��d�e@�           �@                            @vy���@�            �u@������������������������       �\F���@t            �f@������������������������       ���M�@e            @d@                          �1@gg�f'@�           p�@������������������������       ��7�$k
@,            �R@������������������������       ��ԧ�5@�           �@                           �?�}�3@�           |�@                          �9@��;��@            X�@                          �1@�O~�t@�           x�@������������������������       ��O_	{�@p            �e@������������������������       ��`�+\�@n            �@                           @�X��U@B             W@������������������������       �h#���@3            �Q@������������������������       ��|K��@             5@                          �6@z�P���@v           ̕@                          �2@�V�3��@V            �@������������������������       �R�`�Խ@           @}@������������������������       ��{!)w@;            @                           �?p*���@            �z@������������������������       ����@             h@������������������������       ��R�H#�@�            �m@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       @t@     �_@     �W@     pt@     �B@     `~@      @     @k@      =@     p}@     �W@     �L@      D@      T@     �n@     �K@     �w@      t@     �{@     @T@     @`@     �R@      P@     `b@      ;@     @c@      @     @\@      6@     �b@      @@     �@@      7@     �M@      Z@      >@     �b@     �a@     @g@     �B@     �D@      .@      9@      K@             �R@       @      5@       @     �J@      &@      &@      @      .@      C@      (@      K@     �F@     @U@      "@      D@      "@      9@      J@             @Q@       @      1@      @     �D@      "@      &@       @      &@      B@      &@     �H@      D@     �S@      "@       @      �?      @      5@              9@              @       @      $@      @      �?       @      �?       @       @      &@      $@      @@      @      @@       @      5@      ?@              F@       @      &@      @      ?@      @      $@              $@      <@      "@      C@      >@      G@      @      �?      @               @              @              @       @      (@       @              @      @       @      �?      @      @      @                       @                               @              @       @       @      �?               @      @      �?      �?      �?              �?              �?      @               @              @              �?              @      �?              @              �?              @      @      @             @V@     �M@     �C@     @W@      ;@      T@      �?      W@      ,@     �W@      5@      6@      0@      F@     �P@      2@     �W@     �W@     @Y@      <@      7@      5@      1@      9@      @      7@              A@      �?     �E@      @      @      @      ,@      6@       @     �E@      4@     �@@      @      @      0@       @      2@       @      (@              &@              ?@      @      �?      @      @      *@      �?      7@      $@      ,@      @      0@      @      "@      @      @      &@              7@      �?      (@       @       @              "@      "@      �?      4@      $@      3@      @     �P@      C@      6@      Q@      6@     �L@      �?      M@      *@      J@      0@      3@      (@      >@      F@      0@      J@     �R@      Q@      5@      @      �?       @      &@              *@               @              @              @      @               @                      @      &@             �M@     �B@      4@     �L@      6@      F@      �?      I@      *@     �G@      0@      0@      @      >@      E@      0@      J@      Q@     �L@      5@     @h@      J@      ?@     �f@      $@     �t@      �?     @Z@      @     0t@     �O@      8@      1@      5@     �a@      9@     �l@     �f@     @p@      F@      R@      *@      $@      L@      @     �b@              @@              `@      6@      "@      @      @      J@      @      T@      P@      ]@      7@     @P@      (@      $@      J@      �?     �`@              >@              ]@      4@      @              @     �G@      �?      R@      M@      [@      .@       @                      @      �?     �G@               @             �@@              @                      "@      �?      .@      $@      =@      @     �L@      (@      $@     �G@             �U@              6@             �T@      4@       @              @      C@             �L@      H@     �S@      $@      @      �?              @      @      .@               @              (@       @      @      @      �?      @      @       @      @       @       @       @                      @      @      ,@               @              @               @      @      �?      @      @      @      @      @       @      @      �?                              �?                              @       @      �?                       @              �?      �?       @             �^@     �C@      5@      _@      @     �f@      �?     @R@      @     `h@     �D@      .@      ,@      0@      V@      4@     �b@      ]@      b@      5@      P@      :@      0@     @W@      �?     �a@             �K@       @     �b@      8@      (@      &@      @     �K@      $@     �Z@     �S@     @Y@      &@      B@      "@       @      H@              M@              A@             �V@      "@       @      @       @      7@      @     �J@     �@@     �I@      @      <@      1@      ,@     �F@      �?     �T@              5@       @      N@      .@      $@      @      @      @@      @     �J@     �F@      I@      @      M@      *@      @      ?@      @      E@      �?      2@      @      F@      1@      @      @      "@     �@@      $@     �E@      C@     �E@      $@      B@      @              ,@       @      8@      �?       @      @      0@      @                              3@      @      .@      .@      .@      @      6@      @      @      1@      @      2@              $@              <@      (@      @      @      "@      ,@      @      <@      7@      <@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��bhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�۝�ٳ@�	           ��@       	                   �4@B�-@�           �@                           @7nW�v�@D           �@                           �?�M9�@[           Ё@������������������������       ��3���@�            �v@������������������������       ���;�@�             j@                           @���So7@�           8�@������������������������       ��p��m	@�            px@������������������������       ��wo�N2@�             x@
                           �?«ܛ�'@�           ��@                          �;@�V]H�Q@A            @������������������������       �\*BD�@�            �x@������������������������       �5�TT�@B             Y@                           �?�t(��6@r           @�@������������������������       �)hٛ%�@�            @x@������������������������       ����#�@u            �@                           �?�h�:�@�           @�@                          �?@��i@�           ��@                           �?���9P�@�           ��@������������������������       ��F)Y��@�            �j@������������������������       �;���-@            z@                           �?���8�@             �M@������������������������       ��x�2�@
             4@������������������������       �����%	@            �C@                           @���`�@
            z@                          �1@"� r@�            ps@������������������������       ������8@#             J@������������������������       �\f(��k@�            0p@                           �?��9c@F            @Z@������������������������       ��l����	@"            �J@������������������������       ��Gq���@$             J@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       Pt@      a@     @Y@     �v@     �G@     0|@      @     �p@      A@     �z@     �Z@     �P@     �A@     @R@      j@      L@     �u@     �s@     �}@      Q@     �l@      Y@      J@      r@      8@     0u@       @     �e@      6@     Pu@     �P@      F@      4@      H@      c@      D@      o@     �i@     �v@      G@     �S@      @@      2@     �c@       @      g@             �V@       @     @g@      :@      ,@      @       @     �R@      *@     �Y@     @\@      j@      7@      C@      (@      *@      U@       @     �L@              A@      @     @P@      1@      "@      �?      @      >@      $@      B@      K@      T@      1@      <@      (@      &@     �G@       @     �B@              6@      @     �D@      &@       @      �?      @      4@       @      *@     �@@      J@      *@      $@               @     �B@              4@              (@              8@      @      �?               @      $@       @      7@      5@      <@      @     �D@      4@      @     �R@              `@              L@      @     @^@      "@      @      @      �?      F@      @     �P@     �M@      `@      @      $@      $@       @     �F@             �S@              6@             �Q@      �?      @              �?      5@       @      <@      8@     �Q@      �?      ?@      $@      @      >@              I@              A@      @      I@       @      �?      @              7@      �?      C@     �A@     �L@      @     �b@      Q@      A@     ``@      6@     @c@       @     @U@      ,@     `c@     �D@      >@      .@      D@     �S@      ;@     `b@     �V@     �c@      7@      F@      ,@      1@      >@      @     @Q@      �?      ;@              J@      .@       @      @      &@      8@      @     �L@      @@      P@      .@      C@      "@      $@      :@      @     �K@      �?      7@              C@      "@      �?              $@      4@       @     �J@      ;@      L@      .@      @      @      @      @       @      ,@              @              ,@      @      @      @      �?      @       @      @      @       @             @Z@      K@      1@     @Y@      1@     @U@      �?      M@      ,@     �Y@      :@      6@       @      =@     �K@      7@     �V@     �M@     @W@       @     �G@      "@      @      E@      "@      C@      �?      5@       @     �E@      ,@      @      @      @      8@      ,@     �G@      9@      8@      �?      M@     �F@      (@     �M@       @     �G@             �B@      @      N@      (@      0@      @      6@      ?@      "@     �E@      A@     @Q@      @     @X@     �B@     �H@     @S@      7@      \@      �?     @V@      (@     @V@      D@      7@      .@      9@      L@      0@     @Y@      [@      \@      6@     �M@      7@     �B@      C@      5@     �O@      �?     �N@      (@     �@@      9@      4@      *@      6@     �A@       @     @P@     �R@     �P@      (@      I@      .@      ?@     �A@      3@     �N@      �?      N@      (@      @@      7@      4@      @      3@     �A@       @      O@      P@     @P@      &@      9@      @      &@      $@       @      5@              4@      @      $@       @      @      �?      @       @       @      7@      8@      6@       @      9@      &@      4@      9@      &@      D@      �?      D@      "@      6@      .@      .@      @      *@      ;@      @     �C@      D@     �E@      "@      "@       @      @      @       @       @              �?              �?       @              @      @                      @      $@      �?      �?              @                                              �?                       @              @                              �?       @      �?              "@      �?      @      @       @       @                              �?                      �?      @                       @       @              �?      C@      ,@      (@     �C@       @     �H@              <@              L@      .@      @       @      @      5@       @      B@      A@      G@      $@      >@      (@      &@      =@       @      F@              2@             �C@      *@                              *@       @      <@      6@      B@      @      @      �?       @      @              ,@               @              (@       @                                              @      �?      �?              7@      &@      "@      9@       @      >@              0@              ;@      &@                              *@       @      6@      5@     �A@      @       @       @      �?      $@              @              $@              1@       @      @       @      @       @               @      (@      $@      @      @                      @              @              @              @              �?                      @               @      "@      $@      @      @       @      �?      @              �?              @              $@       @       @       @      @      @              @      @              �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�#�$hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@ʂڵ��@�	           ��@       	                    �?����x�@b           x�@                          �2@ `w�ev@W           ��@                            @1Bq��?@
           �z@������������������������       ��]F��	@�            `s@������������������������       ��/��@D            @^@                           �?Q�J*H
@M            ``@������������������������       �	��:�@            �H@������������������������       ��B���B@.            �T@
                            �?�{�r�@           `�@                          �2@M�O
@�            `n@������������������������       ��/��	@w            @g@������������������������       ���j�V=@%            �L@                           �?�ø@o           ȁ@������������������������       ���z8�@            �G@������������������������       ��EC�@X           P�@                           �?h��5e@?           ֣@                          �:@���#@	           h�@                           @����	@(           P�@������������������������       ��Sd@�           ��@������������������������       �1���@�             o@                            �?�s �@�             w@������������������������       �V�@t             h@������������������������       ��h�aHd@m            �e@                            �?iT��]$@6           D�@                          �;@���Ө�@�            �w@������������������������       ���R&`@�            �t@������������������������       � A��ɗ
@            �E@                           @�A�)@M           ��@������������������������       �i]���@X           ��@������������������������       �B�0F.@�             x@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        x@     �_@     �W@     �u@     �A@      ~@      "@     �k@      :@      |@     @Z@      Q@      D@      M@      i@     �O@     pv@     pt@      z@     �X@      ^@      9@      4@     @b@      @      k@      �?     @R@       @     �f@      ;@      7@       @      (@     �S@      ,@      \@      Z@     �g@      5@     @P@       @      "@     �I@      @      W@             �C@      �?     �S@      (@      @      �?      @      >@       @     �C@      ?@      W@      @     �G@      �?       @      >@      @     �S@              @@      �?      L@      @      �?      �?      @      4@       @     �@@      =@     @R@      @      :@      �?      @      :@       @     �N@              .@      �?     �G@      �?      �?              �?      3@              8@      6@     �L@      @      5@              @      @      �?      2@              1@              "@      @              �?       @      �?       @      "@      @      0@       @      2@      �?      �?      5@              *@              @              7@      @      @                      $@              @       @      3@              @      �?      �?      �?              @              @              *@      @      @                       @                              (@              ,@                      4@              "@              @              $@       @                               @              @       @      @             �K@      7@      &@     �W@      @     @_@      �?      A@      �?     �Y@      .@      1@      �?      "@      H@      (@     @R@     @R@     @X@      0@      .@      @              A@             �B@              @              B@      @      @                      (@              8@      ,@      F@      $@      ,@      �?             �@@              ?@              @              @@      @      @                      @              0@      &@      ;@      @      �?      @              �?              @               @              @                                      @               @      @      1@      @      D@      3@      &@     �N@      @      V@      �?      <@      �?     �P@      &@      ,@      �?      "@      B@      (@     �H@     �M@     �J@      @      �?      @              @              1@                               @                              �?                              $@                     �C@      .@      &@     �K@      @     �Q@      �?      <@      �?      M@      &@      ,@      �?       @      B@      (@     �H@     �H@     �J@      @     �p@     @Y@     �R@     �i@      <@     �p@       @     `b@      8@     �p@     �S@     �F@      C@      G@     �^@     �H@     �n@     �k@     �l@     @S@     �Z@      K@      K@     �X@      1@     �X@      @     �V@      0@     @\@      D@      A@      8@      A@      M@      9@     @]@     �[@     �Z@      C@     �T@     �@@      A@      O@      ,@     �V@      @      M@      ,@     @T@      ?@      :@      "@      :@      F@      ,@      V@     �Q@     �O@      >@     �O@      5@      5@      J@      @     �R@      @     �H@       @      H@      >@      *@      @      .@      =@      @      O@     �I@     �H@      8@      4@      (@      *@      $@       @      1@              "@      @     �@@      �?      *@      @      &@      .@      "@      :@      3@      ,@      @      7@      5@      4@     �B@      @       @      @     �@@       @      @@      "@       @      .@       @      ,@      &@      =@      D@      F@       @      @      $@      @      2@               @       @      9@      �?      2@      @      @      (@      @      @      @      *@      4@      7@       @      0@      &@      *@      3@      @              �?       @      �?      ,@       @      @      @      @      &@      @      0@      4@      5@             �c@     �G@      5@     @Z@      &@     �d@       @      L@       @     �c@      C@      &@      ,@      (@      P@      8@     @`@     @\@     �^@     �C@     �F@      ,@      $@      C@      �?     �L@              .@              ?@      "@      @      @      @      :@       @      <@     �C@      A@      @      E@      ,@       @      C@              G@              ,@              ?@      @      @       @      @      8@      @      9@      A@      =@      @      @               @              �?      &@              �?                       @              @      �?       @       @      @      @      @             @\@     �@@      &@     �P@      $@     @[@       @     �D@       @     @_@      =@      @      @       @      C@      0@     �Y@     �R@      V@      @@     �Q@      4@      @      ?@       @      N@              2@       @     @V@      0@       @       @       @      8@      @     �M@      J@      K@      7@     �E@      *@       @      B@       @     �H@       @      7@      @      B@      *@      @      @      @      ,@      "@     �E@      6@      A@      "@�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��]hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���@�@�	           ��@       	                    �?�$��@�           `�@                            @B��_�~@X           P�@                           @lÍ@�            �t@������������������������       ��[{臧@�            `k@������������������������       �C#5���@E            @\@                          �:@�4.��:@�            �k@������������������������       �7hU�Pj@p            @f@������������������������       �?�nF$q@             F@
                          �1@�8�J#�@�           ��@                           �?�ys,��@>            @X@������������������������       �`��9�@             3@������������������������       �ֶ!�V�@/            �S@                          �@@V��Ô�@b           h�@������������������������       ��EIj�@O           @�@������������������������       �6����@            �B@                          �2@�4m�˓@�           �@                            @~yn��@�           8�@                          �1@����@�           X�@������������������������       �[�5��
@�            Px@������������������������       ����
@�            �l@                          �1@�v��l�@`            �c@������������������������       �e+�Y��
@7             U@������������������������       ���(ї@)             R@                          �9@��"�[:@�           ��@                           @/�G:�@�           ��@������������������������       �I�.%�=@�           �@������������������������       �X�`�{y@N           �@                           @(���2@�            @t@������������������������       ��s��@�            �m@������������������������       ��r|ԭ@9            �U@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       0u@     @a@     �W@     �v@     �@@     `}@      @      k@      C@     �{@      \@      N@     �B@     �R@     `l@      T@     Pv@     �s@     p{@     @R@     �a@     �N@     �O@      e@      ;@     �a@      @     �Y@      9@     ``@      I@     �@@      3@      D@      V@      G@      b@      a@     �d@     �B@      L@      &@      :@     �I@      *@     �M@      @     �F@      @     �B@      *@      @      @      ,@      >@      0@      H@      G@     �L@      (@      3@       @      ,@      8@      "@     �B@       @      A@       @      :@       @      @       @      @      0@      *@      =@      8@      E@      &@      @      @      "@      *@      @      A@       @      :@       @      3@      @      @       @      �?      @      @      4@      .@      <@      @      ,@      @      @      &@       @      @               @              @      �?      �?              @      "@      @      "@      "@      ,@      @     �B@      @      (@      ;@      @      6@      �?      &@      @      &@      @      �?       @      @      ,@      @      3@      6@      .@      �?      =@       @      "@      5@       @      6@              @      @      $@      @      �?              @      ,@      @      3@      0@      "@      �?       @      �?      @      @       @              �?      @       @      �?      �?               @      �?                              @      @              U@      I@     �B@     �]@      ,@     �T@       @     �L@      2@     �W@     �B@      ;@      .@      :@      M@      >@     @X@     �V@     �Z@      9@      @               @       @      @      (@       @      @       @      @      �?      @                      (@       @      @       @      .@                               @      @                                       @      �?                                      �?      �?               @      @              @              @      @      @      (@       @      @              @      �?      @                      &@      �?      @      @      $@             �S@      I@      =@     �[@      $@     �Q@              J@      0@      V@      B@      7@      .@      :@      G@      <@     �W@     �T@      W@      9@     �S@      E@      8@     �Z@      $@     �Q@              J@      0@      T@     �A@      3@      ,@      9@      G@      <@      W@     �S@      W@      9@               @      @      @                                               @      �?      @      �?      �?                       @      @                     �h@     @S@      @@     @h@      @     �t@             �\@      *@     `s@      O@      ;@      2@     �A@     `a@      A@     �j@      f@     0q@      B@      L@      .@      "@     @Q@             �^@              G@             ``@      $@      $@      @      @      G@       @     �O@     �F@     �_@      @      @@      ,@      @      K@             @W@             �@@             �[@      @       @      @      @     �C@      @     �I@     �C@     @]@      @      5@      @      @      :@              Q@              0@              P@      @      @      �?      �?     �@@      @      ;@      @@     @R@      @      &@      @       @      <@              9@              1@              G@      @      @      @       @      @              8@      @      F@              8@      �?       @      .@              =@              *@              5@      @       @              @      @      @      (@      @      $@       @      "@      �?       @      @              7@              @              "@       @       @              @      @              (@      @      �?       @      .@                      $@              @              @              (@      �?                              @      @              @      "@             �a@      O@      7@     @_@      @     �i@             @Q@      *@     `f@      J@      1@      ,@      <@     @W@      :@     �b@     �`@     �b@      =@     �\@     �K@      1@     �Z@       @     �d@             �F@      &@     �b@      C@      $@       @      0@     �P@      2@      ]@     @]@      \@      6@      P@      C@      "@      L@       @     @V@              <@       @      V@      3@       @       @      @      @@      2@     �P@      N@     �M@      .@     �I@      1@       @      I@             �S@              1@      @     �N@      3@       @              "@      A@             �H@     �L@     �J@      @      <@      @      @      3@      @     �C@              8@       @      >@      ,@      @      @      (@      ;@       @     �@@      .@      B@      @      ,@      @      @      &@       @      C@              $@       @      ;@      *@      @      @      &@      9@      @      3@       @      ;@      @      ,@      �?      @       @       @      �?              ,@              @      �?                      �?       @      @      ,@      @      "@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ!��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@#��]P�@�	           ��@       	                    �?���b�@           ��@                          �5@�os:S�@$            �@                            �?^X:<@�           ��@������������������������       �CUB0@�            `n@������������������������       �~����@C           �@                            @�D�=@L            �[@������������������������       �!��^Y	@'             N@������������������������       �6+�l�<@%            �I@
                            �?�	��E�@�           l�@                           �?��/Ś�@A           ��@������������������������       �I~� �,@�            �t@������������������������       ��7dW	I@r           P�@                            @�����@�           @�@������������������������       �_�����
@�            �u@������������������������       ������@�            �r@                           �?��p^�@�           8�@                           @�B^��O@w           p�@                          �9@.��?5N@K           0�@������������������������       ��0�*]@�            @q@������������������������       �-�(v
@�            @n@                            �?�;V�@,             R@������������������������       �s��R��@            �I@������������������������       �Lfb!:�@             5@                          �;@��ذ#�@6            �@                           @��S���@�           ��@������������������������       �1R�S�l@a           x�@������������������������       �
R?N�@'            @P@                          �<@k����@�             q@������������������������       ���g>D@+             O@������������������������       �P�m�{�@�            @j@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@      a@     �W@     0u@     �H@     �}@      @     �o@      >@      }@     @W@     �L@      G@     @Q@     �j@      R@     �v@     �r@      |@     @S@     �g@     �P@     �M@     �j@      :@     �v@             `c@      *@     �t@     �H@     �C@      *@      8@     @_@     �A@      o@     @c@     0r@      B@     �U@      8@      <@     �S@      4@     �X@             �O@       @     �U@      5@      0@       @      1@      H@      $@     �S@     �L@     �Y@      2@     @U@      ,@      9@     �Q@      1@     �S@             �J@       @      R@      1@      .@      �?      (@      G@       @     @Q@     �K@     �V@      1@      .@       @      @     �@@       @      2@              6@      @      @@      @      @      �?      @      6@      @      1@      (@      >@      &@     �Q@      (@      3@     �B@      .@     �N@              ?@      @      D@      ,@      $@               @      8@      @      J@     �E@      N@      @       @      $@      @      "@      @      4@              $@              ,@      @      �?      �?      @       @       @      "@       @      *@      �?      �?              �?      @              *@              @              @                      �?      @      �?       @      @              (@      �?      �?      $@       @      @      @      @              @              @      @      �?               @      �?               @       @      �?             @Y@      E@      ?@     �`@      @     �p@              W@      @     `n@      <@      7@      &@      @     @S@      9@     @e@     @X@     �g@      2@      L@      =@      2@     @S@       @     `a@             �E@      @      a@      5@      .@      &@       @      E@      (@     @X@     @Q@      `@      *@      1@      @      @     �A@      �?     �M@              :@      �?      J@      @                              2@       @     �A@      5@     �D@      @     �C@      8@      *@      E@      �?      T@              1@       @     @U@      .@      .@      &@       @      8@      $@      O@      H@      V@       @     �F@      *@      *@      M@      @     @_@             �H@       @     �Z@      @       @              @     �A@      *@     @R@      <@     �M@      @      3@      @      @      =@      �?     �S@              9@       @      L@      @       @              @      6@             �F@      ,@      A@      �?      :@      "@      @      =@      @     �G@              8@              I@      @                       @      *@      *@      <@      ,@      9@      @      b@     �Q@     �A@     @_@      7@     �[@      @     @X@      1@      a@      F@      2@     �@@     �F@     �U@     �B@     �\@     �a@     �c@     �D@      R@      0@      0@     �I@       @     �D@      @      D@      *@      N@      3@       @      "@      @      C@      0@      I@      M@     �K@      .@     @P@      $@      &@      I@       @      @@      @      C@      *@     �H@      .@       @      "@      @     �B@      0@     �D@      J@     �F@      .@      D@      @      @      <@      �?      4@              4@       @     �B@       @      �?              @      8@      @      6@      ?@      ,@      @      9@      @      @      6@      @      (@      @      2@      @      (@      @      �?      "@      @      *@      &@      3@      5@      ?@      &@      @      @      @      �?              "@      �?       @              &@      @                              �?              "@      @      $@              @      @      @                      "@               @              "@      @                                              "@               @                       @              �?                      �?                       @                                      �?                      @       @             @R@     �K@      3@     �R@      .@     @Q@       @     �L@      @     @S@      9@      0@      8@      C@     �H@      5@      P@      U@      Z@      :@     �G@      ;@      (@      H@      @      N@       @     �D@      @      O@      5@      $@      ,@      <@     �A@      3@     �J@     �I@     �P@      2@      F@      2@      (@      H@      @      K@       @      C@      @     �L@      3@       @       @      :@     �@@      $@     �G@     �E@     �P@      2@      @      "@                       @      @              @              @       @       @      @       @       @      "@      @       @                      :@      <@      @      :@      "@      "@              0@              .@      @      @      $@      $@      ,@       @      &@     �@@      C@       @      �?       @              @                              @              @      �?      @              @       @              �?      @      &@      @      9@      4@      @      4@      "@      "@              "@              "@      @       @      $@      @      (@       @      $@      ;@      ;@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�wwhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @&r�xA�@�	           ��@       	                    �?eW\�Դ@           ��@                            �?^��W�@&           l�@                           �?�ܮ9�@N           �@������������������������       �+�K�B�@h            �f@������������������������       �(F��"?@�            �v@                          �?@w�<�+�@�           ��@������������������������       �.�i�@�           ܐ@������������������������       ���J5��@,            �Q@
                          �7@��ÎV�@Y           ��@                            �?���\�@�            @x@������������������������       ���� [@E             ^@������������������������       �]��u��@�            �p@                            �?��,�@u             g@������������������������       ��1�k@H            �[@������������������������       ��K'*@-            @R@                          �6@��BY�@           ș@                           @�,j0�@�           �@                           @'�r�o@�           ��@������������������������       ��Ti�9
@_           8�@������������������������       �o�T�>@�            �m@                           @RO%@�            w@������������������������       ���P�@@            @X@������������������������       ��ųLڇ@�             q@                          �:@�˸�o�@3           �~@                          �9@D�J�<Q@�             s@������������������������       ��5��@�             p@������������������������       �CJ�(i�
@!             I@                           �?�64hG�@l            @g@������������������������       ���bs
@1            �U@������������������������       ����[�@;             Y@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        u@     �a@     @V@     �u@     �D@     �z@      "@     @m@      7@     �}@     �[@     �Q@      C@     @Q@     �l@      N@     `y@     @t@     �y@      S@      g@     �V@     �Q@     `j@      @@     �g@      "@      c@      .@     �n@      T@      J@     �@@      J@      `@      G@     @j@     �h@     @j@     �K@     �`@      Q@     �O@     �d@      <@      _@      "@     �_@      (@     �e@     �M@     �C@      6@      F@     �W@      >@      c@     @b@      d@     �E@     �@@      >@      ,@      O@      (@      H@      @      J@       @      I@       @       @      @      ,@      B@      @      B@     �F@     �P@       @      .@       @      @      6@      �?      3@              2@              ;@      @       @      @       @      (@              "@      0@      4@              2@      <@       @      D@      &@      =@      @      A@       @      7@       @      @      @      (@      8@      @      ;@      =@     �G@       @     �X@      C@     �H@     �Y@      0@      S@      @     �R@      $@     �^@     �I@      ?@      .@      >@     �M@      :@      ]@     @Y@     �W@     �A@     @W@      <@     �D@     @X@      0@     �R@      @     @R@      $@     �]@     �H@      <@      (@      ;@     �M@      9@     @[@     @V@      W@      A@      @      $@       @      @              �?              �?              @       @      @      @      @              �?      @      (@       @      �?      J@      7@      @      G@      @     �P@              :@      @      R@      5@      *@      &@       @     �@@      0@      M@     �I@     �H@      (@      ;@      ,@      @     �@@             �E@              *@      �?      I@      ,@      (@      @      @      0@      $@     �J@     �F@      @@      @      @      �?      @      &@              @              @              2@              "@      @      @      @       @      *@      3@      "@      @      7@      *@       @      6@              B@              $@      �?      @@      ,@      @      @       @      $@       @      D@      :@      7@              9@      "@              *@      @      8@              *@       @      6@      @      �?      @      �?      1@      @      @      @      1@      @      1@      @              @      @      .@              @       @      *@      @              �?              &@      @      @      @      0@               @       @               @              "@               @              "@      @      �?      @      �?      @      @      �?       @      �?      @     @c@     �H@      3@     �`@      "@     `m@             �T@       @      m@      >@      3@      @      1@     @Y@      ,@     �h@     �_@     �h@      5@     �U@      @@      *@      W@      @     �g@             �Q@       @     �e@      3@      0@       @      �?      O@      "@     �`@      V@     �b@      $@     �O@      (@       @     �I@      @     �^@             �N@      �?      a@      0@      @      �?      �?     �F@       @     �W@     �I@     @Z@      "@     �@@       @      @     �@@      @     @Z@              B@              X@      @      @                      8@       @     @S@      B@      T@      @      >@      $@      �?      2@              1@              9@      �?      D@      &@      �?      �?      �?      5@              2@      .@      9@      @      8@      4@      @     �D@       @     @Q@              $@      �?     �B@      @      &@      �?              1@      @      C@     �B@     �F@      �?      @      $@      �?      @              "@              @              3@      �?      @                       @      @      &@      &@      *@      �?      4@      $@      @      B@       @      N@              @      �?      2@       @      @      �?              .@      @      ;@      :@      @@             �P@      1@      @     �D@       @      F@              &@      @     �M@      &@      @      @      0@     �C@      @     �O@     �C@     �H@      &@     �L@      (@       @      =@              >@              @      �?     �B@      @               @      @      <@      @      :@      8@      <@      &@      G@      &@       @      9@              <@              @      �?      A@      @                      @      8@      �?      7@      7@      4@      @      &@      �?              @               @               @              @                       @              @       @      @      �?       @      @      $@      @      @      (@       @      ,@              @      @      6@      @      @      �?      $@      &@       @     �B@      .@      5@              �?      �?       @      @       @      @              @      @      (@       @                      @      @       @      3@      *@      @              "@      @       @       @               @              �?              $@      @      @      �?      @      @              2@       @      2@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�̇BhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                              @��� �@�	           ��@       	                    �?�&��g@�           �@                          �7@�sa�X@d           Ў@                           �?.�|��5@z           Ђ@������������������������       ����v�Z@�             j@������������������������       �������@�            �x@                           @�{}���@�             x@������������������������       �$���@�            �u@������������������������       ��ϲ���
@            �B@
                          �3@Z��ɂ@�           ��@                          �0@V�h���
@�           Ȉ@������������������������       �;�:97@V            ``@������������������������       �>?�^@�           ��@                           �?�\Sш<@�           L�@������������������������       ����@;            @������������������������       ����7��@e           �@                           �?�Z��\@�           �@                           �?�*��$@&           �}@                          �1@{/��]�@g            @e@������������������������       �S�m�?�@             ?@������������������������       �;�[XF�@V            `a@                           �?�@*��@�            Ps@������������������������       ��7B���@c            �c@������������������������       ������	@\            �b@                           @�G��{�@�            �@                          �3@[�	��@k           0�@������������������������       �V��Q/@h            `c@������������������������       ��±6�@           �x@������������������������       ����j~�@'             O@�t�bh�h5h8K ��h:��R�(KKKK��h��B        �s@      a@      T@     �u@      H@     �~@      "@      l@     �B@     �|@     @X@     �G@     �I@      P@     �m@     �M@     v@     Pr@     �~@      R@     �i@      X@      G@     �o@      8@     �w@      "@      b@      2@     Pv@      M@      D@      B@      G@      f@      B@     �p@     @h@     `x@      I@      L@     �F@      ?@      X@      *@     @V@      @     �P@      (@     @\@      4@      5@      *@      7@     �N@      2@     �U@     �M@      a@      5@      B@      .@      ,@      M@       @      S@              C@      &@     �P@      @      *@      @      *@     �C@      $@     �J@      C@      W@      ,@      @      @      @      *@      �?     �B@              *@              1@              @      �?      @      0@              7@      (@      G@      @      =@      &@      "@     �F@      @     �C@              9@      &@      I@      @       @       @      "@      7@      $@      >@      :@      G@      $@      4@      >@      1@      C@      @      *@      @      <@      �?      G@      0@       @      $@      $@      6@       @     �@@      5@     �F@      @      3@      <@      ,@     �B@      @       @      @      :@      �?      F@      0@       @       @      @      6@       @      :@      2@      E@      @      �?       @      @      �?              @               @               @                       @      @                      @      @      @             �b@     �I@      .@     �c@      &@     �q@      @     �S@      @     �n@      C@      3@      7@      7@      ]@      2@     @f@     �`@     �o@      =@      E@      ,@      @      P@             �b@              D@      �?      ^@       @       @      @      @      I@      @     �S@      D@     �b@      "@      @      �?              "@             �D@              @              1@                                      $@      �?       @      @      @@             �B@      *@      @     �K@             �[@              B@      �?     �Y@       @       @      @      @      D@      @     �Q@     �B@     @]@      "@      [@     �B@      (@     �W@      &@      a@      @     �C@      @      _@      >@      &@      3@      3@     �P@      &@     �X@     �W@      Z@      4@     �N@      0@      @     �E@      @     @R@      @      &@      @     �I@      8@       @      &@      @      B@      @     �D@     �G@      E@      $@     �G@      5@       @     �I@      @     �O@              <@             @R@      @      "@       @      *@      >@       @      M@      H@      O@      $@      [@     �D@      A@     @W@      8@     �\@              T@      3@     @Z@     �C@      @      .@      2@     �M@      7@     @V@     �X@     �Y@      6@     �L@      &@      (@      G@      (@     �L@              ?@      "@      E@      1@      @      @      @      6@      @      6@      G@     �Q@      @      .@      �?      @      ,@       @      :@              .@      �?       @       @      �?       @      �?      ,@      �?      @      2@      5@      @      �?              �?              @      @                               @      @                              �?              @      @              �?      ,@      �?      @      ,@       @      3@              .@      �?      @       @      �?       @      �?      *@      �?      @      .@      5@      @      E@      $@      @      @@      @      ?@              0@       @      A@      "@       @       @      @       @      @      0@      <@     �H@       @      2@      @      @      &@      @      0@               @       @      "@      "@               @      @      @      @      @      &@      >@       @      8@      @              5@              .@               @              9@               @                      @      �?      "@      1@      3@             �I@      >@      6@     �G@      (@     �L@             �H@      $@     �O@      6@      @      &@      *@     �B@      1@     �P@     �J@      @@      .@     �F@      :@      5@     �D@      &@     �J@             �G@      $@     �M@      6@      @       @      *@      ;@      &@      N@     �G@      >@      .@       @      @      @      *@      @      3@              *@              :@      "@       @              @      @      �?      $@      1@      ,@             �B@      7@      .@      <@      @      A@              A@      $@     �@@      *@       @       @      $@      4@      $@      I@      >@      0@      .@      @      @      �?      @      �?      @               @              @                      @              $@      @      @      @       @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ- �yhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�@7���@�	           ��@       	                     �?���2@�           �@                           �?؎)6xl@H           �@                           �?h�G�@�           ��@������������������������       ���	���
@E             ]@������������������������       �y�x�@�           �@                           @3�׳��@~           ,�@������������������������       ��_�t��@           Ѓ@������������������������       �e�h��@�           ��@
                           �? ��M�@�           �@                          �:@��5fǕ@K             _@������������������������       ���
n�
@9             X@������������������������       �,�9	�@             <@                           �?�$���P@O           0�@������������������������       ����'@�            @m@������������������������       ��s�M�@�            �q@                          �6@����@�           �@                           �?5�%�{[@�           ��@                           �?����
@�            0r@������������������������       ���V��@[            �b@������������������������       �I��1@Z            �a@                          �1@�0����@�            Pu@������������������������       �.tFs��
@5             T@������������������������       ���Uvw�@�            Pp@                           �?�J4�^@)           �|@                          �9@�l���e@,            �P@������������������������       ����͵�	@             ?@������������������������       ��8�F�W@            �A@                          �?@U�>@3@�            �x@������������������������       ���8�$@�            �u@������������������������       �a�B��
@              H@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �r@     `a@     �V@     t@     �E@     p}@      *@     `k@      C@     �~@     @W@     �P@     �B@      Q@     @n@      J@     �v@     t@     |@     @X@      j@     @X@      L@      p@      8@     `v@      "@     �`@      6@     x@     �L@      E@      =@      D@     �f@      A@     0p@     �k@     �u@      N@     �e@     @V@     �I@      h@      2@     �l@      "@     �Z@      .@     �r@      J@      ?@      7@      ;@     �`@      <@     `h@     `e@      r@     �I@      M@      7@      1@     �T@      $@      X@             �F@      @     ``@      (@      @      @       @      J@      @     �N@     �@@     �Z@      $@      &@      �?      �?      0@              $@              @      @      &@      �?      @      �?              @       @       @      $@      >@             �G@      6@      0@     �P@      $@     �U@             �C@       @      ^@      &@      @      @       @     �F@       @     �M@      7@      S@      $@     �\@     �P@      A@     �[@       @     �`@      "@     �N@      $@     �d@      D@      8@      2@      9@     @T@      8@     �`@     @a@      g@     �D@      M@      =@      (@     �A@      �?     @R@      "@      ?@       @     �V@      1@      "@      "@      @      A@       @      L@      F@      T@      7@      L@     �B@      6@     �R@      @      N@              >@       @     �R@      7@      .@      "@      2@     �G@      0@     �S@     �W@      Z@      2@      B@       @      @      P@      @      `@              <@      @     @V@      @      &@      @      *@     �G@      @      P@      I@     �M@      "@      "@      @              1@      @      *@              @              ;@              �?              @      &@              @      "@      "@       @      "@      @              &@      @      *@              @              7@                              @      @              �?       @      @       @               @              @                              @              @              �?                      @              @      �?       @              ;@      @      @     �G@      @      ]@              5@      @      O@      @      $@      @      @      B@      @     �M@     �D@      I@      @      "@       @      �?      :@       @     �K@              "@      @      7@      @       @      @      @      $@      �?      0@      8@      >@       @      2@      �?      @      5@      �?     �N@              (@       @     �C@      �?       @       @      @      :@      @     �E@      1@      4@      @     �V@      E@      A@     @P@      3@     @\@      @     @U@      0@      [@      B@      9@       @      <@      O@      2@     �Y@      Y@      Y@     �B@     �M@      ;@      2@     �B@      $@     @V@      �?     �G@      @     @Q@      ,@      &@              $@      D@      &@     �P@      J@      L@      &@     �C@      @       @      9@      @      E@              5@              ;@      @      @              �?      .@       @      8@      <@      @@       @      =@      @      @      &@      @      2@              "@              @      @      @              �?      @              (@      3@      *@      @      $@      �?      �?      ,@              8@              (@              4@              �?                      $@       @      (@      "@      3@      @      4@      6@      $@      (@      @     �G@      �?      :@      @      E@      "@      @              "@      9@      "@     �E@      8@      8@      @      @      �?       @      �?              $@      �?       @              3@              @               @       @              @       @       @              ,@      5@       @      &@      @     �B@              2@      @      7@      "@      �?              @      1@      "@      B@      0@      6@      @      ?@      .@      0@      <@      "@      8@      @      C@      *@     �C@      6@      ,@       @      2@      6@      @      B@      H@      F@      :@      @      @      @       @       @      @      @       @       @      @      @      �?              �?       @              *@      @       @      �?                      @       @       @      @              �?      �?      �?      @      �?                                       @       @      �?              @      @                               @      @      @      �?       @       @                      �?       @              @       @      �?      �?      <@      (@      (@      :@      @      2@              >@      &@      B@      0@      *@       @      1@      4@      @      7@      F@      E@      9@      :@      &@       @      4@      @      2@              <@      &@      ?@      *@      *@      @      &@      3@      @      6@     �@@      D@      9@       @      �?      @      @                               @              @      @              @      @      �?              �?      &@       @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ��bhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�G��@�	           ��@       	                    �?�u?�fT@b           ��@                           �?Y��J�@p           ��@                           �?g=���@�             m@������������������������       �Z����@9            �Z@������������������������       ������B@P            �_@                           �?<��w�p@�            �x@������������������������       �v��\@Y            `b@������������������������       �I/��6@�            �n@
                            @U*���@�           �@                           @s�psw@d           �@������������������������       ���`�@�           p�@������������������������       �Ɯ9Z��@�            �j@                           @:����	@�            �j@������������������������       ����@9L@p            `d@������������������������       ��ނ�8@            �I@                          �9@�'��xN@1           >�@                          �6@�>Xg�@c           8�@                            @�)���<@�           p�@������������������������       �.����C@%            |@������������������������       ��+S�i�@r            �e@                           @U$9��@�            �@������������������������       ���d>�x@�           `�@������������������������       �����@
@2             U@                           @.ۣ��@�           ��@                           @�(�w�@�           ��@������������������������       ��d[ߨ@C           p~@������������������������       �BkS$bZ@?            �Z@                            �?���ї�@L            �_@������������������������       ���u�H@-             R@������������������������       ��1]���
@            �K@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       pu@     �b@     �S@     �t@      A@     �|@      @     @o@      =@     �}@     �\@     �J@      E@     �K@      n@      M@     0v@     s@     �{@      U@     `a@     �C@      >@     @e@      1@     �n@             @]@      "@     �l@      H@      6@      &@      $@     �Z@      3@      e@     �b@     �p@      B@      L@      .@      0@     �K@      0@     �M@             �B@      @     @Q@      2@      ,@       @      "@      K@      @      D@      I@     @T@      6@      6@      @      �?      ,@       @      9@              0@              C@      @      @      �?      �?      3@      �?      5@      0@     �A@      @      $@              �?      @      �?      "@              @              3@      @       @              �?      *@      �?       @      @      4@       @      (@      @              "@      �?      0@              $@              3@       @      @      �?              @              *@      &@      .@       @      A@      "@      .@     �D@      ,@      A@              5@      @      ?@      *@      "@      �?       @     �A@      @      3@      A@      G@      2@      0@      @      @      1@      @      1@              @       @      @       @      @               @      @      @      *@      0@      1@      $@      2@      @      &@      8@      $@      1@              1@      @      8@      &@      @      �?      @      =@      �?      @      2@      =@       @     �T@      8@      ,@     �\@      �?     @g@              T@       @      d@      >@       @      "@      �?     �J@      ,@      `@     �X@     `g@      ,@      L@      ,@      "@      X@             �c@              L@       @     �a@      8@      @      "@              H@      @      [@      U@     �d@      &@      C@      @      @     �T@             @`@              G@             @[@      .@      @      @              C@      @     @S@     @R@     �`@      "@      2@      "@      @      ,@              <@              $@       @     �@@      "@               @              $@      �?      ?@      &@      >@       @      ;@      $@      @      3@      �?      <@              8@              3@      @      �?              �?      @      @      4@      .@      7@      @      :@      $@       @      *@      �?      5@              ,@              3@      @                              @      @      3@      @      *@       @      �?              @      @              @              $@                              �?              �?      �?              �?      "@      $@      �?     �i@     �[@     �H@     �d@      1@      k@      @     �`@      4@     `n@     �P@      ?@      ?@     �F@     �`@     �C@     `g@     �c@     `f@      H@      a@     �R@      :@     �[@      "@     `d@       @     �R@      *@      g@      D@      $@      ,@     �C@     �R@      8@     ``@      Y@     @X@      B@     �M@     �D@      ,@     �D@       @     @W@       @     �B@      @     �V@      *@       @      @      *@      9@      &@     �O@     �E@     �D@      ,@      E@      :@      @      B@       @      Q@       @      6@      @     �P@      $@      @      @      "@      5@      "@     �F@      :@      A@      &@      1@      .@       @      @              9@              .@              9@      @      @              @      @       @      2@      1@      @      @     @S@     �@@      (@     @Q@      @     �Q@              C@      @     �W@      ;@       @      $@      :@     �H@      *@      Q@     �L@      L@      6@      R@      7@      &@     �P@      @     �P@             �@@      @     �T@      8@       @      @      9@     �A@      "@      M@     �I@     �K@      6@      @      $@      �?       @      @      @              @              &@      @              @      �?      ,@      @      $@      @      �?              Q@     �B@      7@     �K@       @     �J@      @      M@      @      M@      :@      5@      1@      @      N@      .@      L@      L@     �T@      (@     �E@      @@      4@      H@      @     �G@      �?     �L@      @      H@      6@      ,@      (@      @     �G@      ,@      E@      H@     @Q@      &@     �D@      @@      1@     �B@      @     �B@      �?      G@      @     �B@      .@      ,@      (@      @     �F@      &@      ?@      =@      M@      $@       @              @      &@      @      $@              &@      �?      &@      @                      �?       @      @      &@      3@      &@      �?      9@      @      @      @      �?      @       @      �?              $@      @      @      @      �?      *@      �?      ,@       @      *@      �?      ,@      @      @      @      �?      @              �?               @       @      @                       @      �?      "@       @      $@      �?      &@                      @              @       @                       @       @      �?      @      �?      &@              @      @      @        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJjm�shG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@!�P�@�	           ��@       	                     @�qڋ��@           8�@                           �?xr��?1@w           @�@                           @�����@�           H�@������������������������       ��� �`@�            v@������������������������       ��P�M�x
@�            �r@                           �?^� 5E�@�           �@������������������������       ���>��@�            �u@������������������������       ���u@�           @�@
                           �?~��Tܕ@�           `�@                           �?�;|}=@�            �u@������������������������       ���M��@G             [@������������������������       �!�_~@�            @n@                          �1@�	-莇@�            �r@������������������������       ��(eU�n
@6            �T@������������������������       �7h0��K@�            �k@                           �?��%��@�           ��@                          �@@�w��&@�           ��@                            @3B��@�           0�@������������������������       ��!��ڸ@	           �y@������������������������       �i��a��@�            �r@                           @��B3�Y@            �E@������������������������       �ފӘc�@             <@������������������������       ��w��@@
             .@                           @`�^�e�@�           ��@                           @��$p�@            z@������������������������       �nD�'@�            �o@������������������������       ���mC@j            `d@                           �?!��?ܥ@�            �q@������������������������       ���@T            �`@������������������������       ��|�@@_             c@�t�b�?     h�h5h8K ��h:��R�(KKKK��h��B`       ps@      c@     �U@     �v@      A@     �|@      @     `j@      ;@     �~@     �\@      Q@     �E@     @T@     �m@     @Q@     �u@     0r@      {@      V@     @f@      S@     �F@      n@      0@     �v@      �?      _@      *@     �s@      K@      F@      7@      <@     �a@      9@     �l@      g@     �r@     �K@     @\@     �L@      >@     @g@      @      r@             �T@      (@     `l@     �@@      =@      5@      .@     @Y@      .@     �e@     @`@     @o@      E@      K@      &@      "@     �L@      �?     @[@             �B@       @     �X@      $@      @               @     �B@              L@      G@      W@      2@      ;@      @      @      <@      �?      K@              ,@      �?      L@       @      @              @      6@              D@      0@      H@      ,@      ;@      @      @      =@             �K@              7@      �?      E@       @                      �?      .@              0@      >@      F@      @     �M@      G@      5@      `@       @     `f@              G@      $@      `@      7@      9@      5@      @      P@      .@     @]@      U@     �c@      8@      5@      0@      .@     �G@      �?     �A@              5@       @      =@      @      "@      @      @      0@      @      5@      <@      I@      *@      C@      >@      @     �T@      �?      b@              9@       @      Y@      3@      0@      1@      �?      H@       @      X@      L@      [@      &@     @P@      3@      .@      K@      *@     �R@      �?     �D@      �?     �V@      5@      .@       @      *@      E@      $@     �K@     �K@     �I@      *@     �A@       @      "@      4@      (@      A@      �?      2@      �?      E@      4@      &@       @      &@      0@      @      B@      C@      8@      @      (@      @      �?      &@      �?      @              @      �?      ,@       @      @                      @      @       @      (@      $@      @      7@      @       @      "@      &@      <@      �?      &@              <@      2@       @       @      &@      &@      �?      <@      :@      ,@      �?      >@      &@      @      A@      �?     �D@              7@             �H@      �?      @               @      :@      @      3@      1@      ;@      @      "@       @       @      &@      �?      .@              @              4@              @               @      @              @       @      �?       @      5@      "@      @      7@              :@              3@              =@      �?      �?                      6@      @      .@      .@      :@      @     �`@      S@     �D@      ^@      2@      Y@      @     �U@      ,@     @e@      N@      8@      4@     �J@      X@      F@     @^@     �Z@     ``@     �@@     �G@      G@      ?@     �L@      $@     �B@      @      P@      $@     �R@     �A@      0@      (@     �A@     �E@      3@     �R@      J@     @R@      *@     �G@     �A@      <@     �J@      $@     �A@      @      O@      $@     @R@      =@      .@       @     �@@     �D@      1@     @R@     �I@     @R@      *@      =@      ;@      0@      @@      @      6@      @      =@       @      L@      *@      &@      @      (@      7@      $@     �B@      ;@      E@       @      2@       @      (@      5@      @      *@      �?     �@@       @      1@      0@      @      @      5@      2@      @      B@      8@      ?@      @              &@      @      @               @               @               @      @      �?      @       @       @       @      �?      �?                              "@      @      �?                               @                       @      �?      @       @       @       @                                               @              @               @                               @      @                                              �?      �?                     �U@      >@      $@     �O@       @     �O@       @      7@      @     �W@      9@       @       @      2@     �J@      9@     �G@      K@      M@      4@      N@      4@      @      A@      @     �F@              2@             �O@      &@      @      @      @      =@      @      8@      @@      B@      &@      @@      $@      �?      4@      @      >@              2@              B@      @      @      @      @      3@      @      &@      0@      6@      $@      <@      $@      @      ,@              .@                              ;@       @      �?      �?              $@              *@      0@      ,@      �?      :@      $@      @      =@      @      2@       @      @      @      @@      ,@       @      @      *@      8@      2@      7@      6@      6@      "@      4@      @              1@      @      @       @      @      @      (@      @      �?                      ,@      @      "@      *@      @       @      @      @      @      (@              *@               @              4@      "@      �?      @      *@      $@      (@      ,@      "@      1@      �?�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�J2hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?aN�s�w@�	           ��@       	                   �?@��V��@           ��@                           �?�Fb
�E@�           �@                          �8@z+����@[           H�@������������������������       ��#��jR@           �z@������������������������       ��[�	0�@T            �_@                            @�v���Q@s           ��@������������������������       �o�ʁ�@R           ��@������������������������       ��"�n��@!            |@
                           @,D����@C             Z@                            @��Y��
@!            �J@������������������������       ��ַ�@             =@������������������������       �&6G@�9	@             8@                           �?��4���@"            �I@������������������������       ��}ZG�@             &@������������������������       ��Z7[��	@             D@                           @Өc=[@�           С@                          �2@5���J#@|           H�@                           @�r�Eޤ@e             e@������������������������       ������
@C            �Z@������������������������       � M�vB�@"            �N@                          �5@q�?��@           |@������������������������       �;�5B�@j             d@������������������������       ���)є�@�            r@                           �?�־=�@           ��@                           @Hš�:@           H�@������������������������       ��Q��@�            �t@������������������������       �BрW@<            �@                            �?�����>@           ��@������������������������       �*F_�,@�            �i@������������������������       ���U�R@�           H�@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �v@     �\@      X@      v@      E@     @}@      @     �n@      <@     0}@      W@      K@     �@@      M@     �m@     �P@     @w@     s@     �{@      S@     @a@     �I@      Q@     �b@      ?@     �b@      @     �^@      2@     `d@     �B@      9@      1@     �B@      X@      C@     �a@     �a@      e@      A@      `@     �A@      L@     �a@      ;@     @b@      @     �]@      2@     �c@     �@@      8@      &@      @@     �W@     �@@     @a@     ``@      d@      A@      J@      (@      5@     �L@      @     �M@      @     �C@       @     �H@      0@      @      @      @      >@      4@      J@     �C@      Q@      ,@      E@      &@      2@      G@      @      H@              7@       @     �B@      *@      @       @      @      *@      4@      F@      ?@     �J@      (@      $@      �?      @      &@      �?      &@      @      0@              (@      @       @      @      �?      1@               @       @      .@       @      S@      7@     �A@     �U@      7@     �U@      @      T@      0@     �[@      1@      2@      @      ;@     @P@      *@     �U@      W@     @W@      4@      F@      0@      3@      J@       @     �I@       @      A@      $@      S@      @      @      @       @      E@      "@     �B@     �E@      L@      "@      @@      @      0@      A@      .@      B@      �?      G@      @      A@      *@      ,@       @      3@      7@      @     �H@     �H@     �B@      &@      $@      0@      (@       @      @      @              @              @      @      �?      @      @      �?      @      @      "@      @              @      ,@      &@       @      @       @               @                      �?      �?      �?      @      �?      @      �?       @      �?                      "@      @      �?               @               @                              �?               @      �?      @                                      @      @      @      �?      @                                              �?              �?      �?                      �?       @      �?              @       @      �?      @               @               @              @      @              @       @              �?      @      @      @                      �?              �?                               @                      @              �?                      �?              �?      �?              @      �?      �?      @               @                              @                      @       @                      @      @      @             �k@     �O@      <@     `i@      &@     �s@             @^@      $@      s@     �K@      =@      0@      5@     �a@      =@     �l@     �d@      q@      E@     �Q@      2@      @     �I@      @     �U@              B@      @     @R@      7@      @      @      @      I@      *@     �K@     �F@     �F@      1@      @               @      =@              6@              @              8@      @                      @      "@      @      9@      *@      @      @      @               @      *@              ,@              @              .@      @                              "@              8@      @      @      @       @                      0@               @                              "@      @                      @              @      �?       @      @              P@      2@      @      6@      @     @P@              =@      @     �H@      1@      @      @       @     �D@      @      >@      @@      C@      $@      *@      @      @      $@      �?      3@               @              2@       @       @      @              3@      �?      1@      1@      3@      �?     �I@      (@       @      (@       @      G@              5@      @      ?@      .@      @      @       @      6@      @      *@      .@      3@      "@      c@     �F@      5@      c@       @     �l@             @U@      @     �l@      @@      7@      "@      .@     �V@      0@     �e@      ^@     `l@      9@      T@      4@      "@     �T@       @     �`@              A@      @     @^@      @       @      @      @      G@      @     �R@      Q@      ^@      ,@      <@      &@      @      =@      @     �D@              (@      @     �H@       @      @       @      @      ,@      @      A@      <@      H@       @      J@      "@      @     �J@      @      W@              6@      �?      R@      @      @       @      �?      @@              D@      D@      R@      @     @R@      9@      (@     �Q@             �X@             �I@      �?     �[@      9@      .@      @      &@      F@      &@     @Y@      J@     �Z@      &@      (@      $@      @      9@              7@              *@              :@      @      @                      1@      @      0@      @      C@       @     �N@      .@      @     �F@             �R@              C@      �?      U@      5@      (@      @      &@      ;@      @     @U@     �H@     @Q@      "@�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�ĠhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��-��@�	           ��@       	                     @���w�@9           ��@                            �?��2TJ@k           ��@                          �:@k��XӾ@>           �@������������������������       �:1S��=@�            �y@������������������������       ������@?             X@                            �?X�蜺R@-           �}@������������������������       �I=7@�            �u@������������������������       �o�$�b�@R            �_@
                           @ �
k.@�           H�@                          �9@ l��@�           ��@������������������������       �(˓�x
@5           �}@������������������������       �<�6��@e            @c@                           @X��j�@4            �T@������������������������       �x�iz.@+            �Q@������������������������       ����@	             (@                          �6@m���z@�           P�@                           @���_@�            �@                          �1@�N#@�           @�@������������������������       ��W:�F
@�            �v@������������������������       ���[0�@	           �@                            �?�5d6v(@�            �w@������������������������       ��?-k2�@6            @W@������������������������       �51r�LB@�            �q@                           @j�M@�            �@                          �7@��� @7           �}@������������������������       �*��ăx
@A            �Y@������������������������       ���}���@�            �w@                          �:@�2�+��@x             h@������������������������       ������@R            �a@������������������������       �H�p
�
@&             J@�t�bh�h5h8K ��h:��R�(KKKK��h��B`        t@     �]@     @V@     �v@     �F@     �}@      @      i@      @@     `{@      X@     �R@     �D@     �R@     �o@     �R@     �x@     �r@     �{@     �S@     �`@     �L@     �M@     `d@     �@@     �`@      @     �Z@      3@     �d@      J@      D@      3@      L@     �\@      ?@      a@      c@     �f@     �B@     �P@     �@@      <@     @Y@      .@     �S@       @      P@       @     �\@      :@      9@       @      :@     �P@      7@     �Q@     �S@      `@      6@      ;@      3@      ,@      H@      &@      C@       @      D@      @     �L@      @      *@      @      2@      A@      2@      ?@      D@      Q@      *@      ;@      (@      @      B@      &@      A@       @      =@      @      J@      @      $@       @      &@      :@      *@      9@     �@@     �N@      &@              @      @      (@              @              &@              @      �?      @      @      @       @      @      @      @      @       @     �C@      ,@      ,@     �J@      @     �D@              8@      �?      M@      3@      (@       @       @     �@@      @     �C@      C@      N@      "@     �@@      @      ,@      E@      �?      =@              ,@      �?      A@      0@      $@       @      @      8@      @      >@      ?@     �E@      @      @      @              &@      @      (@              $@              8@      @       @              @      "@              "@      @      1@      @     �P@      8@      ?@      O@      2@     �K@      @      E@      &@      J@      :@      .@      &@      >@     �G@       @     �P@     �R@     �J@      .@     �L@      1@      >@      L@      .@      I@      @      D@      &@      E@      6@      ,@      $@      9@     �A@      @     �M@     @R@      J@      ,@     �F@      "@      4@      A@      *@      H@       @      9@      &@      B@      4@      *@       @      1@      6@      @     �G@     �K@      A@      *@      (@       @      $@      6@       @       @       @      .@              @       @      �?       @       @      *@              (@      2@      2@      �?      $@      @      �?      @      @      @               @              $@      @      �?      �?      @      (@      @       @       @      �?      �?      @      @      �?      @      @      @              �?              $@      @      �?      �?      @      "@      @      @      �?      �?      �?      @       @                                              �?                      �?                              @              �?      �?                     �g@     �N@      >@     �h@      (@     �u@             �W@      *@     �p@      F@      A@      6@      3@     �a@      F@      p@      b@     @p@     �D@      Z@     �A@      3@     �b@      �?     0q@              M@       @     �i@      5@      9@      .@      "@     �U@      6@     �g@     �X@     �h@      5@     @S@      2@      1@      ]@      �?      i@             �J@       @     �e@      .@      2@      (@      @     @Q@      ,@     @`@     @P@      d@      3@      3@      �?      @      =@      �?     �S@              ;@              O@      �?      @              @       @      @      G@      5@      I@      @      M@      1@      $@     �U@             �^@              :@       @     @\@      ,@      .@      (@      @     �N@       @      U@      F@     �[@      .@      ;@      1@       @      @@             �R@              @      @      @@      @      @      @      @      2@       @     �N@      A@     �C@       @      @      @              ,@              @                              "@      �?      �?                      @              4@      ,@      *@              6@      $@       @      2@             @Q@              @      @      7@      @      @      @      @      ,@       @     �D@      4@      :@       @     @U@      :@      &@     �H@      &@     �Q@              B@      @      P@      7@      "@      @      $@     �J@      6@     @P@     �F@     �N@      4@      L@      2@      $@      ?@      $@     �O@              8@      @      G@      ,@      "@      @      "@     �C@      $@      F@      <@     �F@      ,@      8@      �?      @      $@              "@                      @      "@      �?                              (@              (@       @      @      @      @@      1@      @      5@      $@      K@              8@             �B@      *@      "@      @      "@      ;@      $@      @@      4@      E@      &@      =@       @      �?      2@      �?      @              (@              2@      "@              @      �?      ,@      (@      5@      1@      0@      @      5@       @              .@              @              @              ,@      @              @              *@      &@      $@      .@      $@      @       @              �?      @      �?                      @              @      @                      �?      �?      �?      &@       @      @      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�A9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?';y]�@�	           ��@       	                    �?f��
@           0�@                           @q*l�&@Z           x�@                          �9@�M<7�.@�             n@������������������������       �'�L���@z            �g@������������������������       �\���ٕ@%            �I@                           �?�z)��@�            �q@������������������������       �����
!@>            �X@������������������������       ������@}            �g@
                           @���[�@�           ��@                           @�nc2�@�           ��@������������������������       �!��b�'@�           ��@������������������������       �K7��/@�            pp@������������������������       �R�֯�$@             8@                           �?��<,�@�           ��@                          �<@U*GP�r@=           ��@                            �?b��a@$            �@������������������������       ��^wj+�
@3           �}@������������������������       �q"���s@�            �x@                            �?Qq���@            �F@������������������������       �"Bv�@             ?@������������������������       �^,Eal�@             ,@                           @@�a��@k           ��@                          �6@§�Yu�@l           ��@������������������������       �m��:3@            y@������������������������       ����5Vt@l            �d@                           @a�u�.@�           ��@������������������������       ��V�E@�           ��@������������������������       ����.@t            �f@�t�bh�h5h8K ��h:��R�(KKKK��h��B        Pv@      c@     �T@     �v@      @@     �~@      &@     �k@     �@@     �|@      Y@      K@      B@      M@     `o@     �M@      u@     �t@     `y@     �T@     �`@     @T@      L@     @b@      :@      a@      &@      [@      8@     �b@      I@      @@      5@     �C@     �X@      >@     �\@     @c@     `d@      D@     �H@      2@      8@     �D@      @     �I@      @      >@      "@      I@      2@      @      @      @      ?@      *@      ?@     �I@      S@      "@      :@      @       @      7@       @      >@       @      2@      "@      ,@      $@      @      @      @       @      $@       @      5@      @@      @      3@      �?       @      2@       @      ;@       @      &@       @      *@      $@      @               @      @      "@      @      .@      ?@       @      @      @              @              @              @      �?      �?               @      @      �?      @      �?      @      @      �?       @      7@      ,@      0@      2@       @      5@       @      (@              B@       @      �?       @      @      7@      @      7@      >@      F@      @      (@      @       @      �?              @                              0@              �?              @      @       @      @      (@      2@      @      &@      &@       @      1@       @      1@       @      (@              4@       @               @              0@      �?      0@      2@      :@       @     @U@     �O@      @@     @Z@      6@     �U@      @     �S@      .@     �X@      @@      :@      0@      @@     �P@      1@     �T@     �Y@     �U@      ?@     �T@     �K@      @@     @Z@      5@     �U@      @      S@      .@     �X@      >@      :@      0@      @@      O@      1@     �T@     @Y@     �U@      ?@      K@      F@      8@     @R@      2@     �L@      @     �M@      *@     �Q@      9@      0@      (@      9@      I@      &@     @R@     �T@      O@      7@      =@      &@       @      @@      @      =@              1@       @      <@      @      $@      @      @      (@      @      "@      3@      8@       @       @       @                      �?                       @                       @                              @              �?       @      �?             �k@     �Q@      ;@      k@      @     v@             �\@      "@     Ps@      I@      6@      .@      3@      c@      =@     �k@      f@     `n@     �E@      S@      0@      &@      S@             �f@              J@      �?     @_@      .@      @      �?      @     �K@      @     �V@     �P@     �\@      3@     �R@      0@      &@      S@              e@              J@      �?      ]@      .@      @              @     �I@       @     �V@      O@     @[@      1@     �D@      *@      @     �F@             �T@             �A@      �?     �Q@      @                      �?      5@      �?     �I@      >@     �P@      @     �@@      @      @      ?@             �U@              1@              G@      (@      @              @      >@      �?     �C@      @@     �E@      $@       @                                      ,@                              "@                      �?      �?      @       @              @      @       @       @                                      "@                              @                              �?      @       @              �?      @                                                      @                               @                      �?              �?                      @               @     `b@     �K@      0@     �a@      @     @e@             �O@       @      g@     �A@      3@      ,@      ,@     �X@      9@     �`@     �[@      `@      8@     �O@      6@      @      P@             �P@              >@      @     �X@      &@      @      @      @      D@       @     �E@     �F@     �F@      *@      <@      "@      @      H@             �K@              =@              R@      @      @      @              >@       @      A@      ;@     �A@      (@     �A@      *@              0@              &@              �?      @      ;@      @      �?      �?      @      $@              "@      2@      $@      �?      U@     �@@      $@      S@      @      Z@             �@@      @     @U@      8@      *@      "@      &@      M@      7@     @V@     @P@     �T@      &@     �O@      ;@      @      Q@      @     �T@              8@      @     �Q@      2@      "@      @      &@     �A@      0@     @P@      G@      R@      &@      5@      @      @       @      �?      6@              "@              .@      @      @      @              7@      @      8@      3@      &@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ|��qhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�6gl�@�	           ��@       	                    �?����@           t�@                          �:@���N��@b           @�@                          �9@2.U�|C@)           p~@������������������������       ��0a+�K@           �|@������������������������       �ϓiI@             ?@                          �=@(d��t�@9            @X@������������������������       ��@"`�@!            �N@������������������������       �B1�8�@             B@
                           �?�1�=@�           T�@                          �3@o�|�W@�            �t@������������������������       ��_�+	@D            �Z@������������������������       �ߴ�m@�            �l@                            @D]�"!T@�           0�@������������������������       �B�V+�S@�            �z@������������������������       ��t��@�            �u@                          �6@�n��f�@�           X�@                           @����+@�           ��@                          �4@e|��@            ؊@������������������������       ����@�           ��@������������������������       �G���#�@�             i@                           �?��u��@�           ��@������������������������       ��`VN�@�            @q@������������������������       ��ůyD@�             x@                           �?@vC2�@�           �@                          �9@�|��@�            0v@������������������������       ��'P��@w             i@������������������������       ��v`p��@b            @c@                           @�P���S@�            �u@������������������������       ��z.�@�            �h@������������������������       �y��T�
@a            �b@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       `t@     `b@      X@     Pu@      G@     @|@      "@     �o@      >@     Pz@      U@     @P@     �B@     �Q@     @n@      T@     Pv@     r@     �|@     �Y@     �a@     �S@      N@      c@      >@     �`@      "@     @`@      7@     �d@     �I@     �@@      7@     �G@      V@     �C@     @`@     �^@     �f@     �I@     �F@      8@      2@     @P@      @      J@       @      ?@      @     �P@      3@      @      @      *@      =@      4@     �D@     �D@      U@      *@      F@      4@      *@      M@      @      F@              8@      @     �J@      *@      @      �?      $@      9@      2@     �B@      D@      Q@       @      C@      .@      *@     �J@      @      D@              5@      @     �J@      *@      @      �?      $@      6@      2@     �B@     �C@      P@       @      @      @              @              @              @                                                      @                      �?      @              �?      @      @      @               @       @      @              ,@      @       @      @      @      @       @      @      �?      0@      @              �?      @      @               @       @      @              @      @      �?      @       @      @              @              ,@      @      �?      @              @              @              �?              "@      @      �?              �?      �?       @              �?       @       @     @X@     �K@      E@     �U@      ;@     �T@      @     �X@      2@     �X@      @@      <@      0@      A@     �M@      3@     @V@     @T@     �X@      C@      5@      .@      (@      8@       @      3@              D@      @     �B@      ,@      @      @      &@      6@      �?     �D@      1@      >@      .@      @      @      @       @      �?      &@              (@              2@       @              �?              &@               @      "@      2@              2@      (@      @      6@      �?       @              <@      @      3@      (@      @      @      &@      &@      �?     �@@       @      (@      .@      S@      D@      >@     �O@      9@      P@      @     �M@      .@      O@      2@      7@      $@      7@     �B@      2@      H@      P@     @Q@      7@     �B@      ;@      ,@      D@      "@      :@      @      =@      $@      E@      @      *@      @      (@      9@      0@      7@      =@      F@      .@     �C@      *@      0@      7@      0@      C@       @      >@      @      4@      (@      $@      @      &@      (@       @      9@     �A@      9@       @      g@      Q@      B@     �g@      0@     �s@              _@      @     �o@     �@@      @@      ,@      8@     @c@     �D@     `l@     �d@     �q@      J@     �T@      D@      6@     @_@       @     �o@             �W@      @      f@      4@      <@      (@      (@     �[@      7@     `d@      \@      i@      >@      F@      6@      (@     �T@      @     ``@              G@      @      U@      .@      7@       @      @     �P@      6@      X@     @R@     @X@      5@      =@      ,@       @     @R@      @      X@             �A@             @Q@      &@      3@      @       @      G@      .@      R@     �N@     �U@      *@      .@       @      @      $@      �?     �A@              &@      @      .@      @      @      @      @      4@      @      8@      (@      $@       @     �C@      2@      $@      E@       @      _@             �H@       @      W@      @      @      @      @      F@      �?     �P@     �C@     �Y@      "@      5@      @      @      5@      �?     �G@              ;@       @      >@                              @      ;@      �?      6@      *@     �H@       @      2@      .@      @      5@      �?     @S@              6@              O@      @      @      @              1@             �F@      :@      K@      @     @Y@      <@      ,@      P@       @      O@              =@       @     �S@      *@      @       @      (@      F@      2@      P@     �K@      T@      6@      M@      &@      "@     �A@      @      ?@              0@       @      F@      $@      @              �?      8@      &@      5@      :@      @@      0@     �@@      @      @      ;@              4@               @      �?      ;@      @                              3@               @      2@      .@      "@      9@      @      @       @      @      &@               @      �?      1@      @      @              �?      @      &@      *@       @      1@      @     �E@      1@      @      =@      @      ?@              *@             �A@      @      �?       @      &@      4@      @     �E@      =@      H@      @      5@      &@       @      9@      @      1@              $@              4@      @      �?       @      @      &@      @      4@      .@      5@      @      6@      @      @      @              ,@              @              .@                              @      "@              7@      ,@      ;@       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJXlJ3hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?}[�ߘ�@�	           ��@       	                     @��B�I@?           ̔@                          �;@���fN�@u           p�@                          �1@�=�*@K           @�@������������������������       ��{��,
@~            �i@������������������������       ��?�OX@�           І@                            �?܌�vY{@*            �Q@������������������������       �q��Up�@"             N@������������������������       �q�y	O�@             $@
                          �9@��	z@�            Pt@                          �5@M�
2�@�            pq@������������������������       ��p�u�@i            �d@������������������������       ���l)@B            @\@                           �?F�@             G@������������������������       �!.�ߵ
@             <@������������������������       ��xb嫯@             2@                          �;@�p W.=@V           ,�@                           �?�1OJ��@y           f�@                           @���q�@+           �@������������������������       ��Ib.f?@a           ��@������������������������       �������@�            @t@                            �?�Rj�X@N           D�@������������������������       ��a�4@�           ��@������������������������       �K���8�@o           ��@                           @�C���@�            0v@                          �?@���.�@�            `r@������������������������       ��㔇Ҫ@|            @h@������������������������       ������@?             Y@                           @�����@"            �N@������������������������       �p�Ͷ��@
             4@������������������������       �֛�U�	@            �D@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �t@     �^@     @V@     �t@     �C@     �~@       @     `k@      @@     }@     �[@     @Q@     �F@     @R@     `m@      O@     �y@      q@     {@      T@      Y@      5@      7@     @Z@      "@     �f@      �?     �U@      @     �e@     �C@      *@      "@      2@     �T@      @      c@     @U@      g@      ?@     �R@      2@      0@     �V@      @     @b@              O@      @     `a@      3@      &@       @      "@     �O@      @     @[@     �P@      b@      1@     @R@      0@      &@     @U@      @     @a@              O@      @      `@      ,@      $@      �?      @      M@       @     @Z@     �N@     `a@      1@      "@              @      "@      �?      >@              "@      @     �C@      �?       @                      0@      �?      3@      3@     �E@       @      P@      0@       @      S@      @      [@             �J@      �?     �V@      *@       @      �?      @      E@      �?     �U@      E@      X@      .@      �?       @      @      @               @                              $@      @      �?      @       @      @      @      @      @      @              �?      �?      @      @              @                              $@      @              @       @      @      @      @      @      @                      �?                              @                                              �?       @                              �?      �?                      :@      @      @      ,@      @     �B@      �?      9@       @      B@      4@       @      �?      "@      4@       @     �E@      2@      D@      ,@      7@       @      @      "@      @      B@              8@      �?     �@@      2@              �?      "@      0@       @     �C@      *@      C@      @      0@              @      @      @      <@              &@      �?      (@      "@              �?      @      (@      �?      1@      @      >@      @      @       @               @               @              *@              5@      "@                      @      @      �?      6@      "@       @      @      @      �?       @      @       @      �?      �?      �?      �?      @       @       @                      @              @      @       @      @      @      �?       @      @                      �?      �?      �?                                              @              @      @       @      �?                              �?       @      �?                              @       @       @                      �?                                      @     �l@     @Y@     �P@     �k@      >@     0s@      @     �`@      :@      r@     �Q@      L@      B@     �K@      c@     �K@     0p@     `g@      o@     �H@     `h@     @P@     �I@     @i@      6@     �r@      @     @Z@      7@     �o@     �N@     �I@      ;@      C@     @a@      H@     `m@     �b@      k@      E@      R@      6@      .@     @U@      $@     �_@       @     �A@      @     @Y@      5@      0@      $@      @      H@      &@     �Y@     @P@     �Y@      0@     �D@       @      @     �J@      "@      V@       @      9@       @     �R@      (@      $@      $@      �?      4@      &@     �J@      @@      S@      $@      ?@      ,@      $@      @@      �?     �C@              $@      �?      ;@      "@      @               @      <@             �H@     �@@      :@      @     �^@     �E@      B@     @]@      (@     �e@       @     �Q@      4@      c@      D@     �A@      1@     �A@     �V@     �B@     �`@     �U@     �\@      :@      S@      ;@      4@     �R@      @      V@              >@      (@     �V@      3@      ;@      @      7@     �E@      ;@     �I@     �H@      T@      4@     �G@      0@      0@      E@      "@     @U@       @      D@       @      O@      5@       @      &@      (@     �G@      $@     �T@     �B@      A@      @      B@      B@      .@      5@       @      @      @      ;@      @     �B@      $@      @      "@      1@      ,@      @      8@      B@     �@@      @      =@      <@      $@      4@      @      @      �?      ;@      @     �A@       @      @      @      &@      $@      @      2@      A@      5@      @      4@      (@      @      2@      @      @      �?      4@      @      :@      @      @      @       @      "@      @      .@      (@      .@      @      "@      0@      @       @              @              @              "@      @      �?      @      @      �?      @      @      6@      @      @      @       @      @      �?       @               @                       @       @               @      @      @              @       @      (@               @       @                                                                                       @               @              @      �?       @              @              @      �?       @               @                       @       @                      @       @              @      �?      $@        �t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�X*hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@~�B��@�	           ��@       	                     @����<�@           �@                           �?�c$;�@s           �@                          �3@c����}@K            �@������������������������       ��z����@�            �o@������������������������       �$�%x�@�            �p@                            �?���pi*@(           ԓ@������������������������       �._w��4@R           X�@������������������������       �Q��k�@�            �t@
                          �0@D���*@@�           P�@                           �?( ��	@!            �N@������������������������       �4hSU�@             9@������������������������       �}�+2t�@             B@                           �?d\��2@y           h�@������������������������       ��OG�@�            �t@������������������������       ���Ԥ_@�            0p@                           @� ��N�@�           �@                           �?�=���@�           �@                           �?s��ɚJ@d           ��@������������������������       ��s�/%@�            �k@������������������������       �P)��,B@�            `u@                           @ ����@G           8�@������������������������       ���Э@l            �d@������������������������       � D9Ed@�             v@                           @0k����@�            �x@                          �9@��0dZ@�            @r@������������������������       ���w�@O             `@������������������������       � IY�y6@n            �d@                           @��}E
@A            �Y@������������������������       �yX�y�@             <@������������������������       ��Sy�	@0            �R@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@     `b@      V@     �v@     �E@     �@      (@     �m@      @@     �z@     �Y@     �P@      >@     �P@     �n@     �L@     0w@     Ps@      y@     �P@     @i@      W@      G@     @l@      2@     �x@      @     �a@      (@     pq@      J@     �D@      "@      ;@     �a@      =@     �m@     @g@     �p@      @@      `@     �N@      <@     `f@      @     �r@      �?      Y@      &@      k@     �B@      @@       @      @     �Y@      9@     �e@     @`@     �k@      9@     �G@      1@      ,@     �P@      �?      K@      �?      @@      @     �M@      &@      3@       @      @      7@      0@     �C@      D@      K@      $@      4@      $@      "@      @@      �?      4@              .@       @      7@      @      (@      �?      �?      0@      @      $@      ?@     �B@      @      ;@      @      @     �A@              A@      �?      1@      @      B@      @      @      �?      @      @      (@      =@      "@      1@      @     �T@      F@      ,@      \@       @     @n@              Q@      @     �c@      :@      *@      @       @      T@      "@     �`@     �V@     �d@      .@     @Q@     �D@      (@     @V@      �?      d@             �F@             @^@      3@       @      @      �?      M@      "@     �X@     �Q@     �^@      &@      *@      @       @      7@      �?     �T@              7@      @      B@      @      @      �?      �?      6@             �B@      4@      F@      @     @R@      ?@      2@     �G@      .@      X@       @     �D@      �?     �O@      .@      "@      �?      4@     �B@      @      P@      L@      I@      @      $@       @      @      @              *@       @                      &@      �?                       @       @              �?      @      �?      �?                                              &@                              @                               @      �?              �?      @              �?      $@       @      @      @               @       @                      @      �?                              @                              �?             �O@      =@      .@      F@      .@     �T@             �D@      �?      J@      ,@      "@      �?      2@      =@      @     �O@     �J@     �H@      @      >@      5@       @      3@      *@      D@              ;@      �?      6@      @       @      �?      1@      2@              B@     �A@      7@      @     �@@       @      @      9@       @     �E@              ,@              >@       @      �?              �?      &@      @      ;@      2@      :@      �?     �a@     �K@      E@      a@      9@      \@      "@      X@      4@      c@      I@      :@      5@     �C@      Z@      <@     �`@     �^@     @`@      A@     �X@      @@      >@     �Z@      ,@     �X@      "@     �Q@      1@      Z@     �F@      9@      "@     �@@     @Q@      ,@     �W@     �W@     @W@      ;@     �B@      5@      6@      K@      @     �@@      "@      F@      (@      D@      B@      4@      @      1@     �A@      &@      L@     �E@     �H@      *@      @      @      @      .@      �?      ,@       @      4@      @      5@      4@      &@       @      �?      6@      @      ;@      3@      .@      "@      ?@      2@      .@     �C@      @      3@      @      8@      "@      3@      0@      "@      @      0@      *@      @      =@      8@      A@      @      O@      &@       @      J@      "@     @P@              :@      @      P@      "@      @       @      0@      A@      @     �C@     �I@      F@      ,@      0@      @              *@      @      @@              $@      �?      0@      @       @       @       @      &@       @      @      .@      .@       @      G@      @       @     �C@      @     �@@              0@      @      H@      @      @              ,@      7@      �?     �@@      B@      =@      @      F@      7@      (@      >@      &@      ,@              :@      @      H@      @      �?      (@      @     �A@      ,@      C@      =@     �B@      @      >@      6@      (@      5@      &@       @              9@      @      ;@      @      �?      (@      @      7@      "@      >@      ,@      >@      @      "@      &@       @      (@      @      @               @      @      $@      @              $@      �?      *@      �?      1@      @       @      �?      5@      &@      @      "@      @      @              1@              1@              �?       @      @      $@       @      *@      $@      6@      @      ,@      �?              "@              @              �?              5@       @                              (@      @       @      .@      @       @      @                      @              �?              �?              @       @                                       @      @      @                      "@      �?              @              @                              1@                                      (@      @      @      $@      @       @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�;OhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?'*�r�@�	           ��@       	                     �?�����@�           |�@                          �4@�;��@+           �|@                           �?��(��@k            �f@������������������������       ��c���0
@1            �V@������������������������       �������
@:            @W@                           �?v=���@�            `q@������������������������       ���R$X5@>             W@������������������������       ��	�^X6@�            @g@
                          �:@#BT�m�@�           H�@                          �8@����s@6           (�@������������������������       �l��Az�@�           �@������������������������       �q���}@S            @`@                           �?d����@�            �m@������������������������       ��*�b��@/            @Q@������������������������       ��9׵�@d             e@                           �?V&"��N@�           ԡ@                          �4@��U�Y@            P�@                            �?E.0�L�
@2           �}@������������������������       �έ�7�@P             _@������������������������       ��;p#��	@�            �u@                            @�n�+D@�            �t@������������������������       �J��[@�            0q@������������������������       �l�Uy�@%             N@                          �6@a�-O��@�            �@                          �5@�hv|�@x           ��@������������������������       ��a�@            8�@������������������������       �p�U��j
@X            `a@                            �?�2gF@>           �~@������������������������       �A�ZlT@�            �q@������������������������       ����?�@�            `j@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       �u@      b@     �S@     �u@      D@     ��@      @     @k@      =@     P{@     @Z@     �M@      E@     �L@     �o@     @S@     `u@     �t@      y@     �Q@     �`@     �T@      G@      a@      :@     �e@      @      \@      8@     �`@     �H@      A@      6@     �D@      Y@      @@     �a@     �b@     �b@     �A@      7@      8@       @      C@      $@     �J@       @      A@      @      E@      $@      @      @      ,@      >@      @      7@      H@     �P@      0@       @               @      0@      �?      6@              ,@              8@      @      @      �?      �?      0@              @      0@     �B@      @      �?               @       @              $@              @              "@      @      @                      @              @      @      :@      @      �?              @       @      �?      (@              @              .@      @              �?      �?      (@               @      (@      &@              5@      8@              6@      "@      ?@       @      4@      @      2@      @      �?      @      *@      ,@      @      0@      @@      >@      "@      @      $@              @              *@              @       @      @      �?               @      @      @      �?      @      *@      &@       @      2@      ,@              .@      "@      2@       @      0@      @      *@       @      �?      @      @      @       @      &@      3@      3@      @     �[@     �M@      C@     �X@      0@     �^@      @     �S@      3@     �V@     �C@      =@      0@      ;@     �Q@      =@     @]@     �Y@      U@      3@     �V@      B@      <@     @T@      ,@      \@             �M@      2@     @S@      >@      6@      (@      3@     �L@      0@     @Z@     �S@      N@      2@      T@      ?@      6@      S@      *@     �W@              E@      ,@     �P@      >@      4@      (@      1@      C@      0@     �U@     �R@     �J@      1@      $@      @      @      @      �?      2@              1@      @      &@               @               @      3@              2@      @      @      �?      5@      7@      $@      2@       @      $@      @      3@      �?      ,@      "@      @      @       @      *@      *@      (@      7@      8@      �?      @      @       @       @              @      @       @      �?      "@       @       @       @      �?      �?              @      @      (@      �?      2@      0@       @      0@       @      @       @      1@              @      @      @       @      @      (@      *@      @      1@      (@             `j@     �N@      @@     `j@      ,@     `v@             �Z@      @      s@      L@      9@      4@      0@      c@     �F@     @i@     `f@      o@      B@     �L@       @      0@      T@      @     �a@              G@              ]@      6@       @      �?      @     �G@      "@     @R@     �M@      X@      7@      ?@      @      @      N@      �?     �V@              <@              Q@      1@                       @      .@      @      D@      >@     �Q@      @      $@              �?      0@              .@              @              6@      @                              "@      @      "@      &@      (@      @      5@      @      @      F@      �?      S@              5@              G@      ,@                       @      @      �?      ?@      3@     �M@              :@      @      "@      4@      @      J@              2@              H@      @       @      �?      @      @@      @     �@@      =@      9@      2@      7@      @      @      0@      @      H@               @              F@      @      �?      �?      @      8@       @      >@      :@      6@      "@      @               @      @       @      @              $@              @       @      �?                       @       @      @      @      @      "@     @c@     �J@      0@     ``@       @     �j@              N@      @     �g@      A@      7@      3@      $@     @Z@      B@      `@      ^@      c@      *@     �T@      :@      &@     @V@      @     �d@              G@      �?      `@      6@      5@      "@      @     �O@      5@     �X@      R@     �[@      @     @P@      :@      @      R@       @     �_@              E@              ^@      2@      2@      "@      @      I@      5@     �U@     �P@      Y@      @      2@              @      1@      �?     �B@              @      �?      "@      @      @                      *@              (@      @      $@      �?     �Q@      ;@      @      E@      @     �I@              ,@      @     �M@      (@       @      $@      @      E@      .@      >@      H@     �E@       @      H@      ,@      @      5@      �?      A@              @      @      :@      (@      �?      @      @      ;@      @      5@      :@      :@      @      7@      *@       @      5@      @      1@               @             �@@              �?      @      @      .@      (@      "@      6@      1@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJPFHhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?:M�]�@�	           ��@       	                     @c��	�@"           ԙ@                          �6@i�6�t@k           �@                          �4@�ʼ�v@C            @������������������������       �ܔ2���@�            @u@������������������������       ���:���@g            �c@                            �? {t@(           �|@������������������������       ���h���@           Py@������������������������       ���fIV	@!             K@
                          �9@nff��(@�           ��@                           @O�/�!�@J           ��@������������������������       ����9;�@(           �|@������������������������       �>)?R}�@"            @P@                           �?Ֆ���@m             e@������������������������       ��OA�e�
@            �A@������������������������       �R�˫��@Y            �`@                           �?�Ğ��<@�           ��@                           �?=߄.�I@           �@                            @���q@�           h�@������������������������       �����@�           �@������������������������       ���;+�@X             b@                           @�X�+��@5             U@������������������������       �/�F��@#            �J@������������������������       ���Y	�@             ?@                          �5@�F ��@�           L�@                           @�@�8��@           @�@������������������������       ���iH @�            �u@������������������������       �p����@-           �~@                          �6@�lkp�@u           X�@������������������������       �5b$8@N             ^@������������������������       ���mJT�@'           0}@�t�bh�h5h8K ��h:��R�(KKKK��h��B`       s@     �`@     �Y@     @v@      8@     �~@      @     �l@     �B@      {@      ]@     �O@      A@     @R@     �o@     �Q@     �u@     �r@     �|@     �Q@     �_@     @Q@      P@     �`@      3@     �a@      @      _@      =@     `b@      M@     �@@      7@     �H@      _@     �B@     �_@      a@     �e@     �@@     @P@      E@     �@@     �U@      @      U@      @     �P@      (@      Y@      8@      0@      (@      6@     �R@      =@     �S@     �N@     �^@      5@     �C@      $@      0@     �J@       @      K@              <@      (@     �K@      "@      @      @      .@      :@      ,@      >@      @@      T@      .@      >@      @      *@     �A@      �?     �@@              0@      @      D@      "@       @       @      @      6@      "@      2@      7@      M@      .@      "@      @      @      2@      �?      5@              (@      @      .@              @      �?      &@      @      @      (@      "@      6@              :@      @@      1@     �@@      @      >@      @      C@             �F@      .@      &@      "@      @      H@      .@      H@      =@     �E@      @      7@      <@      1@      :@       @      ;@      @      A@              >@      .@      @      "@      @     �E@      .@     �F@      =@     �C@      @      @      @              @      �?      @              @              .@              @                      @              @              @             �N@      ;@      ?@     �G@      ,@      M@       @      M@      1@     �G@      A@      1@      &@      ;@      I@       @     �H@      S@      I@      (@      F@      *@      8@      A@      $@     �K@              H@      "@     �E@      :@      .@       @      6@      C@      @     �F@     �J@      <@      $@     �@@      "@      8@      ?@      $@     �E@             �F@       @     �C@      8@      .@      @      1@      B@      @     �A@      I@      :@      $@      &@      @              @              (@              @      �?      @       @              @      @       @              $@      @       @              1@      ,@      @      *@      @      @       @      $@       @      @       @       @      @      @      (@      @      @      7@      6@       @       @      @      �?                       @       @       @      @               @                      �?       @              �?              @      �?      "@      "@      @      *@      @      �?               @      @      @      @       @      @      @      $@      @      @      7@      1@      �?     `f@      P@     �C@     �k@      @     �u@      �?     �Z@       @     �q@      M@      >@      &@      8@     @`@     �@@     @k@     �d@      r@      C@     �M@      &@      ,@      S@       @     �c@              F@      �?     �Z@      4@      "@      �?      @     �H@      @      Q@      O@     �\@      :@     �H@      $@      *@     �Q@      �?      a@             �D@      �?     �X@      1@       @      �?      @      G@      @      P@      N@     �W@      :@      C@      @      &@      N@      �?     @^@              :@      �?     �T@      @      @      �?       @      D@      @     �J@      L@     �R@      .@      &@      @       @      $@              .@              .@              0@      $@      @              @      @      @      &@      @      5@      &@      $@      �?      �?      @      �?      6@              @               @      @      �?                      @              @       @      3@              @                      @      �?      3@               @              �?              �?                       @              @       @      (@              @      �?      �?                      @              �?              @      @                              �?              �?              @              ^@     �J@      9@     `b@      @     �g@      �?     �O@      @     �f@      C@      5@      $@      3@     @T@      :@     �b@      Z@      f@      (@      H@      ;@      ,@     �T@             @]@              F@      �?     �Z@      .@      1@       @      @      J@      .@      X@     @P@      ^@      @      6@       @      @      @@             �K@              8@             �O@      @      @      @              3@      @      B@      7@      D@      @      :@      3@      $@      I@              O@              4@      �?      F@      &@      (@      @      @     �@@      $@      N@      E@      T@       @      R@      :@      &@     @P@      @     �R@      �?      3@      @     @R@      7@      @       @      ,@      =@      &@      K@     �C@      L@      @      (@              @      0@      @      4@              @       @      2@      @      �?                      @              (@      @      @      �?      N@      :@      @     �H@              K@      �?      (@      @     �K@      0@      @       @      ,@      9@      &@      E@     �A@     �H@      @�t�bubhhubh)��}�(hh.hhhKhK	hKhG        hhMhNhJ�.�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �3@F��v�@�	           ��@       	                    @�4#!Z@n           l�@                           �?r"�;@�           8�@                          �2@,��'@�            �t@������������������������       ���Θ1@�             m@������������������������       �?8� }@C            �Y@                            @Ve���
@�            �@������������������������       �6����	@~           ؂@������������������������       �7�k)�9@g            �d@
                           @�j3�@�            �p@������������������������       �R��Vv�@             3@                           @	L�?�@�            @o@������������������������       �M�q���@y             g@������������������������       ����!�@-            @P@                           �?C�8�Xv@9           ܣ@                            @kX)�" @�            �@                          �?@f��ϖ�@�           ��@������������������������       ��A�ztB@�           @�@������������������������       ��"��[@              K@                           @4�P��1@&            ~@������������������������       � <�w@|             j@������������������������       ������@�             q@                          �7@�E]�T@f           ��@                          �5@�G�M=�@�           ��@������������������������       ��tVͧ�@           p{@������������������������       �{rX�Պ@�            �u@                           @�D���@x           ��@������������������������       ��/"��T@�            0q@������������������������       ��/��@�            �t@�t�bh�h5h8K ��h:��R�(KKKK��h��B        �t@     @a@     �W@     0w@      C@     �}@      "@     @k@      E@     �{@      \@      I@      @@     �M@     �n@      K@     Pw@     pr@     `{@     @V@      S@      @@      5@     �a@       @     �l@      �?      M@       @      h@      9@      3@      @      (@      U@      @     ``@     �W@     `j@      9@     �L@      :@      (@     �X@       @      f@      �?     �G@       @     �e@      4@      1@      @      "@     �O@      @     �[@     @Q@     �f@      6@      0@      "@      "@     �D@      @      ?@      �?      &@       @     �A@      @      @      @      @      6@       @      ?@      <@      M@      $@      @      @      @      >@      @      5@      �?      @       @      8@      @      @      @      @      6@       @      4@      6@      C@      @      &@      @      @      &@              $@              @              &@       @      @                                      &@      @      4@      @     �D@      1@      @     �L@      @      b@              B@             @a@      *@      $@      �?      @     �D@      @      T@     �D@     �^@      (@      4@      1@      �?     �C@      @     @]@              >@             @]@      @      $@      �?      �?     �C@       @     �O@      9@     @[@      @      5@               @      2@              <@              @              5@      $@                      @       @      �?      1@      0@      ,@      @      3@      @      "@     �E@              J@              &@              3@      @       @              @      5@      �?      4@      9@      >@      @                              @                                               @      �?      �?                      @                      @      �?              3@      @      "@     �B@              J@              &@              1@      @      �?              @      0@      �?      4@      6@      =@      @      ,@      @      @     �B@              ;@              $@              *@      @                      @      *@      �?      ,@      0@      4@      @      @      @       @                      9@              �?              @              �?                      @              @      @      "@             �o@     �Z@     �R@     �l@      >@     @o@       @      d@      D@     �o@     �U@      ?@      ;@     �G@     `d@      H@     @n@      i@     `l@      P@     �X@     �L@     �I@     �Z@      3@     �R@       @     �W@      =@     @Y@     �E@      4@      2@      9@      R@      5@     �[@     �W@     �U@      5@      J@      A@      ;@     �Q@      "@      L@      @      I@      @     @R@      6@      *@      "@      &@      D@      &@     �Q@     �C@      M@      (@      I@      8@      3@     @P@      "@      J@      @     �G@      @      R@      6@      $@      @      $@     �C@       @      Q@      C@     �K@      &@       @      $@       @      @              @              @              �?              @      @      �?      �?      @      @      �?      @      �?     �G@      7@      8@      B@      $@      2@       @     �F@      7@      <@      5@      @      "@      ,@      @@      $@      D@     �K@      =@      "@      .@      "@      &@      6@      @      @      �?      @@      ,@      "@      "@      @              @      @      @      (@      9@       @      @      @@      ,@      *@      ,@      @      &@      �?      *@      "@      3@      (@      @      "@      @      9@      @      <@      >@      5@      @     `c@     �H@      7@     �^@      &@      f@             @P@      &@      c@      F@      &@      "@      6@     �V@      ;@     ``@     �Z@     �a@     �E@     @R@      ;@      .@     �R@      @      ^@              =@      @      V@      4@      @      @      @     �L@      $@     �V@     �O@     �O@      =@      7@      4@      @      F@       @      P@              ,@       @      G@      .@      @      @      �?      ;@      @     �I@      F@     �F@      3@      I@      @       @      ?@       @      L@              .@      @      E@      @                       @      >@      @      D@      3@      2@      $@     �T@      6@       @      H@      @      L@              B@      @      P@      8@      @      @      3@      A@      1@      D@      F@     @S@      ,@      C@      (@      @      6@      @      ?@              7@       @     �D@      @      @               @      ,@      @      .@      ,@      A@      @      F@      $@      @      :@      @      9@              *@       @      7@      2@      �?      @      1@      4@      &@      9@      >@     �E@      "@�t�bub�       hhubehhub.