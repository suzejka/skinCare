���&      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C0                                           �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K�
node_count�KU�nodes�hhK ��h��R�(KKU��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B�                             �2@q� ���?s            �\@                           @��_�q�?1            �H@                           @����D�?%            �B@                            @�d��0�?             >@                           �?      �?              @������������������������       �                      @       
                     �?�8��8��?             @       	                    �?      �?              @������������������������       �                     �?������������������������       �                     �?                          �1@      �?             @������������������������       �                     @������������������������       �                     �?                           @���7�?             6@������������������������       �                     ,@                             @      �?              @������������������������       �r�q��?             @������������������������       �                      @                          �1@������?             @                          �0@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �z�G�z�?             @                           @r�q��?             (@                           �?"pc�
�?             &@                            �?      �?             @������������������������       �      �?              @������������������������       �                      @                            �?؇���X�?             @������������������������       �                     @������������������������       �      �?             @������������������������       �                     �?!       L                    @�Ra����?B            �P@"       ?                    @��?��?4             J@#       4                    �?���/<��?#            �A@$       )                     �?~�Q���?             3@%       &                    �?�8��8��?             @������������������������       �      �?              @'       (                    �?      �?             @������������������������       �      �?              @������������������������       �                      @*       -                      @�]�`��?             *@+       ,                    �?�q�q�?             @������������������������       �      �?              @������������������������       �                     �?.       1                    @{�G�z�?
             $@/       0                    �?      �?             @������������������������       �                      @������������������������       �      �?              @2       3                    �?�8��8��?             @������������������������       �      �?              @������������������������       �      �?             @5       >                      @     ��?             0@6       =                    �?d}h���?             ,@7       :                     �?      �?             (@8       9                    6@r�q��?             @������������������������       �                     @������������������������       ��q�q�?             @;       <                    @�q�q�?             @������������������������       �      �?              @������������������������       �      �?             @������������������������       �                      @������������������������       �      �?              @@       E                    �?=[y���?             1@A       D                    @      �?             @B       C                   �5@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @F       G                   �3@�	j*D�?             *@������������������������       �                     �?H       K                    @      �?             (@I       J                    �?z�G�z�?
             $@������������������������       ��q�q�?             @������������������������       �                     @������������������������       �      �?              @M       P                    �?������?             ,@N       O                     �?���Q��?             @������������������������       �                      @������������������������       �                     @Q       T                    @�q�q�?	             "@R       S                     �?      �?              @������������������������       �      �?              @������������������������       ��q�q�?             @������������������������       �                     �?�t�b�values�hhK ��h��R�(KKUKK��hV�B�        *@      :@      &@      ;@      ;@      &@               @      �?      8@      .@      �?              @      �?      8@      @      �?              @              8@      �?                      @              @      �?                       @                                               @              @      �?                      �?                      �?                      �?                                                                      �?                      �?              @                                              @                              �?                                              �?              5@                                              ,@                              �?              @                              �?              @                                               @                              �?      �?              @      �?                      �?                      �?                      �?                                                                      �?              �?                      @                       @                      $@                       @                      "@                      �?                      @                      �?                      �?                                               @                      �?                      @                                              @                      �?                      @                                              �?              *@      2@      $@      @      (@      $@      *@      .@      @      @      (@       @      *@      $@      @       @      @       @      �?      @      @       @      @       @               @              �?      @                      �?              �?                              �?                      @                      �?                      �?                                               @              �?      @      @      �?               @                      �?                       @                      �?                      �?                                              �?      �?      @      @      �?                      �?      @                                               @                                      �?      �?                                               @      @      �?                              �?              �?                              �?      @                              (@      @      �?                              &@      @                                      "@      @                                      @      �?                                      @                                               @      �?                                      @       @                                      �?      �?                                      @      �?                                       @                                              �?              �?                                      @       @      �?      "@                      �?       @      �?                              �?              �?                                              �?                              �?                                                       @                                      @                      "@                      �?                                              @                      "@                       @                       @                       @                      @                                              @                      �?                      �?                      @      @                       @                      @                       @                                               @                      @                                      @                              @              @                              @              �?                              �?               @                              @                                              �?�t�bub�_sklearn_version��1.1.0�ub.