��%     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.1.2�ub�n_estimators�Kd�estimator_params�(�	criterion��	max_depth��min_samples_split��min_samples_leaf��min_weight_fraction_leaf��max_features��max_leaf_nodes��min_impurity_decrease��random_state��	ccp_alpha�t��	bootstrap���	oob_score���n_jobs�NhN�verbose�K �
warm_start��hN�max_samples�NhhhKhKhKhG        h�log2�hNhG        hG        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h5�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C�                                                                	       
                                                               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhKhKhKhG        hh.hNhJ���3hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��h>�f8�����R�(KhBNNNJ����J����K t�b�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFh2�scalar���h>�i8�����R�(KhBNNNJ����J����K t�bC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hK�
node_count�Ks�nodes�h4h7K ��h9��R�(KKs��h>�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hwhZK ��hxhZK��hyhZK��hzh>�f8�����R�(KhBNNNJ����J����K t�bK��h{h�K ��h|hZK(��h}h�K0��uK8KKt�b�B(         <                     @�md&��?�	           ��@                           @$U̚S�?�           F�@                          �2@�9�KL��?N            �@                           @�؁�m��?�            0q@                            �?��A1Z�?�            �i@                            �?�R;����?q            �e@������������������������       ���\m��?G            �Z@������������������������       �n�1�^�?*             Q@	       
                    �?�>U��p�?             ?@������������������������       ��q�q�?             (@������������������������       ����.�?
             3@                          �0@p!`�j��?*            �Q@������������������������       �@�0�!��?
             1@                           �?�fXf��?             �J@������������������������       ��n�MJ��?             E@������������������������       ����k���?             &@                          �8@bQ�@���?�           Ԑ@                           �?�4>�?�           ؄@                           �?�a@]�a�?           �{@������������������������       �d6�M�?�             k@������������������������       ������?�             l@                           �?p�=@`&�?�             l@������������������������       �����tI�?;            �Z@������������������������       �ܶm۶m�?I            �]@                          �@@��h1��?           �y@                           �?L����?�            �w@������������������������       ���r���?:            �X@������������������������       ��t�r�?�            �q@                          �A@�9+�Q�?             =@������������������������       �Iє�?             1@������������������������       �r�q��?             (@        -                    �?�� ���?o           l�@!       &                    @����6�?-           �~@"       #                   �0@F]t�e�?�             v@������������������������       �     ��?             @@$       %                    @�����	�?�             t@������������������������       �Za���L�?y            @h@������������������������       �L�_�B��?L            �_@'       *                     �?�������?V             a@(       )                   �1@�7Ry��?=            @X@������������������������       �
ףp=
�?             4@������������������������       ���p�h��?2            @S@+       ,                   �3@�"c�I�?            �C@������������������������       ���1G���?             *@������������������������       �ݾ�z�<�?             :@.       5                   �3@�C9�r�?B           ��@/       2                   �1@�T M�?�            0t@0       1                    �?�|�j��?V             ^@������������������������       �(�=z��?-            �P@������������������������       �mq�$X�?)             K@3       4                    �?}���&�?�            `i@������������������������       �g\�5�?	             *@������������������������       ���2C��?{            �g@6       9                    @t4]2��?h           ��@7       8                    �?�ORD��?�             w@������������������������       ��H�����?s            @g@������������������������       �1�K36��?~             g@:       ;                   �7@ߏ0P��?w            �g@������������������������       ��vaWN�??            �W@������������������������       �UUUUU��?8             X@=       \                    @�l���?�           ��@>       M                   �7@V�����?           h�@?       F                    �?�&%j�?t           ��@@       C                    @���޺�?�            �o@A       B                   �5@�T����?�             i@������������������������       �.�:�wM�?n             d@������������������������       ����(\��?             D@D       E                    �?�θ�?             J@������������������������       ��ˠT�?             6@������������������������       ��������?             >@G       J                    �?�H����?�             t@H       I                    @)� �f��?S            @`@������������������������       ��,o��?            �D@������������������������       ���sv��?7            @V@K       L                    �?r�qO�?�             h@������������������������       ��8��8��?             8@������������������������       �� � �?r             e@N       U                   �9@���_K*�?�            �p@O       R                    �?�������?E             ]@P       Q                    @��s���?             K@������������������������       ���Q��?             D@������������������������       ��Cc}�?             ,@S       T                    �?��6�/�?'             O@������������������������       ��q-�T�?!             J@������������������������       ��G�z��?             $@V       Y                    �?Y���O��?d            @c@W       X                   �=@θ	j�?E             Z@������������������������       ��k�vC�?,            �P@������������������������       ���X�<�?            �B@Z       [                    @F��_��?             I@������������������������       �������?            �A@������������������������       �<+	���?             .@]       j                    �?p�~fz��?�            �u@^       e                    @���JT�?U             a@_       b                    �?V>�� =�?9            @W@`       a                    8@���.�?             3@������������������������       ���(\���?             $@������������������������       ��<ݚ�?             "@c       d                   �5@��._�?,            �R@������������������������       ��o�����?             ;@������������������������       ���O"�?            �G@f       i                    @���k���?             F@g       h                    @������?             =@������������������������       ��������?	             1@������������������������       ��8��8��?             (@������������������������       �hE#߼�?             .@k       l                   �0@>�Q��?|             j@������������������������       �&�q-�?             *@m       p                    �?c����?t            `h@n       o                    @I���?            �F@������������������������       ����%�?             :@������������������������       �P7�Z�?             3@q       r                   �6@d�2����?Y            �b@������������������������       �S4%t6V�?2            �U@������������������������       �ğӯZ��?'            �O@�t�b�values�h4h7K ��h9��R�(KKsKK��h��BHD       0{@      Q@     �u@     �A@     @Q@      =@     �W@     ��@     ��@      O@     �U@     �b@     ��@     ~@      ,@      P@      J@     ``@     @Q@     `t@     �A@      l@      9@      F@      &@      P@     �z@     �|@      C@     �N@      Y@     pz@     �r@      @      C@      :@     @S@      E@      e@      ,@      a@      .@      @@      &@      F@     �]@     �i@      7@     �E@     �L@     `j@     �c@      �?      3@      *@      H@     �A@     �I@      �?      4@                              @      O@      N@      @      @      @     �E@      5@                              �?       @     �D@      �?      *@                              @     �K@      @@      �?      @      @     �A@      0@                              �?              C@      �?      @                               @      G@      ?@      �?      @       @      ?@      ,@                              �?              7@      �?      @                               @      >@      (@      �?       @      �?      7@      @                              �?              .@              �?                                      0@      3@              �?      �?       @      @                                              @              "@                               @      "@      �?                      �?      @       @                                               @                                                       @      �?                              �?                                                      �?              "@                               @      �?                              �?      @       @                                              $@              @                                      @      <@       @              �?       @      @                                       @                                                              @      ,@                                                                                      $@              @                                      @      ,@       @              �?       @      @                                       @       @              @                                      @      @       @              �?      @      @                                       @       @                                                              @                               @                                                     @]@      *@      ]@      .@      @@      &@      D@     �L@      b@      4@      D@     �J@      e@      a@      �?      3@      *@     �G@     �@@     @V@      @     @P@      @      &@      �?      1@      G@      \@      @      7@      :@      ^@      W@              @      @      8@      .@     �N@      @     �G@              @              $@      ?@     �H@      @      5@      4@     �S@      R@              @      @      0@      .@      ?@      �?      &@                              @      (@      >@      �?      "@      @     �L@     �A@                      �?      @      &@      >@       @      B@              @              @      3@      3@      @      (@      *@      5@     �B@              @      @      &@      @      <@      @      2@      @      @      �?      @      .@     �O@      @       @      @      E@      4@              �?               @               @       @      $@               @               @       @      @@       @              @      9@      &@                              @              4@      �?       @      @      @      �?      @      *@      ?@      �?       @       @      1@      "@              �?               @              <@      @     �I@      (@      5@      $@      7@      &@     �@@      *@      1@      ;@      H@     �F@      �?      *@      "@      7@      2@      :@      @     �H@      "@      5@      $@      7@      &@      >@       @      0@      3@      G@      F@      �?      *@       @      7@      1@      ,@      �?      @       @      @       @      &@       @      .@              �?       @      (@      $@      �?       @      �?      $@              (@      @      F@      @      ,@       @      (@      "@      .@       @      .@      1@      A@      A@              &@      @      *@      1@       @               @      @                                      @      @      �?       @       @      �?                      �?              �?                      �?      @                                      �?      �?      �?      @       @                                              �?       @              �?                                               @      @              �?              �?                      �?                     �c@      5@     @V@      $@      (@              4@     Ps@     �o@      .@      2@     �E@     �j@     �a@       @      3@      *@      =@      @     �E@      @      3@              �?              @     �b@     �Z@       @      $@      *@     �P@     �J@              @       @      @       @      5@      @      0@                               @     @^@      T@      �?      "@      (@      K@      9@              �?               @      �?      �?                                                      =@      �?                              �?                                                      4@      @      0@                               @      W@     �S@      �?      "@      (@     �J@      9@              �?               @      �?      3@      @      ,@                               @      E@      D@      �?      @      "@     �@@      3@              �?               @      �?      �?      @       @                                      I@     �C@               @      @      4@      @                                              6@              @              �?              �?      ;@      :@      �?      �?      �?      *@      <@              @       @      @      �?      "@              @              �?              �?      5@      4@      �?      �?      �?      *@      4@              @       @      �?              @                                                      @      @                      �?                                              �?              @              @              �?              �?      .@      *@      �?      �?              *@      4@              @       @                      *@                                                      @      @                                       @              @               @      �?       @                                                      @       @                                      @                                              &@                                                      @      @                                       @              @               @      �?     �\@      ,@     �Q@      $@      &@              1@      d@     `b@      *@       @      >@      b@      V@       @      (@      &@      8@      @     �E@      @      1@      @                      @     @W@      Q@      @      �?      @     �I@      5@              �?       @      @              0@       @       @                              @      ;@      >@                      @      <@      @                              �?               @                                              @      3@      7@                              $@      @                                               @       @       @                                       @      @                      @      2@      @                              �?              ;@       @      .@      @                      @     �P@      C@      @      �?       @      7@      ,@              �?       @       @              @                                                      �?      @                                       @                                              5@       @      .@      @                      @     @P@      A@      @      �?       @      7@      (@              �?       @       @              R@      $@     �J@      @      &@              &@      Q@     �S@      "@      @      8@     �W@     �P@       @      &@      "@      5@      @      G@      "@      9@      @      @              @      J@     �N@      @      �?       @     @R@     �H@       @      @      @      $@      �?      =@      @      2@              @              @     �@@     �B@       @      �?      @      7@      6@              �?      @      @              1@      @      @      @      @               @      3@      8@      @              @      I@      ;@       @      @              @      �?      :@      �?      <@      @      @              @      0@      2@      @      @      0@      5@      2@              @      @      &@      @      ,@              @               @               @      $@      *@              @      &@      1@       @              �?      �?      @       @      (@      �?      5@      @       @              @      @      @      @      @      @      @      $@              @      @       @       @     @[@     �@@     �^@      $@      9@      2@      >@     �Y@     �a@      8@      9@     �I@     �e@     �f@      &@      :@      :@      K@      ;@     �T@      3@     �T@      "@      2@      ,@      ,@     �U@     �\@      1@      2@      B@     �]@     �]@      @      2@      3@     �@@      4@     �P@       @     �L@      �?      $@      @      @      U@     @U@      $@      &@      3@      X@     @P@      �?      $@      $@      7@      @     �A@      @      6@              "@      @      @      =@      A@      @       @      $@     �A@      A@      �?      @      @      &@      @      @@      @      *@              "@      @              0@      8@      @       @      $@      <@      =@      �?      @      @      &@      @      9@       @      @              @      @              ,@      5@       @       @      $@      <@      9@               @      @      &@       @      @       @      @              @      �?               @      @      �?                              @      �?      �?      @              @      @              "@                              @      *@      $@                              @      @               @                               @               @                                      @       @                               @       @                                              �?              @                              @      @       @                              @      @               @                              @@      @     �A@      �?      �?      �?      @     �K@     �I@      @      "@      "@     �N@      ?@              @      @      (@              "@              ,@                      �?      �?     �A@      5@              @      @      9@      $@              @       @       @              @              @                              �?      $@       @               @      �?      *@      �?              �?              �?              @               @                      �?              9@      3@              �?      @      (@      "@               @       @      �?              7@      @      5@      �?      �?              @      4@      >@      @      @      @      B@      5@               @       @      $@               @      �?      @              �?                              �?       @      @              @      �?                                              5@      @      0@      �?                      @      4@      =@      @      �?      @      >@      4@               @       @      $@              0@      &@      9@       @       @      "@      @      @      >@      @      @      1@      7@      K@      @       @      "@      $@      ,@      @      @      @      �?       @       @      @       @      2@                       @      "@      C@       @       @      @      @               @      @       @              �?                       @      @                      @      @      9@                      �?      @               @      �?                      �?                       @      @                      @      @      5@                              @                      @       @                                              @                                      @                      �?                      @       @      @      �?      �?       @      @              (@                      @      @      *@       @       @      @                      @       @      @              �?       @      @              $@                      @      @      "@               @      @                                              �?                                       @                              �?      @       @                                      $@      @      3@      @      @      @      @      �?      (@      @      @      "@      ,@      0@       @      @      @      @      ,@      @      �?      1@      @      @      @      @              @      @      @      @       @      @      �?      @      @       @      *@      @      �?      (@       @      @      �?      @              @      @              @      @      @              @      �?       @      @      �?              @      @              @                              �?      @      �?       @      �?      �?       @       @              @      @      @       @                      @              �?       @      @              @      @      "@      �?      �?              @      �?      @      @      �?                      @                      @      @              @      @       @      �?      �?              @      �?                      �?                                      �?      @                               @      @                                              :@      ,@      D@      �?      @      @      0@      0@      :@      @      @      .@      K@     �O@      @       @      @      5@      @      (@      @      $@               @       @      @      @      .@       @       @      @      =@      9@              @      @      @      �?      @      @      @               @       @       @      @      (@      �?              @      7@      6@              @      �?       @      �?                                                       @              �?                      �?      "@      @                               @      �?                                                                      �?                      �?      @      �?                               @                                                               @                                              @       @                                      �?      @      @      @               @       @              @      &@      �?              @      ,@      3@              @      �?                      �?               @                                      �?      @      �?              �?      &@       @              @                              @      @      @               @       @               @      @                       @      @      1@                      �?                      @       @      @                              @       @      @      �?       @              @      @               @      @      @              @      �?      @                                       @       @               @               @       @                      @      @               @      �?      @                                       @       @                                                              @      @              @              �?                                                               @               @       @                                                      �?                                      @              �?      �?                      @      �?               @               @              ,@      "@      >@      �?      @       @      &@      &@      &@      @      @      &@      9@      C@      @       @       @      ,@      @                      �?               @                       @                                               @                                              ,@      "@      =@      �?      @       @      &@      @      &@      @      @      &@      9@      B@      @       @       @      ,@      @      "@              @                                              @      @      @      @       @      "@                       @      @       @      @              �?                                              �?      @      @      �?      �?      @                       @      @       @      @               @                                              @                      @      �?      @                                              @      "@      :@      �?      @       @      &@      @      @       @       @      @      7@      ;@      @       @              &@      @      @      @      @      �?              �?      @      �?      @       @              @      5@      4@                               @              �?      @      3@              @      �?      @       @                       @      �?       @      @      @       @              @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�؇ohG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         <                    �?��Fs|��?�	           ��@                          �4@�s����?|           4�@                            @�U���a�?'           ��@                           �?��r�OF�?�           ��@                          �2@U#54c�?�            �p@                           @�����?j            `d@������������������������       �~ឮ:c�?W            �`@������������������������       �;U��j�?             =@	       
                     �?O|��?=            �Z@������������������������       �(����?+            �R@������������������������       �c�=��?             ?@                            �?����?�            0v@                           @G�m���?�            �n@������������������������       ��YK�'��?�            �h@������������������������       ��/�<n�?#            �F@                           @���9�t�?=            �[@������������������������       �      �?             0@������������������������       ��o6A��?5            �W@                           �?�t]Ec��?�             p@                          �2@0�����?             B@������������������������       ������?             6@������������������������       ��Cc}�?             ,@                          �1@�������?�            �k@                           �?�@���?.            �R@������������������������       ���x��?             7@������������������������       ��s�n_�?             J@                           �?`��W�?W            `b@������������������������       ����E�?            �J@������������������������       ��bj*R[�?9            �W@       -                   �9@�݋PB��?U           ،@       &                    �?#��tO�?�           p�@        #                     �?"q[[e�?�            �i@!       "                   �7@_{fI���?N            @_@������������������������       ����{/��?:            �W@������������������������       ��?�P�a�?             >@$       %                   �6@����/��?7            �T@������������������������       ��0�!��?             A@������������������������       ��q�q��?             H@'       *                    @}��R��?           �y@(       )                    @ܩ����?4             W@������������������������       ������j�?             H@������������������������       ���#��Z�?             F@+       ,                    @�`��i�?�            0t@������������������������       ��灐��?w            �f@������������������������       �����1J�?c            �a@.       5                   �<@w��g�?�            �r@/       2                    �?Q����?s            �e@0       1                   �;@;�;��?%             J@������������������������       �T]���b�?            �@@������������������������       ��	"P7��?             3@3       4                   �:@`�e\y�?N            �^@������������������������       ����0�G�?"             K@������������������������       ��}2��?,             Q@6       9                     �?��]��?O            �_@7       8                    @hJ,���?,             Q@������������������������       �*f��N�?            �C@������������������������       �΃�\W�?             =@:       ;                    �?=d��*�?#            �M@������������������������       �n�����?             .@������������������������       ���eP*L�?             F@=       Z                    �?�����?%           x�@>       K                    @0�<�D�?X           ��@?       F                    �?����v�?k           ��@@       C                   �2@7wGͶ�?�            �l@A       B                     �?��Z���?            �D@������������������������       �>
ףp=�?             4@������������������������       ��u]�u]�?             5@D       E                   �3@�c�P��?h            `g@������������������������       �@��Z��?
             7@������������������������       �n�2��?^            �d@G       H                   �0@��5�?�            �v@������������������������       ���!pc�?             &@I       J                   �5@�N~5�?�            0v@������������������������       ��]3����?l            �e@������������������������       �U$?����?u            �f@L       S                    �?�`�i�?�             x@M       P                   �5@��n����?R            @`@N       O                    @Э�*��?%             M@������������������������       �UUUUUU�?             (@������������������������       �#8̺�8�?             G@Q       R                     @��8��8�?-             R@������������������������       ��q�q�?             �I@������������������������       �~VC�1��?             5@T       W                    @    @O�?�             p@U       V                     �?Hrw���?+             O@������������������������       �      �?              @������������������������       �uk~X��?$             K@X       Y                     �?�
�/�$�?p            @h@������������������������       �R�AI-��?(             O@������������������������       �S��a`��?H            �`@[       d                   �5@��M�-L�?�           ��@\       c                    @E�u�I�?�           H�@]       `                    @l��u:�?�           ��@^       _                   �0@VUߘ��?4           �~@������������������������       �     �?!             P@������������������������       ����[�?           �z@a       b                   �3@�^B{	m�?a             b@������������������������       ���X��?A            �W@������������������������       �m���?             �H@������������������������       ��g���e�?             &@e       l                    @�"����?2           �}@f       i                    @mr�)E��?�            �t@g       h                   �9@<����?�            `q@������������������������       �1�=�M�?i            �d@������������������������       ����˸�?G            �[@j       k                    @�a9���?!            �I@������������������������       �pƵHP�?	             *@������������������������       �J�w�"w�?             C@m       p                     @�a�r���?a            �b@n       o                    @59�� �?H            �[@������������������������       �VF�ߎ�?5            @S@������������������������       ��ߋm��?            �@@q       r                    @{�G�z�?             D@������������������������       �N�7��?             =@������������������������       �F]t�E�?             &@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       0}@     @T@     @v@      ?@      R@     �@@     @R@     �@     �@     �L@      R@     `d@     ��@     @y@      ,@     �P@     �L@     �`@      J@      n@      A@     �a@      @      7@      @      ?@      v@     �s@      .@     �@@      P@     �q@     `d@       @      4@      2@      H@      ,@     @]@       @      G@       @       @       @      @     0p@     �c@      @      $@      5@     `b@     �R@              @              7@       @     �R@      �?      5@       @      �?              @     `k@     �_@       @      @      &@     �W@     �J@              �?              @              7@              "@                                     @\@      H@              @      @     �B@      :@                                              0@              @                                     �T@      ?@              @       @      *@      (@                                              (@               @                                     �R@      7@              @              *@      @                                              @               @                                      @       @                       @              @                                              @              @                                      ?@      1@              @      @      8@      ,@                                              @              @                                      0@      "@              @      @      7@      $@                                               @              �?                                      .@       @                              �?      @                                             �I@      �?      (@       @      �?              @     �Z@     �S@       @      �?      @      M@      ;@              �?              @             �C@      �?      @       @      �?              @      N@      O@       @      �?       @      F@      .@              �?              @              @@      �?      @       @      �?              @     �K@      K@              �?       @      :@      (@              �?              @              @               @                                      @       @       @                      2@      @                                              (@              @                                      G@      0@                       @      ,@      (@                              @              @              �?                                               @                              @      @                              @              "@              @                                      G@      ,@                       @      $@      "@                                             �E@      �?      9@              �?       @      @      D@     �@@       @      @      $@      J@      6@              @              0@       @      &@              �?                                       @      @      �?              �?      @      @                              @              @              �?                                      @      @      �?              �?       @                                      @              @                                                      @       @                              �?      @                                              @@      �?      8@              �?       @      @      @@      <@      �?      @      "@     �H@      3@              @              *@       @      2@              @                                      .@      1@      �?                      .@      @                                              @              �?                                      @      $@                              @       @                                              ,@              @                                      (@      @      �?                      (@      �?                                              ,@      �?      2@              �?       @      @      1@      &@              @      "@      A@      0@              @              *@       @      @      �?       @              �?       @              �?      @                              1@      @                              @              @              $@                              @      0@       @              @      "@      1@      $@              @              @       @     �^@      @@      X@      @      5@      @      8@     @W@     �c@      &@      7@     �E@     �`@      V@       @      0@      2@      9@      (@     �S@       @      Q@      �?       @      @      .@     �S@     @]@      @      ,@      A@      V@      O@              $@      (@      .@      @      ?@      @      3@              �?              @      4@     �I@      �?      @       @      C@      .@              @              @      �?      .@              .@                              @      (@      A@      �?      @      @      <@       @                              �?      �?      &@              (@                               @      @      9@      �?      @      @      ;@      @                                              @              @                               @      @      "@                              �?      @                              �?      �?      0@      @      @              �?                       @      1@                      @      $@      @              @              @               @       @       @                                      @       @                              @      @               @              �?              ,@      @       @              �?                       @      "@                      @      @      �?               @               @              H@      �?     �H@      �?      @      @      &@     �M@     �P@      @      &@      :@      I@     �G@              @      (@      &@       @      @              0@                               @      2@      @      �?              @      .@       @              @      @      @               @              .@                               @      �?      �?                      @      "@      @              @       @      �?              @              �?                                      1@      @      �?                      @      @                      @      @             �E@      �?     �@@      �?      @      @      "@     �D@      N@      @      &@      3@     �A@     �C@               @      @      @       @      6@              :@      �?      @      @      @      ,@      9@               @      1@      3@      :@               @      @               @      5@      �?      @              �?              @      ;@     �A@      @      @       @      0@      *@                      �?      @              F@      8@      <@       @      *@              "@      ,@     �C@      @      "@      "@     �F@      :@       @      @      @      $@      "@      9@      1@      $@       @      @              @      ,@      6@      �?      @      @      ?@      2@              �?      @       @      @      (@      @      @      �?                              @      $@              @      @      @      @                      �?      �?              @              @      �?                              @       @                       @      @      @                      �?      �?              @      @                                                       @              @      �?      �?      @                                              *@      ,@      @      �?      @              @      &@      (@      �?      @              ;@      &@              �?      @      @      @      "@      @      @              �?               @      �?      @                              .@      @              �?       @      �?      @      @       @      @      �?       @              @      $@      @      �?      @              (@       @                      �?      @              3@      @      2@              $@              @              1@      @      @      @      ,@       @       @      @       @       @      @      (@      @       @              @              �?              0@               @      @       @      @              �?               @      @      "@      @      �?               @                              @               @      @              @              �?              �?      �?      @              @              �?              �?              $@                               @      �?                              �?      @      @              $@              @               @              �?      @      �?              (@      @       @      @       @               @      @              �?                                                              �?               @                       @                              @              "@              @               @              �?      @                      @      @       @       @       @               @     `l@     �G@     �j@      :@     �H@      ;@      E@     �k@     �r@      E@     �C@     �X@     �s@      n@      (@     �G@     �C@     �U@      C@     @Y@      ;@     @Z@      ,@      <@      6@      3@     �C@      ]@      >@      A@      M@      _@      a@       @      8@      =@     �D@      8@     �Q@      4@      L@       @      3@      *@       @      9@     @U@      $@      3@      ?@     �T@      T@      @      ,@      1@      <@      @      2@      @      3@              @      @      @      1@      B@              @      $@     �A@     �B@              @       @      "@      @      @               @                                      $@       @              �?       @      &@      �?                                              @               @                                      @      @                      �?      @      �?                                              �?                                                      @      @              �?      �?       @                                                      (@      @      1@              @      @      @      @      <@              @       @      8@      B@              @       @      "@      @                       @                                              @               @                      @              @                      @      (@      @      .@              @      @      @      @      7@              @       @      8@      @@                       @      "@       @      J@      ,@     �B@       @      *@      $@      @       @     �H@      $@      (@      5@     �G@     �E@      @      @      "@      3@              "@              �?                                      �?                                                                                             �E@      ,@      B@       @      *@      $@      @      @     �H@      $@      (@      5@     �G@     �E@      @      @      "@      3@             �@@      @      *@       @      @               @       @     �@@       @      $@      @      >@      4@              �?              @              $@      "@      7@      @       @      $@      �?      @      0@       @       @      ,@      1@      7@      @      @      "@      (@              ?@      @     �H@      @      "@      "@      &@      ,@      ?@      4@      .@      ;@      E@     �L@      @      $@      (@      *@      3@      6@              (@              @              @      @      ,@      "@       @      @      1@      .@              @      @      @      @      "@              @                              �?      �?      *@      @              @      @      @                      @      @      @      @                                              �?                                       @               @                      �?               @      @              @                                      �?      *@      @              @      @       @                       @      @      �?      *@              @              @              @      @      �?       @       @      �?      ,@      &@              @       @      �?      @      @              @              �?              @       @      �?       @       @      �?      $@       @              @      �?      �?      @      @              �?              @                       @                                      @      @                      �?                      "@      @     �B@      @      @      "@      @      "@      1@      &@      *@      5@      9@      E@      @      @      @      "@      (@      �?      �?      @                       @       @      �?      @      @      @       @       @      ,@               @      @       @      @                       @                                      �?      �?                                                      �?              �?       @      �?      �?      @                       @       @              @      @      @       @       @      ,@              �?      @      �?      @       @      @      @@      @      @      @      @       @      (@      @       @      3@      7@      <@      @      @              @      @       @              &@      @       @      @      �?              @       @      @       @      @      @               @                      @      @      @      5@      @       @      @      @       @      @      @      �?      &@      2@      6@      @      @              @       @     �_@      4@     @[@      (@      5@      @      7@     �f@     �f@      (@      @     �D@      h@      Z@      @      7@      $@     �F@      ,@     �Q@      @      L@      @       @      �?      (@     @c@     �^@      @      @      *@     @[@      I@              &@      @      *@      &@     �Q@      @      L@      @       @      �?      &@     @c@     �^@      @      @      *@     �Z@     �E@              &@      @      *@      &@      I@       @      G@       @       @      �?      @     �`@     �W@      @      @      $@      V@      A@              @      @      @      @      @                                                      <@      .@                              .@                                                      F@       @      G@       @       @      �?      @     @Z@      T@      @      @      $@     @R@      A@              @      @      @      @      5@       @      $@      �?      @              @      5@      ;@                      @      2@      "@              @       @      @      @      *@       @       @      �?                      @      0@      6@                       @       @      @              @       @      @               @               @              @              @      @      @                      �?      $@      @                              �?      @                                                      �?                                              @      @                                             �K@      0@     �J@      "@      *@      @      &@      <@      M@      "@       @      <@     �T@      K@      @      (@      @      @@      @      D@      $@      8@      @      $@      @      @      9@      H@      @       @      5@     �N@      A@      @      $@       @      1@       @      B@      @      5@      @      $@      @      @      ,@      D@      @       @      4@      E@      A@      @      "@       @      1@       @      8@      @      (@      @      @      �?      @      $@      B@      �?       @      @      =@      1@              @              @       @      (@      �?      "@       @      @      @      �?      @      @      @              ,@      *@      1@      @      @       @      (@              @      @      @                                      &@       @                      �?      3@                      �?                                                                                      @      @                              @                                                      @      @      @                                      @      @                      �?      0@                      �?                              .@      @      =@      @      @              @      @      $@      @              @      6@      4@      �?       @      @      .@      �?      *@      @      :@      @      �?              @      @      @      @              @      (@      1@               @      @       @      �?      $@      @      2@      @      �?              �?       @       @      @              @      @      1@               @      �?      @              @               @                               @      �?       @                      @      "@                               @       @      �?       @      @      @               @               @              @                      �?      $@      @      �?                      @               @       @      �?               @              �?              @                      �?      $@       @                               @                      �?       @                              �?                                                      �?      �?                      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJIp�ohG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKuhnh4h7K ��h9��R�(KKu��hu�B�         <                   �2@�ԓ1��?�	           ��@                           �?LV�`��?�           ��@                           @>�O*�2�?;           �~@                            �?�A�E|��?�            @j@                           �?��I�_�?F             [@                           �?贁N�?*             N@������������������������       ����ލL�?             ;@������������������������       ��"��?            �@@	       
                    @r�qG�?             H@������������������������       �s�	U���?             A@������������������������       �                     ,@                           �?�κ��~�?@            �Y@                          �0@���bo�?(            �Q@������������������������       �<+	���?             .@������������������������       �j�V���?!            �K@                           @     �?             @@������������������������       �9��8���?             8@������������������������       �      �?              @                            @yJ"9�?�            `q@                           @�k�	���?�            `m@                          �1@&	\�O�?r            �f@������������������������       �4S�1�[�?I            �\@������������������������       �.C�d�K�?)            �P@                            �?/
k��?&             K@������������������������       ���(\���?             D@������������������������       ���>4և�?
             ,@                           @Us�k���?            �E@                            @�������?             >@������������������������       ��1G����?	             *@������������������������       ��hJ,��?             1@������������������������       �����W�?             *@        /                    @%�wށ��?X            �@!       (                    @��LE?�?�            �z@"       %                     �?��ǆM�?�            `p@#       $                    �?�&T����?*             Q@������������������������       ���"e���?             B@������������������������       �     P�?             @@&       '                    �?*=8-��?t            @h@������������������������       ��
�GN�?2             V@������������������������       �l<�1�'�?B            �Z@)       ,                     �?-Xm� �?`            �d@*       +                   �1@T���,c�?0            @U@������������������������       �8��d�?$             O@������������������������       �36�v[�?             7@-       .                    @y[��G��?0            �S@������������������������       �HP�s�?             9@������������������������       ��X;�U��?             K@0       7                    @��E���?Z            @c@1       4                    @E%]}��?F            @\@2       3                     �?�	��?+            �P@������������������������       �9��8���?             8@������������������������       �`*�s��?             E@5       6                     �? Q�"T��?            �G@������������������������       �{�/��>�?
             1@������������������������       �؂-؂-�?             >@8       9                     �?(x��:�?            �D@������������������������       �؉�؉��?             *@:       ;                    �?������?             <@������������������������       �F]t�E�?             &@������������������������       �躍`3�?             1@=       Z                    @���Gs��?-           :�@>       M                   �=@IPS!��?G            �@?       F                    �?b�����?�           d�@@       C                    @��T�)D�?�           8�@A       B                     �?����G�?
           �y@������������������������       �����?F            �\@������������������������       ��ѷQC�?�            �r@D       E                     @4�ݦ��?�            �m@������������������������       ����h�*�?`             c@������������������������       �ՙ/,�?8             U@G       J                   �5@������?:           ��@H       I                    @��H9n�?�            0s@������������������������       �`�_A
J�?�            `q@������������������������       ����Kϟ�?             =@K       L                     @8VSK�?n           ��@������������������������       ��c)����?�            �t@������������������������       �%_L
�8�?�            �j@N       S                    �?�&Ͼ�?k            �d@O       P                   �>@     ��?(             P@������������������������       �
ףp=
�?             4@Q       R                     �?ޏ��k��?             F@������������������������       ������?             3@������������������������       ��A`��"�?             9@T       W                   �>@j�«R~�?C            �Y@U       V                    �?f��S�?            �@@������������������������       ������H�?             "@������������������������       ��q�q�?             8@X       Y                     @�j U��?,            �Q@������������������������       ��������?             E@������������������������       �������?             <@[       j                   �:@2�$X�?�           t�@\       c                    �?ǵ�O�?~           ؏@]       `                    @3��Od{�?>           0�@^       _                     �?@Xc,$��?V            @b@������������������������       �{�G�z�?             D@������������������������       �
�rk�B�?>            �Z@a       b                    @`(L�
�?�            @w@������������������������       �     V�?M             `@������������������������       �hg�h��?�            �n@d       g                   �3@��G��o�?@           P@e       f                     �?�����
�?5            @U@������������������������       �      �?             0@������������������������       ���L��s�?(            @Q@h       i                    @ʃg\[�?            z@������������������������       �˕6�#��?C            �[@������������������������       ��� �tY�?�             s@k       r                    @%
|u�?h            @d@l       o                     �?#hT�?X             a@m       n                    @8�q_��?            �@@������������������������       ��������?             1@������������������������       �      �?             0@p       q                    @�"AM�h�?@             Z@������������������������       ����=A�?             C@������������������������       �l�����?$            �P@s       t                    @ݵ�|г�?             9@������������������������       �ףp=
��?             $@������������������������       ��|�j��?
             .@�t�bh�h4h7K ��h9��R�(KKuKK��h��BxE       0}@     @Q@     �t@     �@@     @S@      3@     @Q@     x�@     ��@     �S@      W@     `c@     8�@     �z@      &@      O@      Q@     @^@     �L@     `a@      ,@      N@      �?      @               @     �p@     �m@      &@      @      5@     �d@      V@              "@       @      2@      @     �M@      @      3@                              @      d@     �^@      @      �?      @     �Q@      :@              @              @              A@       @      @                              @     �H@      O@       @      �?      �?      B@      @              @              @              (@       @      @                                      ?@     �F@              �?              &@      �?                               @              @       @       @                                      5@      1@              �?              $@                                                      @               @                                      *@      @                              @                                                      @       @                                               @      *@              �?              @                                                      @              �?                                      $@      <@                              �?      �?                               @              @              �?                                      $@      ,@                              �?      �?                               @                                                                              ,@                                                                                      6@              @                              @      2@      1@       @              �?      9@       @              @              @              (@              @                              @      0@       @      �?              �?      .@       @              @              @              @              �?                                      @                                      @                                                      @               @                              @      &@       @      �?              �?      (@       @              @              @              $@                                                       @      "@      �?                      $@                                                      "@                                                       @      @                              "@                                                      �?                                                              @      �?                      �?                                                      9@      @      *@                                      \@     �N@       @              @      A@      7@                                              2@      @      @                                     �W@      M@       @              @      ;@      7@                                              "@       @      �?                                      U@      F@                              4@      5@                                              @       @      �?                                     �O@      6@                              ,@      @                                               @                                                      5@      6@                              @      0@                                              "@      @      @                                      &@      ,@       @              @      @       @                                              @      @      �?                                      $@       @       @              @      @      �?                                              @               @                                      �?      @                                      �?                                              @              "@                                      1@      @                              @                                                      @              @                                      ,@       @                              �?                                                      �?              @                                      @      �?                              �?                                                      @              �?                                      $@      �?                                                                                      �?               @                                      @      �?                              @                                                      T@      @     �D@      �?      @              @     @[@     �\@      @      @      1@     �W@      O@              @       @      &@      @     �P@      @      9@      �?      @              @     �U@      T@      @      @      "@     �S@     �C@              @       @      @       @      D@      @      $@      �?      @              @     �A@     �I@      @      @       @     �N@      9@              �?       @      @               @                                              �?      ,@      $@      @      �?              9@      @                                              @                                                      @      @              �?              0@      �?                                              �?                                              �?      "@      @      @                      "@      @                                              @@      @      $@      �?      @              @      5@     �D@       @      @       @      B@      3@              �?       @      @              6@      �?       @              @               @      $@      7@       @               @      ,@      @                                              $@      @       @      �?       @              �?      &@      2@              @      @      6@      *@              �?       @      @              ;@       @      .@                              �?     �I@      =@                      �?      2@      ,@              @              �?       @      7@       @                                              4@      5@                      �?      @       @               @              �?              0@      �?                                              1@      3@                      �?      @                                      �?              @      �?                                              @       @                                       @               @                              @              .@                              �?      ?@       @                              &@      @              �?                       @       @               @                                      @      �?                              @                                                       @              @                              �?      8@      @                              @      @              �?                       @      *@              0@                                      7@      A@       @       @       @      .@      7@              �?      @      @      @      "@              $@                                      0@      <@                      @      &@      1@              �?      @      @      @      @               @                                      @      3@                              @      0@                              @      @      @              @                                      �?      @                              �?      @                                              �?               @                                       @      (@                              @      (@                              @      @      @               @                                      *@      "@                      @      @      �?              �?      @      @              @                                                      @                                      �?      �?              �?      @       @                               @                                      $@      "@                      @      @                                      �?              @              @                                      @      @       @       @      @      @      @                                      �?                       @                                      @                              @              @                                      �?      @              @                                      @      @       @       @              @      @                                              @               @                                                       @                      @                                                                       @                                      @      @               @              �?      @                                             �t@     �K@      q@      @@     �Q@      3@     �N@     p@     �x@      Q@     @U@     �`@     0|@     `u@      &@     �J@      N@     �Y@      I@     �f@      C@      f@      .@     �I@      2@     �D@     @S@     �i@      F@     �M@      W@      p@     �j@      @     �D@     �C@     �Q@      D@     �d@      A@     �d@      "@     �E@      *@      D@     @S@      i@      @@     �F@      R@     �n@      i@      �?      A@      9@     �M@     �@@     �P@      .@      Q@      @      "@      @      &@     �D@     �Z@      @      5@      <@     �`@     �T@              &@      (@      5@      &@     �C@       @     �C@      �?      @      @       @      ?@     �S@       @      *@      1@     @Q@      N@               @      "@      .@      @      "@              @      �?      @              @      @      ;@              @      @      3@      1@               @       @      $@      �?      >@       @      A@                      @      @      :@      J@       @       @      (@      I@     �E@              @      @      @      @      ;@      @      =@       @      @      @      @      $@      ;@      �?       @      &@      P@      6@              @      @      @      @      6@      @      2@              @              �?      @      1@      �?      @              F@      1@              @              @       @      @      �?      &@       @       @      @       @      @      $@               @      &@      4@      @                      @       @       @      Y@      3@     �X@      @      A@      @      =@      B@     �W@      =@      8@      F@     �\@     �]@      �?      7@      *@      C@      6@     �H@      @     �B@              @      �?       @      .@      I@      @      @      2@     �A@      F@              @      @      1@      �?      G@      @      ?@              @      �?      @      .@     �H@      @      @      0@      >@     �D@              @      @      0@      �?      @              @              �?              @              �?       @               @      @      @                              �?             �I@      (@     �N@      @      >@      @      5@      5@     �F@      8@      2@      :@     �S@     �R@      �?      3@      @      5@      5@      B@      "@     �A@              *@      @      &@      2@      :@      (@      (@      *@     �P@      B@      �?      (@      @      ,@      "@      .@      @      :@      @      1@      @      $@      @      3@      (@      @      *@      (@      C@              @      @      @      (@      .@      @      &@      @       @      @      �?              @      (@      ,@      4@      "@      ,@      @      @      ,@      &@      @      ,@      �?      �?              @              �?              @       @      @      @      @      @      �?      @      @      @      �?       @                                                                              @      @      �?                      �?              �?              @      �?      �?              @              �?              @       @      @              @      @      �?       @      @       @      �?      �?      �?                                      �?              @       @      @                      @                       @       @              @              �?              @                                                              @      @      �?       @      @              �?      �?      @      $@      @      @      @                              $@      @      ,@       @       @      @      @      "@       @      @              @      @      �?      @       @                                      @              �?      @              @      �?      @                      @      �?              �?                                                              �?       @                      �?                                      @      �?       @       @                                      @                       @              @              @              �?              @      @       @      @                              $@       @      ,@      �?      @      @      �?       @      @      @                      @      @       @       @                              @      �?      "@      �?       @              �?      @      @              �?                       @              �?                              @      �?      @               @      @               @              @     `b@      1@     �W@      1@      4@      �?      4@     �f@     �g@      8@      :@      E@     `h@      `@      @      (@      5@     �@@      $@     @`@      *@     �R@      0@      2@              0@     �e@     �e@      ,@      1@      >@     �e@     �Z@      @      &@      .@      9@      "@     @P@      @      ?@      @      @              @     �\@     �W@      (@      $@      (@     �T@      L@               @      @      &@       @      =@              @      @       @              @      3@      8@      @              @      8@      .@                      �?      @       @      @              @      @                      �?      @      $@       @               @      @      @                                              9@              �?               @              @      0@      ,@       @              @      5@       @                      �?      @       @      B@      @      9@              @                     �W@     �Q@       @      $@      @     �M@     �D@               @      @      @               @              2@                                      D@      1@       @      @      @      6@      $@                      @      �?              <@      @      @              @                     �K@      K@      @      @      @     �B@      ?@               @       @      @             @P@      "@     �E@      *@      *@              "@     �M@      T@       @      @      2@     �V@     �I@      @      "@      "@      ,@      @       @      �?      @      @                       @      @      @@               @      @      @      &@               @       @               @      �?      �?      �?       @                              @       @               @              @                                                      @              @      @                       @      @      >@                      @      �?      &@               @       @               @     �L@       @     �C@       @      *@              @      J@      H@       @      @      .@     �U@      D@      @      @      @      ,@      @      (@              0@       @      @                      8@      @               @      @      4@      *@              �?               @      �?     �F@       @      7@      @      "@              @      <@     �D@       @      @      "@     �P@      ;@      @      @      @      (@      @      1@      @      5@      �?       @      �?      @      @      ,@      $@      "@      (@      6@      5@      �?      �?      @       @      �?      (@      @      1@      �?              �?      �?      @      (@      $@      "@      (@      6@      *@      �?      �?      @       @              @      �?      �?                              �?       @       @      @              @              @                      @       @              @      �?      �?                              �?      �?       @      @                              �?                               @              �?                                                      �?               @              @              @                      @                       @      @      0@      �?              �?              @      $@      @      "@      "@      6@       @      �?      �?      �?      @               @      �?      @                                              @       @      @       @      ,@      �?      �?              �?      �?              @       @      (@      �?              �?              @      @      �?      @      @       @      @              �?              @              @              @               @              @               @                                       @                                      �?      @                               @                                                                      @                                               @              @                              @               @                                      @                                      �?�t�bub�R"     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJb8khG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKohnh4h7K ��h9��R�(KKo��hu�BH         >                   �5@?���=��?�	           ��@                           @�R��W��?U           �@                           �?��Qw��?�            �@                          �2@�t3ޝD�?�           ��@                            @K�q�#�?�            �u@                           �?�ߎ ��?{            �g@������������������������       �6g*͸�?1            �Q@������������������������       �mT$�0�?J            �]@	       
                    �?B	Y����?b            �c@������������������������       �c���?-            �S@������������������������       �ڽ���?5            @S@                            �?Vn�*�?           �{@                           �?������?O            ``@������������������������       ���K�[��?              O@������������������������       ��*2S�?/            @Q@                            @�`�n6q�?�            �s@������������������������       ����NV��?D            @Z@������������������������       ��o5;/Z�?�            `j@                            �?˒����?�             s@                           @��j+���??             Y@                           @��İ2�?/            @S@������������������������       ��b�b�?%             O@������������������������       ��A��S�?
             .@������������������������       �t���?             7@                          �3@L���(`�?�            �i@                            @��$�5�?S            �`@������������������������       ��b����?2             U@������������������������       ���{�P�?!             I@                           �?�\$����?1            �Q@������������������������       �?,R�n�?             B@������������������������       ���¤�h�?             A@        /                     @�%�N���?�           �@!       (                    �?VjѡL�?           @�@"       %                   �0@���� �?           @|@#       $                    �?z~Riv�?&             M@������������������������       �l��[B��?             =@������������������������       ���Ϧ���?             =@&       '                    @e�a����?�            �x@������������������������       �az��?�            �q@������������������������       ������?G             \@)       ,                    @5�1	4�?�            @z@*       +                    �?���>j7�?�            �q@������������������������       �ʫ֮f��?=            @X@������������������������       �F���v��?s            �g@-       .                     �?�sEi�?O            �`@������������������������       ���WV��?!             J@������������������������       ��� ����?.            @T@0       7                    �?@�M���?�            �j@1       4                   �2@���>4��?5             U@2       3                    �?u���?             E@������������������������       ��袋.��?             6@������������������������       ���Q��?             4@5       6                   �4@��|�`��?             E@������������������������       ��*�{72�?             ;@������������������������       �؂-؂-�?             .@8       ;                   �3@     M�?Q             `@9       :                    �?��|���?8             V@������������������������       �r�O��?            �C@������������������������       ��lB1rq�?             �H@<       =                    �?�(\����?             D@������������������������       ��9����?             6@������������������������       ��)O�?	             2@?       ^                   �<@�M�]�?I           �@@       O                    �?��f��+�?z           ̕@A       H                   �6@L�XTU��?~           ��@B       E                    @�6����?V            �_@C       D                    �?s��?c�?,            @P@������������������������       ����x�?             7@������������������������       ���?"md�?             E@F       G                    @�c�1��?*             O@������������������������       �-)���?             =@������������������������       ���3cڟ�?            �@@I       L                    @nD;��?(           @}@J       K                   �7@��`����?�            �v@������������������������       ��F.��9�?=            @Y@������������������������       �ρ�M��?�            �p@M       N                    @'�J�?A            �Y@������������������������       ���!pc�?             &@������������������������       ��i#��?;            �V@P       W                   �8@M�O�t�?�            �@Q       T                    �?�	&��9�?*           @}@R       S                     �?Pm.<b)�?�            �i@������������������������       ��յ� c�?,            @P@������������������������       ��;J�L��?Y            �a@U       V                    @�L�����?�            `p@������������������������       �I��͸(�?q            �e@������������������������       �{v�X�?4             V@X       [                    @H��|O]�?�            �t@Y       Z                    �?�&���`�?~            �g@������������������������       �Ĝ�-�?             =@������������������������       ��v�b^m�?j            @d@\       ]                     @L!vѩ�?T            �a@������������������������       �nb����?:            �W@������������������������       ����,d!�?             G@_       j                    @�L��Ԫ�?�             u@`       e                    @vpJ����?�            pr@a       d                   �A@��4\5��?�            `m@b       c                   �@@Q�J7���?�            �k@������������������������       �t���P��?}             i@������������������������       ��(\����?             4@������������������������       �d}h���?             ,@f       i                    @�a�r���?*             N@g       h                    �?�a��d�?             �G@������������������������       �����X�?	             ,@������������������������       ����%��?            �@@������������������������       �ݾ�z�<�?
             *@k       l                    �?�C�_�;�?            �E@������������������������       �x9/���?             ,@m       n                   @@@��`���?             =@������������������������       �n,�Ra�?	             6@������������������������       �������?             @�t�bh�h4h7K ��h9��R�(KKoKK��h��B�A       @~@     �W@     �u@      D@      S@      7@     �W@     Ȁ@     8�@      O@      Y@     `d@     (�@     0y@      $@      K@     �I@     ``@     �H@     �s@      5@     �c@      (@      3@      @      ?@     �z@     �y@      .@      @@      R@     �u@      i@              2@      *@      P@      *@      f@      ,@     �V@      @      ,@      @      2@     �`@     `h@      &@      4@      E@     �f@      ^@              &@      "@     �D@      @     @`@      (@     �Q@       @      (@       @      *@     �U@     �\@      $@      3@      A@      a@      W@              &@       @      @@      @      F@      @      >@              @              @     �I@      J@      @      "@      0@      Q@      =@              @      @      1@      @      >@              ,@              �?               @      ?@     �B@       @       @      "@     �E@      *@                               @      @      1@              @                                      1@      0@                      @      &@      @                                              *@              &@              �?               @      ,@      5@       @       @      @      @@      "@                               @      @      ,@      @      0@               @              @      4@      .@       @      @      @      9@      0@              @      @      .@              @      �?      @                              @      .@      @       @              @      0@       @              @               @              $@      @      &@               @                      @      "@              @      �?      "@       @              �?      @      @             �U@      @      D@       @      "@       @       @      B@     �O@      @      $@      2@     @Q@     �O@              @      @      .@      @      9@       @      &@       @                      �?      @      7@              @       @      @@      2@                              @              1@              @                                      @      "@              @              5@      �?                                               @       @      @       @                      �?      �?      ,@              �?       @      &@      1@                              @             �N@      @      =@              "@       @      @      >@      D@      @      @      0@     �B@     �F@              @      @      $@      @      8@              "@              @              @      4@      $@              @      @      @      *@              @              @      �?     �B@      @      4@              @       @      @      $@      >@      @      �?      &@      ?@      @@               @      @      @       @     �G@       @      5@       @       @      @      @     �G@      T@      �?      �?       @      G@      <@                      �?      "@      �?      2@              @       @                              3@      A@      �?               @      "@      @                              @      �?      0@              @                                      1@      4@      �?               @      "@      @                              @      �?      $@              @                                      *@      2@                       @      "@      @                              �?      �?      @                                                      @       @      �?                                                               @               @                       @                               @      ,@                                      �?                               @              =@       @      2@               @      @      @      <@      G@              �?      @     �B@      6@                      �?      @              8@              *@               @                      7@      :@              �?      @      7@      *@                      �?      @              ,@              "@                                      0@      3@                      �?      (@      $@                      �?       @              $@              @               @                      @      @              �?      @      &@      @                              �?              @       @      @                      @      @      @      4@                      �?      ,@      "@                              �?               @       @                              @               @      *@                      �?      @      @                              �?              @              @                              @      @      @                              "@       @                                             �a@      @     �P@       @      @              *@     0r@     �k@      @      (@      >@     �d@      T@              @      @      7@      @      [@      @     �D@       @      @              &@     �o@     �g@       @      @      8@     �`@     �O@              @      @      0@      @      D@       @      1@      �?      �?              @      c@     �Z@       @              &@     @T@      >@                               @               @               @                                     �@@      $@                              &@                                                       @               @                                      4@       @                              @                                                                                                              *@       @                               @                                                      C@       @      .@      �?      �?              @     �]@      X@       @              &@     �Q@      >@                               @              4@      �?      (@      �?                      @     @X@      P@      �?              @     �I@      5@                               @              2@      �?      @              �?                      6@      @@      �?              @      3@      "@                                              Q@      @      8@      �?      @              @      Y@     �T@              @      *@      K@     �@@              @      @      ,@      @     �F@      �?      3@                                      V@     �L@              @      @      >@      5@              �?               @      @      @              @                                      C@      <@               @       @       @      @                                              C@      �?      ,@                                      I@      =@              @      @      6@      ,@              �?               @      @      7@      @      @      �?      @              @      (@      9@              �?      @      8@      (@              @      @      @              @      @      �?      �?      �?              @      @      &@                       @      (@      @                              @              3@              @              @                      @      ,@              �?      @      (@       @              @      @      @              A@      �?      9@      @                       @     �C@      @@       @      @      @      ?@      1@               @      �?      @       @      *@              (@      @                      �?      "@      @               @       @      1@      (@                              @      �?      @              (@                                      @      @               @      �?      "@                                                       @              @                                      @      @                              @                                                      @              @                                       @                       @      �?      @                                                      @                      @                      �?      @      �?                      �?       @      (@                              @      �?      �?                      @                      �?       @      �?                      �?      @      "@                                      �?      @                                                       @                                      �?      @                              @              5@      �?      *@       @                      �?      >@      9@       @      @      @      ,@      @               @      �?      @      �?      $@              $@       @                              8@      8@              @      �?      @      @               @              �?      �?      "@              @                                      $@      @              @              �?      @                                              �?              @       @                              ,@      2@                      �?      @      �?               @              �?      �?      &@      �?      @                              �?      @      �?       @              @       @      �?                      �?       @              @                                              �?      @               @                      @      �?                      �?       @               @      �?      @                                              �?                      @       @                                                     �d@     �R@     `g@      <@     �L@      2@      P@      \@      i@     �G@      Q@     �V@      m@     `i@      $@      B@      C@     �P@      B@     �a@      N@     �b@      7@      B@      $@      I@      Z@     �d@      A@     �E@     �P@     �j@     �c@      @      <@      <@     �I@      ;@     @P@      <@      Q@      @      @      @      7@      I@     @Z@      "@      *@      ,@      X@      Q@              @      "@      .@      @       @      �?      3@              @      �?       @      .@     �@@                              9@      ,@                       @      @              @      �?      3@              @      �?       @      @      $@                              ,@      @                      �?                      �?               @                                      �?      @                              @      �?                                              @      �?      &@              @      �?       @      @      @                              @      @                      �?                      @                                                      &@      7@                              &@       @                      �?      @                                                                      $@      (@                               @      @                      �?                      @                                                      �?      &@                              "@      @                              @             �L@      ;@     �H@      @      @      @      5@     �A@      R@      "@      *@      ,@     �Q@      K@              @      @      &@      @     �G@      3@     �E@      @      @      @      5@      2@      J@      @      "@      ,@     �N@     �C@              @      @      $@      @      3@      @      @              @               @      "@      *@      @      @      @      3@      "@                      �?      �?              <@      (@     �B@      @      �?      @      3@      "@     �C@              @      $@      E@      >@              @      @      "@      @      $@       @      @       @                              1@      4@      @      @              $@      .@               @              �?      �?      �?              �?                                      "@                                                                                              "@       @      @       @                               @      4@      @      @              $@      .@               @              �?      �?      S@      @@      T@      0@      =@      @      ;@      K@      O@      9@      >@     �J@     �]@     �V@      @      5@      3@      B@      4@      O@      ,@      G@      @      0@       @      @     �D@      C@      "@      6@      <@     �L@      O@      @      $@      "@      9@      $@      4@       @      3@      �?      $@       @      �?      *@      (@      @      4@      $@      6@      B@               @      @      "@      "@      ,@       @      @      �?      �?                      @       @      @      @      @      &@      @                      @      �?      @      @      @      (@              "@       @      �?       @      $@       @      0@      @      &@      @@               @      @       @      @      E@      @      ;@      @      @              @      <@      :@      @       @      2@     �A@      :@      @       @       @      0@      �?     �@@      @      0@      @                      @      1@      2@      @       @      @      ?@      7@              @      �?      "@              "@      �?      &@      @      @              �?      &@       @                      *@      @      @      @      @      �?      @      �?      ,@      2@      A@      "@      *@      @      5@      *@      8@      0@       @      9@     �N@      =@      �?      &@      $@      &@      $@      "@      $@      7@      @      &@      @      @      $@      1@      &@      @      &@      A@      @      �?      @      $@       @      @      @                              @      �?              @      �?              �?      �?      $@      �?                      �?       @              @      $@      7@      @       @      @      @      @      0@      &@       @      $@      8@      @      �?      @      "@      @      @      @       @      &@       @       @              0@      @      @      @      @      ,@      ;@      6@               @              @      @      @      @      @       @      �?              @      �?      @      @      @      "@      9@      ,@              @               @      @              @      @              �?              *@       @      @                      @       @       @               @              �?              8@      ,@     �C@      @      5@       @      ,@       @     �@@      *@      9@      8@      2@      F@      @       @      $@      0@      "@      4@      ,@      ;@      @      5@       @      ,@       @      ;@      *@      9@      7@      2@      ?@      @       @      $@      *@      @      (@      ,@      2@      @      0@      @      *@       @      8@      (@      9@      5@      0@      3@      @      @      @      @      @      (@      *@      0@      @      "@      @      *@       @      8@      (@      6@      5@      0@      3@      @      @      @      @      @      (@      *@      .@      @      "@      @      *@       @      8@      (@      5@      *@      *@      3@       @      @      @      @      @                      �?                                                              �?       @      @               @       @               @      �?              �?       @              @      �?                                      @                                                                       @              "@       @      @       @      �?              @      �?               @       @      (@      �?       @      @      @      �?      @              "@       @      @       @      �?              @                       @              "@      �?       @      @      @      �?      �?              @               @              �?              @                                                               @      �?               @              @       @       @       @                                               @              "@      �?       @      �?      @      �?      @                              �?                                      �?                       @      @                              �?              @              (@                                              @                      �?              *@                              @      @                                                                      @                                      @                              �?      @      @              (@                                                                      �?              "@                               @      �?                      &@                                                                                      "@                               @              @              �?                                                                      �?                                                      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ\�yhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         >                   �4@���块�?�	           ��@                          �1@ 'fdC�?i           ��@                           @��_H��?�           H�@                           @z������?�             p@                            �?���P�8�?�            �h@                            �?T�Ɣ��?N            �[@������������������������       ���Hx��?-             R@������������������������       �,r�|��?!             C@	       
                    @�zv�X�?=             V@������������������������       �     ��?#             H@������������������������       �ffffff�?             D@                           @�Q����?'             N@                             @*Uf����?            �C@������������������������       �VUUUUU�?             8@������������������������       ��.�?�P�?             .@                             @�&%�ݒ�?             5@������������������������       ���8��8�?             (@������������������������       �h/�����?             "@                           @J�fF��?�            pt@                          �0@VI��?�            �o@                           @"�%��?4            �T@������������������������       �s����?             >@������������������������       ���/�y�?            �J@                           @;`�&��?k             e@������������������������       ���w���?S            ``@������������������������       ��+r�|�?             C@                           @�@���?4            �R@                            �?�������?+             N@������������������������       �     @�?             0@������������������������       �t�E]t�?             F@������������������������       �VUUUUU�?	             .@        /                   �3@�������?�           ��@!       (                    �?��'f��?�           ��@"       %                     @/�d�<�?�            @x@#       $                     �?�� }J��?�            �p@������������������������       �#8_&�J�?v             g@������������������������       ��"���?3            @T@&       '                    �?�0l��?K            �^@������������������������       ���8��8�?             B@������������������������       ����)k��?2            �U@)       ,                     @f�&���?�            @y@*       +                    �?���f�?�            �p@������������������������       �d�I�R�?;            �W@������������������������       ����tp��?o            �e@-       .                   �2@���]�M�?T            �`@������������������������       �3O�x�?1            �S@������������������������       ��|f59�?#            �K@0       7                    �?�6Wr���?�            �x@1       4                    �?��@W�s�?j            �f@2       3                     �?{�ӉF��?'            �Q@������������������������       �V-��?             9@������������������������       �h����?             G@5       6                     �?v�c�9v�?C            �[@������������������������       �}댯�t�?$             O@������������������������       ��q�q\�?             H@8       ;                    �?��^B{	�?�             k@9       :                     �?�̿0�=�?             ?@������������������������       �.y0��k�?             *@������������������������       ����Hx�?
             2@<       =                    @m�{,U�?v             g@������������������������       �rª���?D            @Z@������������������������       �>
ףp}�?2             T@?       X                    �?���s*�?I           ��@@       I                    �?Z�\��j�?P           ��@A       H                   �=@G9sJ�?�            �r@B       E                     �?�@%�PW�?�            �q@C       D                   �5@�#��9�?.            @S@������������������������       �Ǻ����?             9@������������������������       �s�n_Y��?              J@F       G                   �6@TD� ���?�            �i@������������������������       ��;�64�?8            �V@������������������������       �/�H=��?M            �\@������������������������       �n�����?	             .@J       Q                   �9@�� ���?�           @�@K       N                    @��b�>J�?           |@L       M                    @���i)�?�             p@������������������������       �-)�?�             m@������������������������       ���?��?             :@O       P                   �7@���V-C�?u            �g@������������������������       ��gB����?U            @a@������������������������       ��
Yg��?             �J@R       U                    @�k�y��?�            �h@S       T                     @���nN�?            �C@������������������������       �'��}��?             ;@������������������������       ���8��8�?
             (@V       W                   @@@��(\�r�?j             d@������������������������       �٫~Q$��?[             a@������������������������       �      �?             8@Y       h                     @3Q��b�?�           ��@Z       a                    �?H	�2R�?           @�@[       ^                     �?#����?�            �o@\       ]                   �5@x]��g��?o            @f@������������������������       ��GN��?             F@������������������������       ��q�"��?V            �`@_       `                    @���yZ�?+            �R@������������������������       ����1u��?              M@������������������������       �ZZZZZZ�?             1@b       e                    @5���d�?�           X�@c       d                     �?�ϥ���?�            �t@������������������������       �
���x�?p            �c@������������������������       �v�X��?n             f@f       g                    @>�����?�            �o@������������������������       ����&��?C            @Z@������������������������       ����]4�?_            `b@i       p                    @!j���;�?�             v@j       m                    @z	N��'�?�            �o@k       l                   �7@�/�$�?�             i@������������������������       ��nx��^�?1            �S@������������������������       �*=6�9��?S            @^@n       o                   �8@~4��?            �J@������������������������       �     ��?             @@������������������������       ��ܤ��?
             5@q       t                    @��`}�^�?>            @Y@r       s                    �?f~w��?)            �Q@������������������������       �����k�?             G@������������������������       �46<�R�?             9@u       v                    �?�P�a�r�?             >@������������������������       �
ףp=
�?             4@������������������������       �>
ףp=�?             $@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       @}@      T@     Pu@     �@@      U@     �B@     @Q@     ��@     Ђ@     @P@      S@     �b@     ��@     0}@      .@      R@      L@     �_@      G@     �j@      2@     @^@      "@      *@       @      "@     �x@     �t@      .@      8@     �M@     0t@     �b@              5@       @     �F@      $@      S@      @      .@               @               @     @g@     �^@      @      @      3@     �Y@      A@                              @      @     �D@      �?      $@              �?              �?     �J@      G@      @      @      $@     �M@      3@                              @      @      B@      �?      @              �?              �?      I@      9@       @      @      "@     �H@      &@                               @       @      0@              �?              �?              �?      B@      .@              @      @      9@      @                               @       @      $@                                              �?      8@      @              @       @      5@      @                              �?      �?      @              �?              �?                      (@      "@                       @      @      �?                              �?      �?      4@      �?      @                                      ,@      $@       @      �?      @      8@      @                                              "@      �?                                              @      @       @      �?      @      3@       @                                              &@              @                                       @      @                       @      @      @                                              @              @                                      @      5@      @              �?      $@       @                              @      �?      @              �?                                       @      3@                              @      @                              @               @                                                       @      .@                              @       @                                              �?              �?                                              @                              @       @                              @               @              @                                      �?       @      @              �?      @      @                                      �?      �?                                                      �?       @      @              �?      @                                              �?      �?              @                                                                                      @                                             �A@      @      @              �?              �?     �`@     @S@              �?      "@     �E@      .@                               @              5@      @      @                              �?     �[@     �N@              �?      @      @@      $@                               @               @                                                     �J@      (@                              @       @                              �?              @                                                      *@       @                              @                                                      @                                                      D@      @                              �?       @                              �?              *@      @      @                              �?      M@     �H@              �?      @      9@       @                              �?              &@       @       @                              �?      I@     �D@              �?      @      *@      @                                               @      @       @                                       @       @                              (@       @                              �?              ,@              �?              �?                      6@      0@                      @      &@      @                                              $@              �?              �?                      3@      "@                      @      $@      @                                                                                                      @      @                       @       @      �?                                              $@              �?              �?                      ,@      @                      @       @      @                                              @                                                      @      @                              �?                                                     @a@      (@     �Z@      "@      &@       @      @     �j@     �j@      $@      3@      D@     �k@     �\@              5@       @      C@      @     @U@       @     �S@      @      @              @     �c@     @c@      "@      $@      >@     �^@     �R@              *@      @      :@      @      D@       @      <@      @                       @     @W@     �R@      @      @      3@      M@      F@               @              *@      �?     �@@       @      1@      @                             @R@     �K@      @       @      (@      B@      7@                              @              3@       @      $@      @                              F@      @@      @       @      $@      ?@      6@                              @              ,@              @                                      =@      7@                       @      @      �?                                              @              &@                               @      4@      3@              �?      @      6@      5@               @              "@      �?      @              "@                                       @      �?                              @      @                              @               @               @                               @      2@      2@              �?      @      1@      ,@               @               @      �?     �F@      @      I@      @      @              @     �O@      T@      @      @      &@      P@      ?@              &@      @      *@      @      @@       @     �@@      �?      �?               @      L@      M@       @      @      @     �A@      6@              @      @      @              @              7@      �?                              "@      2@       @      @      @      ,@      $@              �?              @              9@       @      $@              �?               @     �G@      D@                       @      5@      (@              @      @      @              *@      @      1@      @      @              �?      @      6@      �?      @      @      =@      "@              @      �?      @      @      "@      @      @       @                      �?      @      .@              @      @      5@      @                              @      @      @      �?      (@      �?      @                      �?      @      �?      �?       @       @      @              @      �?       @             �J@      @      <@       @      @       @       @     �L@      M@      �?      "@      $@     �X@      D@               @       @      (@      @      7@       @      @              @       @      �?      >@      A@              @             �J@      (@              @              @               @                              �?       @              *@      &@                              ?@      @                              �?               @                                                      �?      �?                              2@       @                              �?              @                              �?       @              (@      $@                              *@       @                                              .@       @      @               @              �?      1@      7@              @              6@       @              @              @               @              �?               @              �?       @      3@              @              &@      @              @                              @       @      @                                      "@      @              @              &@      @                              @              >@       @      5@       @      @              �?      ;@      8@      �?       @      $@      G@      <@              @       @       @      @      @               @                                               @      �?              @      (@       @                       @              �?                                                                      �?                              &@                                              �?      @               @                                              �?      �?              @      �?       @                       @                      9@       @      3@       @      @              �?      ;@      6@               @      @      A@      :@              @               @       @      .@       @      .@                              �?      ,@      $@              �?      @      ,@      6@                              @      �?      $@              @       @      @                      *@      (@              �?      �?      4@      @              @              @      �?     �o@      O@     �k@      8@     �Q@     �A@      N@     �`@     �p@      I@      J@     �V@     �p@     �s@      .@     �I@      H@     �T@      B@     �_@      0@     @V@      @      8@       @      1@     �T@     `c@      .@      3@      A@     `c@     ``@       @      2@      6@      3@      ,@      I@      "@      6@      �?      @               @      .@     �R@      @      @      @      H@      D@       @      @      @      @      �?     �F@      "@      6@      �?      @               @      .@     �R@      @      @      @     �D@      C@       @      @      @      @      �?      (@              �?      �?       @              �?       @      =@      @      �?              *@       @                      @                      @                                                      �?      @              �?              &@       @                                              @              �?      �?       @              �?      �?      8@      @                       @      @                      @                     �@@      "@      5@               @              �?      *@     �F@       @      @      @      <@      >@       @      @              @      �?      (@      @      "@                                       @      4@              �?       @      3@      (@              �?               @      �?      5@      @      (@               @              �?      @      9@       @      @      @      "@      2@       @       @              @              @                                                              �?                              @       @                                              S@      @     �P@      @      4@       @      .@     �P@      T@      $@      ,@      <@     �Z@     �V@              .@      2@      ,@      *@      J@      �?     �D@      �?      @       @      (@     �O@      O@       @      "@      6@      Q@     �R@              @      *@      @       @      B@              ?@      �?      @       @      &@      .@      9@               @      .@      G@     �G@              @      $@      �?       @      <@              <@      �?      @       @      &@      .@      8@              @      (@      C@     �G@              @      "@               @       @              @                                              �?              �?      @       @                              �?      �?              0@      �?      $@              @              �?      H@     �B@       @      �?      @      6@      ;@              @      @      @              .@              @              @                      B@      @@      @      �?      @      2@      (@                      @      @              �?      �?      @                              �?      (@      @       @              @      @      .@              @                              8@      @      :@      @      *@              @      @      2@       @      @      @     �C@      1@               @      @      "@      &@      @              (@              @                      �?               @              @       @       @              @              @      �?       @              $@               @                      �?               @              @      �?      �?               @              @              @               @              �?                                                              �?      �?              @                      �?      3@      @      ,@      @      $@              @      @      2@              @      @     �B@      .@              @      @      @      $@      .@      @      *@      @      @               @      @      2@              @       @      B@      $@               @      @      @      @      @              �?              @              �?                               @      �?      �?      @              �?       @              @      `@      G@     ``@      3@     �G@     �@@     �E@      I@      \@     �A@     �@@     �L@      ]@     `g@      *@     �@@      :@     �O@      6@     @Y@      7@     �X@      *@     �@@      ,@      @@      E@     @T@      >@      ;@     �B@     �V@     @]@       @      ;@      2@      E@      (@      ?@      @      9@      �?      @       @      "@      2@      E@      "@       @      @      5@      F@       @      @      �?      "@      @      7@      �?      2@              @      @       @      0@      8@      "@      @      @      ,@      B@       @      @      �?       @               @              �?                      @      @      @      &@              �?              �?      "@                              �?              .@      �?      1@              @              @      (@      *@      "@      @      @      *@      ;@       @      @      �?      @               @      @      @      �?      �?      @      �?       @      2@              @      @      @       @               @              �?      @      @      �?      @      �?      �?      @               @      0@              @      @      @      @              �?                              @      @                                      �?               @                                      �?              �?              �?      @     �Q@      0@     @R@      (@      =@      @      7@      8@     �C@      5@      3@      ?@     �Q@     @R@              6@      1@     �@@      "@      =@       @     �A@      @      6@      @      3@      *@      6@      .@      .@      (@      :@      G@              3@      (@      7@      @      $@      @      4@      @      "@      @       @      @      &@      @      @      @      *@      :@              "@      @       @      @      3@       @      .@       @      *@              &@       @      &@      (@       @       @      *@      4@              $@      @      .@      @     �D@       @      C@      @      @              @      &@      1@      @      @      3@      F@      ;@              @      @      $@      @      1@      @      9@      @      �?              �?      "@      @      @              $@      $@      (@                       @      @              8@      @      *@      �?      @              @       @      ,@      @      @      "@      A@      .@              @      @      @      @      ;@      7@     �@@      @      ,@      3@      &@       @      ?@      @      @      4@      9@     �Q@      &@      @       @      5@      $@      3@      3@      .@       @      *@      2@      @      @      >@      @      @      ,@      4@     �H@      @      @      @      "@       @      @      .@      .@       @      $@      *@      @      @      5@      @      @      *@      .@     �E@       @      @      @       @       @      @      &@       @       @      @       @       @      @      "@      �?              @      @      @              @      @      @               @      @      @              @      @       @       @      (@      @      @      $@      &@      B@       @       @      @      @       @      *@      @                      @      @       @      �?      "@                      �?      @      @       @              �?      �?              $@       @                                              �?      @                              @      @       @                                      @       @                      @      @       @               @                      �?              �?                      �?      �?               @      @      2@      @      �?      �?      @       @      �?      �?       @      @      @      5@      @              �?      (@       @      @       @      $@              �?                      �?              �?       @      @      @      3@      @              �?      &@       @      @      �?      "@              �?                                      �?       @      @      �?       @      @              �?      @       @              �?      �?                                      �?                                      @      &@                              @              @       @       @      @              �?      @      �?      �?                      �?               @      �?                      �?               @       @      @      @              �?      @      �?                              �?              �?                                              �?              @                               @              �?                                      �?      �?                      �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���}hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKyhnh4h7K ��h9��R�(KKy��hu�Bx         :                   �3@�^e���?�	           ��@                           �?��K��?t           @�@                           @�A!ˏ �?�           �@                          �1@z�oƲ��?&           �|@                           @N�i�7��?�            `j@                            �?�|u��2�?R            @a@������������������������       ��K!�H��?5            �T@������������������������       ��e�� �?            �K@	       
                    @3�X=��?3            @R@������������������������       ��)�c{��?             C@������������������������       ���@z��?            �A@                           @T� Pō�?�            @o@                           @���}�?~            @h@������������������������       �ʊ�-�?P             _@������������������������       �>����\�?.            �Q@                           @�r
^N��?#             L@������������������������       ��e�ݥ��?            �B@������������������������       �~�Q���?             3@                            @���3��?�             j@                           �?����-m�?|            �g@                           @G���H�?5             U@������������������������       ��q�q�?             (@������������������������       �������?-             R@                          �2@>�T ��?G            �Z@������������������������       ���.��?3             S@������������������������       �,�Œ_,�?             >@                           @~X�<��?             2@������������������������       �      �?              @������������������������       ��������?             $@       +                   �0@�������?�           ��@       $                     �?�Q�}e�?A             Z@        #                    @8�Z$���?"             J@!       "                    �?d��E���?             A@������������������������       �����W�?	             *@������������������������       �h5����?             5@������������������������       �x�5?,R�?
             2@%       (                     @\�5��?             J@&       '                    �?AA�?             5@������������������������       �r�q��?             (@������������������������       ��<ݚ�?             "@)       *                    @]"?ӧ
�?             ?@������������������������       �"P7��?             3@������������������������       ��8��8��?             (@,       3                     @۪��	�?�           X�@-       0                    @���?�            P{@.       /                     �?��<ߋ��?s            �h@������������������������       �/��6i��?`            �c@������������������������       �Cȍ�n�?            �D@1       2                    @Pg��(��?�            �m@������������������������       ���k�?a            `d@������������������������       �d��D��?+            �R@4       7                    @2��8X�?�            �j@5       6                   �1@DOs9�D�?e            �d@������������������������       �o�����?0            @S@������������������������       �rr�ϛ�?5            @V@8       9                   �2@�8��8N�?             H@������������������������       ���I!��?            �B@������������������������       ��T�x?r�?             &@;       Z                   �8@I��q�?"           r�@<       K                    �?�*��e�?�           T�@=       D                     @)À����?�           �@>       A                   �6@�/h\B�?C           �@?       @                    �?q�O��?�            @u@������������������������       ��z�<p�?B             Z@������������������������       �+&a�1��?�            �m@B       C                    @/�����?n             e@������������������������       �Lz�Dc�?F            �[@������������������������       �����?(             M@E       H                    �?�l,����?            �h@F       G                   �6@,78�/��?+            �Q@������������������������       ���j�y��?             G@������������������������       ��q�q�?             8@I       J                    @��1k��?T             `@������������������������       �;�NW��?F            �Z@������������������������       ���,d!�?             7@L       S                    @�9,\���?           ��@M       P                     @ �B�>��?m           ��@N       O                    �?K>�:F�?�            �v@������������������������       ���ո��?7            �U@������������������������       �"��HQ4�?�            pq@Q       R                    @���QI��?             i@������������������������       ���^B{	�?7            �V@������������������������       ��U}��`�?H            �[@T       W                    @�3����?�            �q@U       V                   �6@�|�f�?�            �o@������������������������       ����D�R�?k            �d@������������������������       ��*��c�?6            @V@X       Y                   �6@�>�>�?             >@������������������������       �ffffff�?             4@������������������������       ��(\����?             $@[       j                     �?�5����?A            �@\       c                    @���c�?8           �@]       `                    �?��\�q�?�            @w@^       _                    �?j��pX��?0            @W@������������������������       ��z�����?(            �R@������������������������       �����Gc�?             3@a       b                    �?�c�г�?�            pq@������������������������       ����p9W�?/             S@������������������������       ���nd��?�            `i@d       g                    �?p��Ϭ��?W            �a@e       f                    @     ��?&             P@������������������������       �4%���?             1@������������������������       �`!�2���?            �G@h       i                    @6��Z�?1            �S@������������������������       �
^N��)�?             <@������������������������       �Hk�����?             �I@k       r                   �:@��V<f��?	           z@l       o                    �?A����?_            `b@m       n                    @��+��?3             U@������������������������       ��c���+�?!             J@������������������������       �     ��?             @@p       q                    @ۺ/�3�?,            �O@������������������������       ��������?"             H@������������������������       ��|�j��?
             .@s       v                    @��l���?�            �p@t       u                    @�g�>Æ�?�            �j@������������������������       ��pA���?{            �g@������������������������       �+7����?             7@w       x                    �?ÇՊ~��?             �L@������������������������       �k��\��?	             1@������������������������       ��G�z��?             D@�t�bh�h4h7K ��h9��R�(KKyKK��h��B�G       }@     �R@      u@     �B@     @U@      @@     @R@     ��@     ��@     �N@     �T@     �c@     ��@     �|@      $@     @Q@     �F@     �_@     @P@     �f@       @      \@      @      @              "@     �u@     �q@      ,@      5@     �F@     �j@     �\@              (@       @      ?@      $@     @T@      @      A@       @                      �?     `i@     �b@      $@      @      3@      Y@     �E@              @              @      @     �O@      @      >@       @                      �?     @_@     �V@       @      @      ,@     �R@      <@              @              @      @      >@       @      &@                              �?     @R@     �I@      @      @      @      <@      @                                              1@              "@                                     �D@     �C@      @      @      �?      5@      @                                              "@               @                                     �@@      <@              @      �?      @       @                                               @              @                                       @      &@      @                      0@       @                                              *@       @       @                              �?      @@      (@                       @      @       @                                               @       @       @                              �?      ,@       @                               @      �?                                              @                                                      2@      @                       @      @      �?                                             �@@       @      3@       @                              J@      D@      @      @      &@     �G@      6@              @              @      @      4@       @      1@       @                              F@      >@      @       @      @     �A@      5@               @              @      @      &@       @      *@                                      9@      3@              �?       @      <@      .@               @               @      @      "@              @       @                              3@      &@      @      �?      @      @      @                              @              *@               @                                       @      $@       @      �?      @      (@      �?              �?              �?              &@              �?                                      @      @       @      �?      @      @      �?              �?              �?               @              �?                                      @      @                      �?      @                                                      2@              @                                     �S@     �M@       @      �?      @      9@      .@              �?                              .@              @                                      S@     �K@       @              @      5@      *@                                              @               @                                      C@      >@                       @      @      @                                                              �?                                       @                                      �?       @                                              @              �?                                      >@      >@                       @      @      �?                                              &@               @                                      C@      9@       @               @      0@      $@                                              @              �?                                      =@      5@      �?               @      ,@      @                                               @              �?                                      "@      @      �?                       @      @                                              @                                                       @      @              �?      �?      @       @              �?                                                                                      �?       @              �?      �?      @                                                      @                                                      �?       @                              �?       @              �?                             @Y@      @     �S@      @      @               @      b@      a@      @      ,@      :@     @\@     �Q@               @       @      8@      @      8@              @                                      C@      1@                              ,@      @                                              .@              �?                                      &@      *@                              $@       @                                              @              �?                                      @      (@                               @                                                      @              �?                                      �?      @                               @                                                      �?                                                      @      "@                              @                                                       @                                                      @      �?                               @       @                                              "@              @                                      ;@      @                              @      @                                              @                                                      ,@                                       @      �?                                               @                                                      $@                                                                                               @                                                      @                                       @      �?                                              @              @                                      *@      @                               @      @                                              @              @                                       @      @                               @      @                                                                                                      &@      �?                                                                                     @S@      @     �R@      @      @               @     �Z@     �]@      @      ,@      :@     �X@      P@               @       @      8@      @     �L@       @     �C@                              @      V@     �V@      @      @      4@      N@      C@              @      @      ,@      @      A@              <@                              �?      <@      ?@       @      @      ,@      =@      0@               @      �?      @      @      @@              0@                                      1@      <@       @      @      $@      6@      .@               @      �?      @      @       @              (@                              �?      &@      @                      @      @      �?                                              7@       @      &@                              @      N@      N@      �?       @      @      ?@      6@               @      @       @              ,@      �?       @                              @      J@     �E@      �?       @      @      4@      .@                              �?              "@      �?      @                               @       @      1@                      @      &@      @               @      @      @              4@       @     �A@      @      @               @      2@      <@      �?      "@      @     �C@      :@              @       @      $@       @      1@       @      6@      @      @                      $@      8@      �?      "@      @      @@      7@               @       @      @      �?      &@              $@              @                      "@      &@              �?      @      "@      ,@               @      �?      �?              @       @      (@      @       @                      �?      *@      �?       @              7@      "@                      �?      @      �?      @              *@                               @       @      @                       @      @      @               @              @      �?      �?              &@                              �?       @      @                      �?      @                      �?              @      �?       @               @                              �?              �?                      �?              @              �?                             �q@     �P@      l@      ?@     �S@      @@      P@     `k@     0s@     �G@     �N@     �[@     �v@     �u@      $@     �L@     �B@      X@     �K@     �h@      7@     `a@      (@      ?@      *@      =@      f@     �n@      2@     �B@     �J@      n@      m@      @      5@      &@      K@      1@     �U@      @     �I@      @      *@      $@      $@      X@     �b@      @      0@      3@     @^@      V@      �?      @      @      0@      @     �P@      @      B@               @              "@     @R@     @^@       @      ,@      *@     @X@     �I@              @      �?      @       @      E@      @      6@               @              @     �D@     �W@      �?      @      @     @S@      7@              �?      �?      @              .@              *@              @              �?      @      *@              @       @      A@       @              �?              �?              ;@      @      "@              @              @      A@     �T@      �?      @      @     �E@      .@                      �?      @              8@       @      ,@                               @      @@      :@      �?      @      @      4@      <@               @               @       @      .@       @      @                              �?      :@      5@      �?      @      @      *@      (@              �?               @       @      "@              @                              �?      @      @              @       @      @      0@              �?                              5@      �?      .@      @      @      $@      �?      7@      =@      @       @      @      8@     �B@      �?              @      $@      @      .@      �?      �?              @       @              @      ,@                               @      0@      �?                      �?      �?      @                              @       @              @      $@                              @      &@                              �?      �?       @      �?      �?              �?                              @                              @      @      �?                                      @              ,@      @      �?       @      �?      1@      .@      @       @      @      0@      5@                      @      "@      @      @              &@      @      �?       @      �?      0@      .@               @      @      (@      *@                      @      @      @                      @                                      �?              @                      @       @                              @             �[@      0@      V@       @      2@      @      3@      T@     @X@      *@      5@      A@      ^@      b@      @      2@      @      C@      &@     @Q@      &@     �P@       @      $@      @      $@      E@     �K@      *@      3@      :@     @S@     �[@              @      @      :@      @     �H@      @     �E@      @      @               @      C@      D@      @      0@      &@      K@      Q@              @      �?      $@      @      &@       @      1@      �?      �?              @      �?      @              @       @      3@      *@                      �?      �?       @      C@       @      :@      @      @              @     �B@     �@@      @      &@      "@     �A@     �K@              @              "@      �?      4@      @      7@       @      @      @       @      @      .@      @      @      .@      7@     �E@              @      @      0@       @      @      @      @              @       @              @      "@      @       @      @      "@      *@              @      @      .@      �?      ,@      @      0@       @       @      �?       @      �?      @      @      �?      &@      ,@      >@                      �?      �?      �?     �D@      @      6@               @              "@      C@      E@               @       @     �E@     �@@      @      &@              (@      @     �D@      @      ,@              @               @     �A@      D@               @      @     �@@      @@       @      &@              (@      @      ;@      �?       @              @              @      ?@      1@               @      @      3@      6@              $@              @      @      ,@      @      @              @              �?      @      7@                      �?      ,@      $@       @      �?              @                               @              �?              �?      @       @                      �?      $@      �?      @                                                       @              �?                       @      �?                      �?      @                                                                                                      �?      �?      �?                              @      �?      @                                     �U@      F@     @U@      3@      H@      3@     �A@     �E@      N@      =@      8@      M@      ^@      ]@      @      B@      :@      E@      C@     �H@      2@      I@      @      0@      @      9@      =@      ?@      .@      0@      ;@     @P@     @T@              8@      0@      8@      .@      ?@      .@      A@      @      *@      @      6@      (@      5@      "@      &@      7@     �B@      P@              5@      (@      5@      *@      ,@      @      @       @                      @       @      @      �?       @      @      &@      9@                      @      @              ,@      @       @       @                      @              @      �?       @      @      &@      .@                      @      @                              @                              �?       @      �?                                      $@                                              1@      (@      ;@      @      *@      @      .@      $@      ,@       @      "@      4@      :@     �C@              5@       @      0@      *@      @      @      @              @       @              @       @       @      �?      @       @      $@              @      �?      �?      @      $@       @      7@      @      @      @      .@      @      @      @       @      .@      2@      =@              0@      @      .@       @      2@      @      0@      �?      @              @      1@      $@      @      @      @      <@      1@              @      @      @       @      0@      �?      @      �?                      @      @      @              @      @      (@      @                                      �?      @      �?                                      �?       @      @               @       @                                                              &@              @      �?                       @      @      �?              @       @      (@      @                                      �?       @       @      (@              @                      (@      @      @                      0@      $@              @      @      @      �?                      @                                      &@      �?      @                               @                       @      �?               @       @      @              @                      �?      @      �?                      0@       @              @       @       @      �?     �B@      :@     �A@      (@      @@      (@      $@      ,@      =@      ,@       @      ?@     �K@     �A@      @      (@      $@      2@      7@       @       @      ,@       @      @      @      @      (@      &@       @       @      $@      >@      &@      �?      @       @       @      $@      @      @      &@       @                       @      @       @               @      �?      5@      @              @      �?      �?      @      @      �?      &@                                      �?      @               @      �?      *@      @               @      �?      �?       @      �?      @               @                       @      @      �?                               @      �?              �?                      @      �?      �?      @              @      @      @      @      @       @              "@      "@      @      �?      @      �?      �?      @      �?      �?       @               @      @       @      @      @       @              "@      @       @      �?      @              �?      @                      �?              @               @      �?                                       @      @                      �?                      =@      2@      5@      $@      :@      "@      @       @      2@      (@      @      5@      9@      8@      @      @       @      0@      *@      ;@      @      &@      @      :@      @      @       @      0@      (@      @      0@      3@      6@      @      @       @      "@      *@      5@      @      $@      @      7@      @      @       @      0@      (@      @      0@      2@      .@      @      @       @      "@      *@      @      �?      �?       @      @       @                                                      �?      @                                               @      *@      $@      @              @      �?               @                      @      @       @               @              @                      "@                                                                              @      �?       @                              �?               @      @      $@      @              @      �?               @                      �?      @                       @              @        �t�bub�2     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��khG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKmhnh4h7K ��h9��R�(KKm��hu�B�         4                   �3@�������?�	           ��@                           �?2�Y���?r           |�@                            @�&���?�           ��@                           @����?D           x�@                           @ �F����?0           `~@                            �?).�	F��?h            @d@������������������������       �����k�?4            @T@������������������������       �8�N���?4            @T@	       
                    �?p1���?�            @t@������������������������       �������?d            �d@������������������������       �#�4�f�?d            �c@                            �?<��b��?            �D@                            �?�ˠT��?             6@������������������������       �g\�5�?             *@������������������������       ���"e���?             "@������������������������       �^Cy�5�?             3@                          �0@�_.��C�?e            �d@                           @r�q��?             8@������������������������       �9��8���?             (@������������������������       �VUUUUU�?             (@                           @5��A��?Y            �a@                           @��-q��?C            @[@������������������������       ������?&            �L@������������������������       �*D>��?             J@                           @d��E���?             A@������������������������       �l �&��?             7@������������������������       ��9����?             &@       )                     @���7��?�           H�@       $                    @�:�I|M�?-           `@       !                    �?�SJ����?�            t@                            @���_E�?7            �V@������������������������       �2���NV�?+            �Q@������������������������       ����c���?             5@"       #                    @C�B��?�            �l@������������������������       �%>]3S�?f            �e@������������������������       ���m�
�?$            �L@%       &                    �?��!l��?l            �f@������������������������       �������?             :@'       (                   �2@U�_w��?]            `c@������������������������       �b'vb'v�?<             Z@������������������������       ����(A�?!            �I@*       -                   �0@��E��&�?�            `n@+       ,                    @HN�zv�?             6@������������������������       �9��8���?             (@������������������������       ���Q��?             $@.       1                    @��F��?�            �k@/       0                    @��q
��?q            `e@������������������������       ������H�?a             b@������������������������       �'��}��?             ;@2       3                    @��^)�?             I@������������������������       ��ۨ:�?            �A@������������������������       ��|�j��?
             .@5       N                    �?��&sE�?           T�@6       C                    �?�ei�iu�?�           Ȑ@7       >                   �6@�*o��c�?�            �u@8       ;                     @?6�^r��?n            `d@9       :                   �4@9�(	r�?V            �_@������������������������       �Ia�T#�?            �D@������������������������       ��W�$���?7            @U@<       =                   �4@&���S)�?            �B@������������������������       ��G�z�?             4@������������������������       ��t����?             1@?       B                   �=@��,j�?o            �f@@       A                   �8@��~0�?d            `d@������������������������       �kN¾�?.             S@������������������������       �fG1�)��?6            �U@������������������������       �kN¾��?             3@D       K                    @_l�ǚ��?�           Ȇ@E       H                    @���;6��?�           �@F       G                   �7@H�O>��?�            px@������������������������       ��,�F.�?{            �h@������������������������       ��0�1���?~             h@I       J                     �?�=Bf:��?�            �s@������������������������       ��eP*L��?2             V@������������������������       ��8|L9��?�            @l@L       M                   �5@�������?             8@������������������������       ��ˠT�?             &@������������������������       ���]�`��?             *@O       ^                    �?�r]5M�?r           ��@P       W                   �8@A�9F;{�?�           ��@Q       T                    �?�=�_a��?�            Px@R       S                     �?���81��?e            @c@������������������������       ���2(&�?             F@������������������������       �T�����?G            �[@U       V                     @�˅�'��?�            `m@������������������������       ��^a�M�?C            �]@������������������������       ����l��?T            @]@X       [                    �?��N���?�             s@Y       Z                   �<@D�]��0�??            @[@������������������������       �     �?$             P@������������������������       �n����?            �F@\       ]                     �?�&H��?            `h@������������������������       �BQ!���?A            �X@������������������������       �9��8���?>             X@_       f                   �9@�#g����?�           �@`       c                    @�vU[N��?P           ؀@a       b                    @婆�9N�?�            �w@������������������������       ��?.4�r�?�            `n@������������������������       ��������?^            �`@d       e                   �5@�mM���?c            `d@������������������������       �OgםS�?&            @P@������������������������       ��YՏ�m�?=            �X@g       j                    @?�!���?h             e@h       i                     �?�������?             H@������������������������       �'��л��?             =@������������������������       �Dy�5��?             3@k       l                    @�7�&��?I             ^@������������������������       ���E$���?#            �J@������������������������       �%�m��L�?&            �P@�t�bh�h4h7K ��h9��R�(KKmKK��h��B�@       |@     @V@      v@      >@      T@      :@     �S@     ��@     H�@      F@     @W@      d@     ��@     0|@      "@      R@      E@      a@      M@     �e@      3@     @Y@      @      $@              (@     �v@      r@       @      2@      @@     �l@     @\@              1@      @      B@      @      T@      @     �C@      �?                      @      k@      d@              @      .@      ]@      B@              �?              $@      �?     �N@      @      6@      �?                      @      g@      _@              @      &@     �U@      7@                              @              G@      @      5@      �?                      @     �e@     @^@               @      $@     �S@      7@                              @              8@              &@                                     �D@     �E@              �?       @      :@       @                                              1@              @                                      .@      8@              �?       @      .@       @                                              @              @                                      :@      3@                      @      &@      @                                              6@      @      $@      �?                      @     �`@     �S@              �?       @      J@      .@                              @              &@       @      �?                                      Q@      F@                       @      A@      @                                              &@      @      "@      �?                      @      P@      A@              �?              2@      &@                              @              .@              �?                                      (@      @              �?      �?       @                                                      @              �?                                       @       @              �?      �?      @                                                      @                                                      @                                      @                                                                      �?                                      @       @              �?      �?                                                              $@                                                      @      �?                              @                                                      3@       @      1@                              @      @@      B@              �?      @      >@      *@              �?              @      �?      @                                                      $@      @                              @                                                      @                                                      @                                      @                                                                                                              @      @                              �?                                                      ,@       @      1@                              @      6@      @@              �?      @      9@      *@              �?              @      �?      ,@       @      (@                              @      4@      2@              �?      @      1@      (@                              @      �?      $@       @                                      @      @      @                       @      &@      "@                              @      �?      @              (@                                      ,@      &@              �?      �?      @      @                                                              @                              �?       @      ,@                      �?       @      �?              �?              �?                               @                                              (@                      �?      @                      �?              �?                              @                              �?       @       @                               @      �?                                             �W@      (@      O@      @      $@              @     �b@     @`@       @      ,@      1@     �\@     @S@              0@      @      :@      @     �Q@      @     �@@      @      @              @      _@     @W@      @       @      *@     �P@      F@              @      @      &@      @      D@      @      6@      @      @              @     �V@     �K@      @      @       @     �G@      9@              @      �?      @      @      ,@       @      $@      @      @                      (@      .@      �?       @       @      .@      @               @               @       @      ,@       @      "@                                      @      .@               @      �?      &@      @               @               @                              �?      @      @                      @              �?              �?      @                                               @      :@      @      (@                              @     �S@      D@      @      @              @@      4@              �?      �?      @      �?      3@      @      "@                               @     @P@      ?@      @      @              0@      2@              �?      �?      �?      �?      @              @                              �?      ,@      "@      �?       @              0@       @                               @              >@      �?      &@              �?              �?     �@@      C@      �?      �?      &@      4@      3@              @      @      @      �?      $@               @                                              @      �?              @      @                                                      4@      �?      "@              �?              �?     �@@      ?@              �?       @      1@      3@              @      @      @      �?      (@              @                              �?      ;@      ,@                       @      (@      ,@              @      @      @      �?       @      �?      @              �?                      @      1@              �?              @      @                              @              8@      @      =@              @              �?      8@     �B@       @      @      @     �G@     �@@              $@              .@              �?       @                       @                      @      @                                       @                                              �?       @                                              @                                              @                                                                               @                      �?      @                                       @                                              7@      @      =@              @              �?      4@      @@       @      @      @     �G@      9@              $@              .@              0@      @      ;@              @              �?      0@      ;@      �?      @       @     �D@      ,@              $@              @              (@      @      :@              @                      $@      4@      �?      @       @      C@      ,@              @              @              @              �?                              �?      @      @                              @                      @                              @               @                                      @      @      �?      �?       @      @      &@                              &@               @              �?                                      @      @                       @      @      $@                               @              @              �?                                              �?      �?      �?               @      �?                              @             0q@     �Q@     `o@      :@     �Q@      :@     �P@     �h@     pt@      B@     �R@      `@     �t@      u@      "@     �K@     �B@     @Y@     �J@      _@      5@     @V@      @      6@      @      1@     @_@     @g@      "@     �B@      G@     �d@     �a@      �?      *@      ,@     �@@      7@     �F@      &@      9@       @      @       @      @     �A@     @V@              "@      @      M@      D@      �?      �?              $@      @      *@      �?      (@                       @      �?      3@     �J@              @      �?     �D@      (@                               @      @      "@      �?      &@                              �?      *@      H@              @      �?      @@      @                                      �?      @                                                      "@      *@                              (@      @                                      �?      @      �?      &@                              �?      @     �A@              @      �?      4@      @                                              @              �?                       @              @      @                              "@      @                               @       @       @                                       @              @      @                              @      @                                               @              �?                                      �?      �?                              @      @                               @       @      @@      $@      *@       @      @              @      0@      B@              @      @      1@      <@      �?      �?               @       @      8@      $@      *@       @      @              @      0@      B@              @      @      &@      :@      �?      �?               @       @      "@      @      @              �?              @      &@      *@              �?       @      @      1@      �?                               @      .@      @      @       @       @                      @      7@               @       @      @      "@              �?               @               @                                                                              @              @       @                                             �S@      $@      P@       @      3@      �?      *@     �V@     @X@      "@      <@     �D@     �Z@     �Y@              (@      ,@      7@      2@     @S@      $@      N@       @      1@      �?      (@     �V@     @W@      @      <@     �D@     �Y@     �Y@              &@      (@      7@      2@     �D@      @     �H@      �?      "@      �?       @      8@     �@@       @      1@      >@      M@     �P@              @      &@      1@      "@      ?@      �?      6@              @      �?      @      4@      7@              &@      *@     �A@      ;@               @               @              $@      @      ;@      �?      @               @      @      $@       @      @      1@      7@      D@              @      &@      .@      "@      B@      @      &@      �?       @              @     �P@      N@      @      &@      &@      F@      B@              @      �?      @      "@      1@              @                              �?      $@      2@                       @      &@      4@              @              �?              3@      @      @      �?       @              @      L@      E@      @      &@      "@     �@@      0@              �?      �?      @      "@       @              @               @              �?              @      @                      @                      �?       @                                                       @              �?               @      @                       @                                                       @              @                                               @                               @                      �?       @                     �b@     �H@     @d@      6@      H@      7@      I@     �R@     �a@      ;@      C@     �T@     �d@     `h@       @      E@      7@      Q@      >@     �N@      =@     @T@      &@      B@      1@      >@      4@     �K@      0@      <@      H@     �S@      X@      @      8@      $@      8@      8@      D@      0@     �H@      @      .@      @      (@      ,@      A@      "@      1@      8@      G@     @R@              @      @      *@      $@      0@      @      4@      �?      @              @      @      *@      @      @      $@      =@      6@              �?       @      @      @                      @      �?      �?              �?       @      @                      @      .@      @                               @      �?      0@      @      ,@              @              @      @      @      @      @      @      ,@      2@              �?       @      @      @      8@      (@      =@      @       @      @      @       @      5@      @      *@      ,@      1@     �I@              @      �?       @      @      1@       @      1@              �?              @      @      *@      @      "@      @      @      9@              @      �?      @      @      @      $@      (@      @      @      @      @       @       @       @      @      "@      *@      :@                               @      @      5@      *@      @@      @      5@      &@      2@      @      5@      @      &@      8@     �@@      7@      @      4@      @      &@      ,@      $@       @      $@              (@      �?      @      @      @       @      @      @      3@      "@               @       @      @      @      $@      @      @              @      �?              @      @       @      �?      @      0@      @              �?                      @              @      @               @              @               @               @       @      @      @              �?       @      @      �?      &@      @      6@      @      "@      $@      (@       @      0@      @       @      2@      ,@      ,@      @      2@      @       @      @      @      �?       @      @      @      @      "@       @      @      @      @      $@      "@      @      �?      .@       @      @      @      @      @      ,@      @      @      @      @              (@       @      @       @      @      "@      @      @      @      �?      @     �V@      4@     @T@      &@      (@      @      4@      K@     �U@      &@      $@      A@      V@     �X@      @      2@      *@      F@      @     @S@      2@     �L@      "@      @              0@      H@      T@      @      $@      3@     @R@     �Q@      @      &@      @      :@      @      L@      (@     �B@      @       @              &@      B@     �Q@       @      $@      ,@      L@     �D@      �?      @       @      (@      �?      A@      @      @@      @       @              "@      6@      >@       @      @      &@      C@      A@              @               @      �?      6@      @      @      @                       @      ,@      D@              @      @      2@      @      �?      @       @      @              5@      @      4@      @      @              @      (@      $@       @              @      1@      =@       @      @      @      ,@      @      *@              @              @              @      "@      @                       @      @      $@              @               @      @       @      @      0@      @      �?               @      @      @       @              @      &@      3@       @              @      (@              *@       @      8@       @      @      @      @      @      @      @              .@      .@      =@      �?      @      @      2@       @       @              @                       @      �?      �?       @      �?               @       @      &@      �?      �?      @      $@      �?                      @                       @                              �?              �?       @       @                      @      "@      �?       @                                              �?      �?       @                      �?              "@      �?      �?              �?              &@       @      1@       @      @      @      @      @      @      @              *@      *@      2@              @       @       @      �?      @       @      &@       @      @      @              �?      �?      @              @      @      @              �?       @      @               @              @              �?              @      @      @                       @      $@      *@              @              @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ/�J\hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         8                    �?>�季��?�	           ��@                           �?��G?*�?           ��@                            �?���T��?%           �|@                          �6@�qUp�f�?X            �`@                           �?NI8d�?5            �R@                           �?     0�?             @@������������������������       �V�Lt�<�?             3@������������������������       ��	j*D�?             *@	       
                    �?�������?             E@������������������������       �s
^N���?
             ,@������������������������       �����S�?             <@                          �8@���}"c�?#            �M@������������������������       �r�q��?             (@                           �?�K2���?            �G@������������������������       �9��8���?             2@������������������������       ���𡌢�?             =@                           �?=��o���?�            �t@                            �?���ml�?P            �`@                           �?�������?"             N@������������������������       ��q�q�?             8@������������������������       �_B{	�%�?             B@                           �?�&�?.            @R@������������������������       �8�V�Ɓ�?            �B@������������������������       ��n���?             B@                            �?�"�ᛊ�?}            �h@                           6@IPolg��?!            �H@������������������������       �n۶m۶�?             <@������������������������       ����H��?             5@                          �3@�U~����?\            `b@������������������������       ���^)�?             I@������������������������       �=u�P��??            @X@        +                   �2@��~�(�?�           l�@!       (                    @�~\�L7�?�            @m@"       %                    �?��S���?�            �i@#       $                   �1@�矆�1�?4            �T@������������������������       �ԍx�V�?             C@������������������������       �Ra���i�?             F@&       '                    �?�e���n�?P            �^@������������������������       ��^B{	��?             B@������������������������       ��i-x|e�?7            �U@)       *                    �?t�@�t�?             >@������������������������       �Iє�?
             1@������������������������       �������?             *@,       3                   �@@��<YBG�?G           ��@-       0                    �?����6�?4           ��@.       /                    @����P�?�            ps@������������������������       ��Ƈ�4y�?y             h@������������������������       ��)_�5m�?M            �]@1       2                    �?��׻gf�?n           ؂@������������������������       ��ѳ�w�?            �I@������������������������       ���4�|p�?T           @�@4       5                   @A@�+O�?             ?@������������������������       ��������?             $@6       7                     @Cu��?             5@������������������������       ��T�6|��?             *@������������������������       �      �?              @9       X                   �2@ŜA4k��?�           ��@:       I                     �?qOƈ�V�?�           @�@;       B                    @W!����?�            @l@<       ?                    @wG���?\            �b@=       >                    @�b�b�?#             O@������������������������       �z�i���?            �D@������������������������       ��%7)��?
             5@@       A                    �?80�B��?9            @V@������������������������       �_L
�8Y�?!            �J@������������������������       �{	�%���?             B@C       F                    @�V�u)9�?-            �R@D       E                   �0@��Kh/�?             B@������������������������       �        	             ,@������������������������       �*L�9��?             6@G       H                    @�(�Tw��?            �C@������������������������       �      �?              @������������������������       �/�E���?             ?@J       Q                    �?ӈ�)�?9           `~@K       N                     @ǫ��u�?�            p@L       M                    @\ʉ����?�            �h@������������������������       ��U]E��?H            �]@������������������������       �
ףp=��?;             T@O       P                    �?a���{�?+             M@������������������������       �������?             1@������������������������       �1OxJ'�?            �D@R       U                     �?8-����?�            �l@S       T                   �1@fffff&�?3             T@������������������������       �0�S�v�?             �I@������������������������       ���-�?             =@V       W                    @�l���?X            �b@������������������������       �A�>�)
�?"             G@������������������������       ��]����?6            �Y@Y       h                   �:@�W�T8��?�           `�@Z       a                    �?���|,�?K           ��@[       ^                   �8@�~R��w�?�           `�@\       ]                    @=¢�9�?a           ��@������������������������       ��۷c��?[           p�@������������������������       ���(\���?             $@_       `                    @	�kv�"�?8             U@������������������������       ���T���?/            �Q@������������������������       �^N��)x�?	             ,@b       e                    �?��ˇ��?�           ��@c       d                   �8@���}��?�            @j@������������������������       ��l����?u            @g@������������������������       ��������?             8@f       g                    @xsK��?.            ~@������������������������       �ɕ����?1            �R@������������������������       �uG��?�            �y@i       p                    �?��@M^�?�             o@j       m                   �=@z�:���?<            @U@k       l                     �?ʃg\��?$             J@������������������������       ��
t�F��?	             1@������������������������       ����v��?            �A@n       o                    @��u��?            �@@������������������������       �p=
ףp�?             $@������������������������       �l �&��?             7@q       t                    @���w�?a            `d@r       s                    @��Yi��?A             [@������������������������       ����eP*�?             F@������������������������       �     ��?(             P@u       v                     �?j�V���?             �K@������������������������       �l+�2���?             ?@������������������������       �9��8���?             8@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       �}@     �V@     u@      <@     �R@      A@      R@     �@     �@      R@     �S@     �g@     P�@     Pz@      0@     @Q@      A@     �`@     �K@      j@      F@      d@      (@     �G@      ;@      @@     �_@     @f@     �A@     �F@      \@     �l@     �i@      &@      E@      8@     �N@      C@      W@      .@      A@      �?      ,@      @      "@     �B@     �K@      @      @      4@      M@     �J@      @      *@       @      6@       @      <@              (@              @               @      $@      1@      @              $@      *@      *@      @               @      *@              3@              @              �?              �?      "@      ,@                      @      "@      @                      �?      �?              @              @                              �?      @      @                      �?      @      @                      �?                      @              @                                      @      @                               @      @                                               @              �?                              �?       @      @                      �?       @                              �?                      (@              @              �?                      @       @                      @      @      @                              �?               @               @              �?                      @                               @      @                                                      $@              �?                                               @                      @       @      @                              �?              "@              @              @              �?      �?      @      @              @      @      @      @              �?      (@              �?               @                              �?      �?              @                               @                      �?                       @              @              @                              @      �?              @      @      @      @                      (@              @                                                              @                              @      @                              @               @              @              @                                      �?              @      �?       @      @                      "@              P@      .@      6@      �?      $@      @      @      ;@      C@      �?      @      $@     �F@      D@              *@      @      "@       @      4@      @      "@              �?               @      .@      5@              @      @      2@      3@               @      @      �?      @      @      @      �?                               @      @      (@               @       @      "@      &@              @                      @      �?      @      �?                                       @      @                              @      @                                      �?      @                                               @       @      @               @       @      @      @              @                       @      ,@               @              �?                      &@      "@               @      @      "@       @              @      @      �?      �?      &@              @                                      @      @                      �?      @       @               @              �?              @              @              �?                      @      @               @       @      @      @              �?      @              �?      F@      (@      *@      �?      "@      @      @      (@      1@      �?       @      @      ;@      5@              @      @       @      @      2@       @      @               @              @      @      �?                              @      @                              �?      �?      ,@              @                                      @      �?                              @                                              �?      @       @       @               @              @                                              �?      @                              �?              :@      $@       @      �?      @      @              @      0@      �?       @      @      7@      1@              @      @      @      @       @       @       @              �?                       @      $@              �?               @      $@                              @              2@       @      @      �?      @      @              @      @      �?      �?      @      .@      @              @      @      �?      @     @]@      =@     �_@      &@     �@@      4@      7@     �V@     �^@      =@     �C@      W@     �e@      c@      @      =@      0@     �C@      >@      ?@       @      2@              �?               @     �I@      F@      @      @       @      E@      6@                      �?      @      �?      5@       @      .@              �?               @     �G@     �E@       @       @      @      D@      2@                      �?      @               @       @      �?                              �?      8@      7@                       @      .@      @                              �?              @                                                      .@      *@                              @      �?                                              @       @      �?                              �?      "@      $@                       @      &@      @                              �?              *@              ,@              �?              �?      7@      4@       @       @      @      9@      *@                      �?      @              @              @                                      @      &@                      �?      @      @                                              "@              @              �?              �?      2@      "@       @       @      @      4@      $@                      �?      @              $@              @                                      @      �?      �?       @       @       @      @                                      �?      @               @                                              �?      �?       @       @       @                                                      @              �?                                      @                                              @                                      �?     �U@      ;@     @[@      &@      @@      4@      5@     �C@     �S@      :@     �A@      U@     @`@     ``@      @      =@      .@     �A@      =@     @U@      ;@     �Z@      &@      ?@      4@      5@     �C@     �S@      :@     �@@     �Q@     @`@     ``@              =@      ,@     �@@      <@      C@      @      <@      �?      $@       @      @      4@      9@      @      @      5@     �Q@      F@              @       @      &@      @      :@      @      9@      �?      "@       @      @      &@      1@      @      �?      ,@     �C@      5@              �?      @      "@       @      (@              @              �?              �?      "@       @      @      @      @      @@      7@              @      @       @      @     �G@      5@     �S@      $@      5@      2@      1@      3@      K@      4@      <@     �H@     �M@     �U@              9@      @      6@      5@              @       @               @                      �?      @       @      @      @       @      4@               @                             �G@      2@     @S@      $@      3@      2@      1@      2@      I@      (@      9@     �F@     �L@     �P@              7@      @      6@      5@      �?               @              �?                                               @      ,@                      @              �?       @      �?      �?              �?                                                              �?      @                       @                       @                              �?              �?                                              �?      &@                      @              �?              �?                      �?                                                                      $@                                      �?              �?                                      �?                                              �?      �?                      @                                     �p@      G@      f@      0@      <@      @      D@     �{@     �z@     �B@      A@      S@     @t@     �j@      @      ;@      $@     �R@      1@      S@      @     �C@              �?              @     �n@     �d@      @      "@      *@     @W@     �B@              @              "@      @      ?@      @      @                               @     �N@      S@      �?       @      @      9@      $@                              @      �?      7@      @      @                                      H@      F@               @       @      1@      @                              �?      �?      *@              @                                      (@      0@               @      �?      &@      @                                      �?      "@              @                                      @      $@               @      �?       @      @                                      �?      @                                                       @      @                              @                                                      $@      @                                              B@      <@                      �?      @      @                              �?              @                                                      8@      2@                      �?      @      @                                              @      @                                              (@      $@                              @      �?                              �?               @                                               @      *@      @@      �?              @       @      @                              @                                                               @      @      8@      �?               @      �?      �?                               @                                                                              ,@                                                                                                                                       @      @      $@      �?               @      �?      �?                               @               @                                                      $@       @                       @      @       @                               @               @                                                              @                      �?       @                                                      @                                                      $@      @                      �?      @       @                               @             �F@       @      B@              �?              @      g@     @V@      @      @      @      Q@      ;@              @              @       @      =@      �?      ,@                                     �\@     �G@      @               @     �A@      (@                                              6@      �?      @                                     @Y@     �A@                       @      9@      "@                                              $@      �?                                              O@      :@                       @      0@       @                                              (@              @                                     �C@      "@                              "@      @                                              @              $@                                      *@      (@      @                      $@      @                                              �?              @                                       @      @                              �?      �?                                              @              @                                      &@      @      @                      "@       @                                              0@      �?      6@              �?              @     �Q@      E@      �?      @      @     �@@      .@              @              @       @      @      �?      @                               @      1@      1@               @       @      0@      @              @               @              @      �?      @                                       @      .@               @       @      (@      �?                              �?               @                                               @      "@       @                              @      @              @              �?              $@              1@              �?              @      K@      9@      �?      @      @      1@       @              �?               @       @      @               @              �?              �?      $@      @      �?      @      @      &@      �?                                              @              .@                               @      F@      2@                              @      @              �?               @       @     �g@     �D@      a@      0@      ;@      @     �@@      i@     `p@      @@      9@     �O@     �l@     @f@      @      7@      $@     @P@      ,@     �d@      7@     �Z@      (@      4@      �?      9@      h@     �o@      4@      5@     �G@      i@     @a@      @      3@      @      H@      (@     @S@       @     �H@      �?      @      �?      @      Z@     �b@      .@      $@      (@      V@     @Q@              @      @      0@      @     �N@      @     �D@      �?      @      �?      @     @X@     �`@      .@      @      $@     @S@     �L@               @      @      .@       @     �N@      @      D@      �?      @      �?      @     @X@     �`@      $@      @      $@      S@     �L@               @       @      .@       @                      �?                                              �?      @                      �?                               @                      0@      @       @              �?              �?      @      *@              @       @      &@      (@               @              �?       @      .@      @       @              �?              �?      @      &@               @       @      &@      "@              �?              �?       @      �?                                                      @       @              @                      @              �?                             @V@      .@     �L@      &@      .@              4@      V@      Z@      @      &@     �A@      \@     @Q@      @      .@      @      @@       @     �@@      �?      1@      @       @              @     �@@      B@      @      �?      @      2@      @@              $@      �?      @      �?      =@      �?      .@      @       @              @      =@      B@              �?      @      0@      >@              @      �?      @      �?      @               @                              @      @              @                       @       @              @                              L@      ,@      D@       @      *@              ,@     �K@      Q@      �?      $@      =@     �W@     �B@      @      @       @      :@      @      (@      @      $@       @      @              @      ,@      $@                              (@       @                              �?              F@      &@      >@      @       @              &@     �D@      M@      �?      $@      =@     �T@     �A@      @      @       @      9@      @      9@      2@      ?@      @      @      @       @       @      $@      (@      @      0@      ?@      D@       @      @      @      1@       @       @      @      @       @      @                      @      @      �?       @       @      3@      0@                              @              @      @      @       @      @                      @      @               @      �?      "@      @                              @              @      @                                               @                                      �?      @                              @                      @      @       @      @                      @      @               @      �?       @                                      @              @               @              �?                      �?      �?      �?              �?      $@      *@                                              �?               @                                                                              @                                                       @                              �?                      �?      �?      �?              �?      @      *@                                              1@      &@      :@       @       @      @       @      �?      @      &@       @      ,@      (@      8@       @      @      @      $@       @      &@      $@      ,@       @       @      @              �?      @      &@       @      ,@       @      .@       @               @       @      �?      @              @      �?       @      @                               @              @      @      @      �?              �?              �?       @      $@       @      �?               @              �?      @      @       @      "@      @       @      �?              �?       @              @      �?      (@                               @              �?                              @      "@              @      �?       @      �?      @              "@                              @              �?                              @      @              @      �?      �?      �?      @      �?      @                              @                                              �?      @                              @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKqhnh4h7K ��h9��R�(KKq��hu�B�         2                   �5@T|R�v��?�	           ��@                          �0@����?u           8�@       
                     �?���?�             i@       	                    @���H��?M            @\@                           �?1�n����?=            �V@������������������������       �����2�?             .@                           �?80\�Uo�?2             S@������������������������       ���{u��?            �C@������������������������       ��-����?            �B@������������������������       �$��Z=;�?             6@                           @�V���?;             V@                            @�%����?            �D@������������������������       ���[r��?             5@������������������������       �      �?             4@                           @@��"��?#            �G@                           �?� =[y�?             1@������������������������       ���E���?             "@������������������������       �      �?              @                           @�&���?             >@������������������������       ��X�C�?             ,@������������������������       �      �?             0@       #                    �?��+�~��?�           L�@                          �1@�p�dg�?�           ��@                           �?�o
��]�?X            �`@                           @�����d�?             K@������������������������       ��B'U�?            �@@������������������������       ��u]�u]�?             5@                           @������?9             T@������������������������       �������?-            �P@������������������������       �����>4�?             ,@       "                    @��"=s�?u           ��@        !                     @F�y^n�?n           P�@������������������������       �F����=�?�            �t@������������������������       ��L&�V�?�            �o@������������������������       �r�q��?             (@$       +                    @�>YѠU�?            ܓ@%       (                     @Hv���?[           @�@&       '                    �?i�Y�B��?�           �@������������������������       �S�0b�M�?�             q@������������������������       �!}��wG�?            �|@)       *                    �?c{�����?�            �l@������������������������       �i�CדS�?D             [@������������������������       ����}��?E            �^@,       /                    �?�������?�            �r@-       .                    �?����1�?J            �\@������������������������       �JC�ɯ�?)            �L@������������������������       �V+�io�?!            �L@0       1                     �?�T�\P�?{            �g@������������������������       ��d�����?&            @P@������������������������       ��+\&p�?U             _@3       R                    �?c>�WU�??           ��@4       C                    �?7�A���?�            �@5       <                     �?��"B���?�             m@6       9                   �:@�>���}�?\            �a@7       8                    @      �?@             X@������������������������       ���>z��?/             Q@������������������������       �?4և���?             <@:       ;                    �?�&EՁ��?            �F@������������������������       ��?�P�a�?             >@������������������������       �؂-؂-�?
             .@=       @                   �7@B���j�?7             W@>       ?                     @'��л��?             =@������������������������       �t�@�t�?             .@������������������������       ��X�C�?             ,@A       B                   �9@��y�
�?(            �O@������������������������       �      �?             @@������������������������       ��+\&p�?             ?@D       K                     �?_@z��?.           p}@E       H                    @     B�?W             `@F       G                    @gL��J�?'             M@������������������������       �J���#��?             6@������������������������       �����K�?             B@I       J                   �;@�r���2�?0            �Q@������������������������       �pΈ����?"             I@������������������������       �\���(\�?             4@L       O                     �?$ ,S!�?�            pu@M       N                    @?~�.�_�?R            ``@������������������������       ��F�!�5�?H            @]@������������������������       ��>4և��?
             ,@P       Q                    @F��')�?�            �j@������������������������       ��P�m
�?a            `c@������������������������       ��4S�1��?$            �L@S       b                    @mm�H�~�?~           h�@T       [                    �?,�`�p�?�           Ȇ@U       X                   �<@�bH�"��?           �x@V       W                     �?�G!�2&�?�            �r@������������������������       ��r@+�?d             c@������������������������       ������?_            �b@Y       Z                     @h����z�?>            �V@������������������������       �Z�9�(l�?%             K@������������������������       �?,R�n�?             B@\       _                   �:@���g��?�             u@]       ^                   �7@S�Te�Z�?�            �j@������������������������       �     ��?B             \@������������������������       �\J����?C            @Y@`       a                     @BՍ���?K            �^@������������������������       �>�X�q��?9             W@������������������������       ���QN�?             ?@c       j                    @��3�?�?�            @q@d       g                    �?�h0M��?l            `f@e       f                   @A@Ǎ�[�/�?T            ``@������������������������       ��I/�u�?N            �]@������������������������       �*D>��?             *@h       i                    @�8��8��?             H@������������������������       �:2��h�?             =@������������������������       ��d�����?             3@k       n                   �8@�F1-C�?A            @X@l       m                    @ �}��?'            �L@������������������������       �x9/���?             <@������������������������       �K�]l���?             =@o       p                    @�z�G��?             D@������������������������       �+f��ӫ�?             5@������������������������       �ԍx�V�?             3@�t�bh�h4h7K ��h9��R�(KKqKK��h��BC       y@     @S@     @u@      =@      S@      5@     �V@     ��@     ��@     �Q@      X@     @g@     `�@     �{@      (@      R@     �G@     @a@     �P@     �p@      ,@     �c@      *@      *@      �?      A@     �|@     y@      4@     �B@     �X@     �v@     �j@              9@      &@      Q@      1@      @@      �?      @                                     @U@      D@              �?              <@      "@                              �?              4@              @                                      C@     �@@              �?              ,@      @                              �?              4@              @                                      A@      5@              �?              &@                                      �?              @              �?                                      @       @                                                                                      1@               @                                      ?@      *@              �?              &@                                      �?              @                                                      6@      @              �?               @                                                      $@               @                                      "@      @                              "@                                      �?                                                                      @      (@                              @      @                                              (@      �?      �?                                     �G@      @                              ,@      @                                              $@      �?                                              2@      �?                              $@      �?                                              @                                                      (@                                      @                                                      @      �?                                              @      �?                              @      �?                                               @              �?                                      =@      @                              @      @                                               @                                                      @       @                               @      @                                               @                                                      @      �?                                      �?                                                                                                       @      �?                               @      @                                                              �?                                      6@      @                               @      �?                                                              �?                                       @      @                               @                                                                                                              ,@      �?                                      �?                                              m@      *@      c@      *@      *@      �?      A@     @w@     �v@      4@      B@     �X@     �t@     �i@              9@      &@     �P@      1@     �X@      @      L@      @      @              @     �V@      X@      "@      7@     �D@      `@     @X@              0@       @     �B@      $@      4@              @              �?                     �@@      &@      @      @      $@      7@      1@                      �?      @       @      (@              �?                                      3@      @      @              @      @       @                              @              @              �?                                      0@              �?              @      @       @                                              "@                                                      @      @       @                                                              @               @              @              �?                      ,@       @              @      @      4@      .@                      �?      �?       @       @              �?              �?                      @      @              @      @      2@      ,@                      �?      �?      �?                       @                                      @      �?                               @      �?                                      �?     �S@      @      J@      @      @              @      M@     @U@      @      3@      ?@     @Z@      T@              0@      @      @@       @      S@      @      J@      @      @              @      M@     @U@      @      3@      =@     @Z@     �R@              0@      @      @@       @     �K@      �?     �@@      @      �?              @     �C@      J@      @      (@      1@      K@      @@              "@              *@      @      5@      @      3@               @              @      3@     �@@      @      @      (@     �I@      E@              @      @      3@      @       @                              �?              �?                                       @              @                                             �`@      @     @X@      "@       @      �?      ;@     �q@     �p@      &@      *@     �L@     �i@     �Z@              "@      @      >@      @     �X@      @     �U@      @       @      �?      1@      m@     �h@      &@      "@     �E@     `d@     �Q@              @       @      0@      @     @Q@      @      K@      @                      ,@     �h@     `d@      &@      @      =@     �[@      M@              @       @      &@      @      2@               @                               @      U@     �R@      @       @      ,@     �G@      3@                                      @     �I@      @      G@      @                      (@     @\@     @V@       @      @      .@      P@     �C@              @       @      &@              =@      �?      @@      @       @      �?      @      B@     �@@              @      ,@      J@      *@                              @       @      1@              (@                      �?              ;@      ,@               @       @      :@      @                              @              (@      �?      4@      @       @              @      "@      3@               @      (@      :@      "@                               @       @      B@      @      &@       @      @              $@      H@     @Q@              @      ,@      E@      B@              @      �?      ,@       @      0@              @              @              @      ,@      5@              �?       @      &@      =@              �?              @      �?      @              @                                      (@      0@              �?       @      @      $@                                              $@              @              @              @       @      @                              @      3@              �?              @      �?      4@      @      @       @       @              @      A@      H@              @      (@      ?@      @              @      �?      &@      �?      @      @       @       @      �?               @      "@      7@                       @      $@                              �?      @              1@               @              �?              @      9@      9@              @      $@      5@      @              @              @      �?      a@     �O@     �f@      0@     �O@      4@      L@     @Z@     �h@      I@     �M@      V@     `l@     �l@      (@     �G@      B@     �Q@     �H@     �O@      9@      S@      @      .@      @      5@      N@     �\@      "@      7@      ?@      X@     �V@      @      ,@      .@      6@      .@      >@      "@      7@      �?      @              @      1@      M@       @      @      @      =@      :@      @      @       @      @      �?       @      @      3@      �?      @              @      &@     �C@       @      @       @      1@      2@                       @       @      �?      �?              2@      �?      �?              @      &@      :@       @      @      �?      (@      &@                               @      �?                      (@      �?      �?              @       @      4@       @      @      �?      &@      @                               @      �?      �?              @                                      "@      @              �?              �?      @                                              @      @      �?               @               @              *@               @      �?      @      @                       @                      @      @                       @              �?               @               @                      @                       @                      �?              �?                              �?              @                      �?      @      �?                                              6@      @      @                                      @      3@                      @      (@       @      @      @              �?              $@      �?      �?                                      @       @                       @      @      �?      @                                       @              �?                                      @       @                       @      @      �?                                               @      �?                                                                                       @              @                                      (@      @      @                                       @      1@                      @      @      @              @              �?              @      �?                                               @      ,@                      �?       @      @               @              �?              @      @      @                                              @                       @      @      @              @                             �@@      0@     �J@       @      (@      @      ,@     �E@     �L@      @      1@      8@     �P@     @P@       @       @      *@      3@      ,@      $@      @      .@                               @       @      *@      �?      @      @      4@      ;@              @      �?      (@       @      �?      @      @                              �?      �?      @              @       @      @      4@               @              "@                      �?      �?                              �?      �?                      �?              @      @              �?              @              �?       @       @                                              @              @       @       @      0@              �?               @              "@       @      (@                              @      �?       @      �?      �?      �?      *@      @               @      �?      @       @       @       @      (@                              @      �?      @      �?      �?      �?      @      @               @              @              �?                                              �?              @                              "@       @                      �?               @      7@      &@      C@       @      (@      @      @     �D@      F@      @      (@      5@     �G@      C@       @      @      (@      @      (@      &@      @      @      �?       @              �?      4@      7@              @      @      ,@      6@              @      @              @       @      @      @      �?       @              �?      1@      5@              @      @      *@      6@              �?      @              @      @                                                      @       @                              �?                       @       @              �?      (@      @      ?@      �?      $@      @      @      5@      5@      @      @      0@     �@@      0@       @      �?      @      @      @      "@      @      7@      �?      "@      @      @      @      0@      @      @      0@      :@      &@       @      �?      @              @      @      @       @              �?                      ,@      @       @       @              @      @                              @             �R@      C@     �Z@      *@      H@      .@     �A@     �F@     �T@     �D@      B@     �L@     ``@     �a@      @     �@@      5@      H@      A@     �G@     �@@     �S@      $@     �A@      ,@      2@     �B@     �Q@     �B@      7@     �@@     @U@     �[@      @      8@      1@      A@      0@      <@      *@     �C@      @      =@      &@      *@      .@      7@      2@      0@      3@      B@      P@      @      *@      (@      3@      .@      ;@      (@      ;@      @      4@      "@       @      *@      3@      .@      $@      *@      B@      M@      �?      @      @      ,@      &@      .@      @      .@      �?      *@       @      �?      &@      @      @      "@      @      8@      5@      �?      @      �?      @      @      (@      @      (@      @      @      @      �?       @      ,@       @      �?       @      (@     �B@               @      @       @      @      �?      �?      (@       @      "@       @      &@       @      @      @      @      @              @       @      @       @      @      @      �?               @      �?      "@               @              @              @      @               @              @      @      @                      �?      @      �?               @      @       @      �?      @       @                      @       @      @      @      �?      @      3@      4@      D@      @      @      @      @      6@     �G@      3@      @      ,@     �H@     �G@      @      &@      @      .@      �?      0@       @      5@       @      @              @      3@      B@       @      @      @      C@      @@      �?      &@              @              &@      �?      *@      �?                      @       @      ,@      @              @      1@      ;@              @               @              @      @       @      �?      @               @      &@      6@      @      @              5@      @      �?      @              @              @      (@      3@      �?      �?      @              @      &@      &@      @      &@      &@      .@       @              @      $@      �?       @      @      3@      �?      �?      @              �?       @      &@      @      @      @       @       @              @      @              �?      @                                               @      @                      @      @      @                              @      �?      ;@      @      <@      @      *@      �?      1@       @      (@      @      *@      8@      G@      =@      �?      "@      @      ,@      2@      ,@      @      3@      @      "@      �?      (@       @      "@      @      *@      4@      3@      (@      �?      @      @      $@      2@      $@      @      2@      �?       @      �?      &@      �?       @      @      *@      ,@      0@      &@      �?      @      @      @      (@      $@      @      2@               @      �?      &@      �?       @      @      *@      "@      0@      &@      �?      @      @      @      @                              �?                                                              @                                                      @      @              �?       @      @              �?      �?      @                      @      @      �?              @              @      @                      �?                                      �?      @                      @      @      �?                              @      @      @                       @      @              �?                                      �?                              @              �?              *@      �?      "@              @              @      @      @      �?              @      ;@      1@               @      �?      @              @      �?      @              @              �?      @      @                      @      *@      @              �?      �?      @              @               @              �?              �?      @      @                              $@      �?              �?              �?              @      �?      @              @                       @                              @      @      @                      �?       @              @               @                              @                      �?              �?      ,@      $@              �?              �?              @                                                                      �?              �?      @      @              �?              �?                               @                              @                                               @      @                                        �t�bub�     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��=hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         8                   �2@����Ǆ�?�	           ��@                          �0@��ֶ��?�           X�@                           @Je�6H�?�            `i@                           �?	Ǳ�,��?e            `c@                            �?�ݷP�*�?:            �U@                           �?Sl �?&            �K@������������������������       ��^�q��?            �@@������������������������       �_�g����?             6@	       
                     @�H���?             ?@������������������������       ��Q����?             .@������������������������       �      �?	             0@                           @ܳ�.���?+            @Q@                           �?�"w����?             C@������������������������       ��Q����?             $@������������������������       �����X�?             <@                            �?8,�̂�?             ?@������������������������       �kN¾��?             3@������������������������       ��q�q�?             (@                           @��8����?              H@                            �?j�J�Z��?            �@@������������������������       �ףp=
�?             4@������������������������       �؉�؉��?             *@                           @n�����?             .@������������������������       �      �?             @������������������������       �VUUUUU�?             "@       )                    �?`I&�;�?           X�@       "                    �? �!�:�?           �{@                           �?��o$%��?O            �`@                           �?~h����?"             L@������������������������       ��2Tv��?             >@������������������������       �8�Z$��?             :@        !                     @��Դ��?-             S@������������������������       ��,o��?            �D@������������������������       ��!�>���?            �A@#       &                     @
{��%s�?�            �s@$       %                   �1@f�6D`��?�            �o@������������������������       ���3E�T�?I            �]@������������������������       ������H�?N            �`@'       (                   �1@`s���?'            �N@������������������������       �     P�?             @@������������������������       �ܷ��?��?             =@*       1                    @	
�fa��?           �|@+       .                   �1@�<��E�?�            �s@,       -                    @)����?b            `d@������������������������       ���[4�?I            �^@������������������������       �L�J��}�?            �D@/       0                    �?�T�,tM�?R            �b@������������������������       ��ؓo�?#             O@������������������������       �|�nol�?/            �U@2       5                    @���h��?Z            �b@3       4                     @�Q����?             D@������������������������       ��U̠ç�?             5@������������������������       �(������?	             3@6       7                   �1@tN��?F            @[@������������������������       ���7����?            �E@������������������������       �~j{3���?'            �P@9       X                   �7@�z#Z���?           �@:       I                    �?�I#/�S�??           h�@;       B                    �?3��E��?�           ��@<       ?                     �?�Z�p��?�            �m@=       >                    �?��[���?,            �P@������������������������       �     p�?             @@������������������������       ����W��?            �A@@       A                     �?ʾ���t�?z            �e@������������������������       �P�����?4            �Q@������������������������       � *4>HR�?F            �Y@C       F                    �?�h�d.�?	           @z@D       E                    �?��?j�/�?W            @a@������������������������       �0)L�?'            �N@������������������������       �Pj(��?0            @S@G       H                    �?��v/
A�?�            �q@������������������������       ���-��?L            @_@������������������������       ����?�?f            �c@J       Q                     @N�끑��?�           �@K       N                   �6@������?           H�@L       M                    @1�%0�n�?�           �@������������������������       �V�U���?X             b@������������������������       �񎴠��?h           ��@O       P                    @�m�1��?U             a@������������������������       �Fi���?9             W@������������������������       ����eP*�?             F@R       U                    �?,�ͬ4��?{            �g@S       T                   �5@j<ⴇ�?/            @U@������������������������       ��Z��L��?&            �Q@������������������������       �������?	             ,@V       W                    @ �����?L            @Z@������������������������       ��V���?             6@������������������������       ��-��-��?>            �T@Y       h                    �?��_^B^�?�           d�@Z       a                     �?*�8�G�?�             q@[       ^                    �?Z4���?.            �P@\       ]                    �?b���i��?            �@@������������������������       ��θ�?             *@������������������������       ���Q��?             4@_       `                   �9@%����?             A@������������������������       �������?             &@������������������������       ��Ӫ�Ep�?             7@b       e                   �;@���cD�?�            �i@c       d                    @�zS��?U            �`@������������������������       �jM�S�??             Y@������������������������       �d �?�*�?            �A@f       g                    @�[�mT�?2            �Q@������������������������       �r�qG�?"             H@������������������������       ��zv��?             6@i       p                   �>@b�~'W�?*           H�@j       m                   �9@Y��T��?�           (�@k       l                    �?�.}*َ�?�            �t@������������������������       ��N8���?T            �_@������������������������       �+@;����?            @i@n       o                    @�&r$�?�            �w@������������������������       �g8�$N>�?�            Pt@������������������������       �����>4�?#             L@q       t                    @��sS]��?Y            �`@r       s                   �@@2��.��?>            �V@������������������������       �a
��F�?$            �J@������������������������       �cT!)��?             C@u       v                    @=��G��?            �D@������������������������       ���1G���?             *@������������������������       ��$I�$I�?             <@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       �{@     @S@     `w@      @@      M@      =@     �U@     �@     8�@     �R@     @V@      e@     p�@      {@      $@     �K@      G@     �Y@      K@      a@      1@     �T@              @              "@     0r@     �k@      @      "@      ;@     �f@      V@              $@      @      1@       @      =@      @      @                                     �R@     �K@              �?              5@      "@                              @              5@      @      @                                     �P@     �@@              �?              .@       @                              @              &@               @                                      F@      3@              �?              "@                                                       @              �?                                      <@      *@              �?              @                                                      @              �?                                      4@      @              �?               @                                                      @                                                       @      "@                               @                                                      @              �?                                      0@      @                              @                                                                                                              "@      @                              @                                                      @              �?                                      @      @                               @                                                      $@      @      �?                                      7@      ,@                              @       @                              @               @      @      �?                                      @       @                              @      @                                                                                                       @      @                               @                                                       @      @      �?                                      @       @                              @      @                                               @                                                      0@      @                              �?      @                              @               @                                                       @      @                                                                      @                                                                       @                                      �?      @                                               @              @                                      @      6@                              @      �?                                              @              @                                              4@                              @      �?                                                                                                              2@                               @                                                      @              @                                               @                              @      �?                                              @                                                      @       @                              �?                                                      �?                                                      @      �?                                                                                      @                                                      @      �?                              �?                                                      [@      *@     �R@              @              "@      k@      e@      @       @      ;@     @d@     �S@              $@      @      ,@       @      J@      @      >@                              @     �^@     �X@      �?      �?      $@      S@      D@              @              @              8@       @      @                                      8@      5@      �?      �?       @      @@      @              @              @              &@       @       @                                      .@      @      �?               @       @      @              �?              @              "@               @                                      @       @      �?               @      @       @              �?              �?               @       @                                              "@      @                              @      @                               @              *@              @                                      "@      .@              �?      @      8@       @              @                              $@              �?                                      @       @              �?      @      $@                                                      @               @                                      @      @                              ,@       @              @                              <@      �?      9@                              @     �X@     @S@                       @      F@     �@@                               @              5@      �?      @                              @      V@     �P@                       @     �@@      =@                               @              (@                                              @      H@     �@@                      �?      ,@      @                               @              "@      �?      @                                      D@      A@                      �?      3@      8@                                              @              2@                                      &@      $@                              &@      @                                               @              @                                      @       @                              "@       @                                              @              (@                                      @       @                               @       @                                              L@      $@     �F@              @              @     �W@     �Q@      @      @      1@     �U@     �C@              @      @      "@       @     �E@       @      B@              @              @      P@      F@       @      @      "@     @Q@      ,@               @              @      �?      :@      �?      ,@              @              �?      C@      6@              @      "@     �A@      @                                      �?      7@      �?      ,@              @              �?      >@       @              @      @      6@      @                                      �?      @                                                       @      ,@                      @      *@                                                      1@      @      6@                              @      :@      6@       @                      A@      "@               @              @              @       @      .@                                      @      1@      �?                      &@      @                              @              *@      @      @                              @      6@      @      �?                      7@      @               @              �?              *@       @      "@                              �?      >@      :@      @      �?       @      1@      9@              @      @      @      �?      �?       @                                              &@      @       @               @      @      @              @      �?                                                                               @      @       @              �?      @      �?                                              �?       @                                              @      @                      �?              @              @      �?                      (@              "@                              �?      3@      3@      �?      �?      @      &@      4@              �?      @      @      �?       @               @                                      &@       @      �?              @      @       @                              @      �?      $@              @                              �?       @      &@              �?      @      @      (@              �?      @       @              s@      N@     @r@      @@     �J@      =@     @S@      p@     �x@      Q@      T@     �a@     p{@     �u@      $@     �F@      E@     @U@      J@      j@      7@      e@      *@      5@      &@      A@     �i@     �q@      @@     �C@     �O@     r@     `h@              2@      3@      F@      8@      U@      ,@      S@      @      &@      "@      (@     �H@      R@      4@      7@      >@     @[@     �T@              &@      (@      :@      ,@      8@       @      9@               @              @      :@      8@      @      @       @     �L@      @@               @      @      @      $@      @      �?      @                                      �?       @              �?       @      <@      @                              @       @      @                                                      �?      @              �?      �?      3@       @                                               @      �?      @                                              @                      �?      "@      @                              @       @      1@      �?      3@               @              @      9@      0@      @      @      @      =@      :@               @      @               @       @              @              �?              @      @      @      @      @              1@      "@              �?                      @      "@      �?      ,@              �?               @      2@      "@      @       @      @      (@      1@              �?      @              @      N@      (@     �I@      @      "@      "@      @      7@      H@      *@      0@      6@      J@      I@              "@      "@      5@      @      >@       @      0@              @      @      @      @      ,@      �?              @      5@      0@              �?      @      "@              0@              "@                               @       @      @                      @      &@      @                              @              ,@       @      @              @      @      �?      @       @      �?              �?      $@      &@              �?      @      @              >@      $@     �A@      @      @      @      @      2@      A@      (@      0@      1@      ?@      A@               @      @      (@      @      1@      @      *@       @      @      �?      �?      *@      5@              @      $@      0@      &@              @       @       @      �?      *@      @      6@      @      �?      @      @      @      *@      (@      &@      @      .@      7@              @       @      $@      @     @_@      "@      W@       @      $@       @      6@     `c@     �j@      (@      0@     �@@     �f@     @\@              @      @      2@      $@      Z@       @     �T@      @      @      �?      .@     �`@     �f@      &@      ,@      8@     `a@      U@              @      @      (@      @     �T@      @     �R@      @      @      �?      (@     �]@     �d@      @      (@      3@     �Z@     �Q@              @      @      "@      @      ,@      �?      7@                      �?      @      1@      E@       @              @      3@      0@                              �?             @Q@      @     �I@      @      @              @     �Y@     �^@      @      (@      .@     �U@     �K@              @      @       @      @      5@      @       @                              @      0@      2@      @       @      @     �@@      *@              @       @      @      �?      ,@      �?      @                                       @      1@      @               @      9@      (@                      �?       @      �?      @       @      @                              @       @      �?               @      @       @      �?              @      �?      �?              5@      �?      $@      @      @      �?      @      4@      =@      �?       @      "@     �D@      =@              �?       @      @      @      0@      �?               @      @      �?       @       @      @                       @      4@      5@                              �?      �?      &@                       @              �?       @       @      @                       @      4@      4@                              �?      �?      @      �?                      @                              @                                      �?                                              @              $@      �?      �?              @      (@      6@      �?       @      @      5@       @              �?       @      @       @       @              @                               @      �?      @              �?      �?      @      �?                              �?              @              @      �?      �?              @      &@      3@      �?      �?      @      1@      @              �?       @      @       @     �W@     �B@      _@      3@      @@      2@     �E@      J@      [@      B@     �D@     �S@     �b@     �b@      $@      ;@      7@     �D@      <@      @@      *@      ;@      @      @       @      0@      1@     �F@      "@      @      ,@      >@      >@      �?      @       @      "@      @      "@              @              �?              @      @      2@       @               @       @      *@      �?                      @              @                                               @      �?      0@                       @      �?      @                               @              @                                                              @                                       @                               @               @                                               @      �?      &@                       @      �?      �?                                              @              @              �?              �?      @       @       @                      �?      $@      �?                       @                              @                              �?      @      �?                                                                                      @                              �?                       @      �?       @                      �?      $@      �?                       @              7@      *@      5@      @      @       @      *@      &@      ;@      @      @      (@      <@      1@              @       @      @      @      4@      @      4@      @              �?      @      &@      4@      �?       @      $@      ,@      *@               @               @       @      *@      @      4@      @              �?       @      @      *@              �?      "@      "@      *@               @               @       @      @      @                                      @      @      @      �?      �?      �?      @                                                      @      @      �?      @      @      �?      @              @      @      @       @      ,@      @               @       @      @      �?      @      @      �?      @      @              @              @      @      @      �?      @       @               @      �?       @                      @                              �?                      @                      �?      "@       @                      �?      �?      �?     �O@      8@     @X@      (@      <@      0@      ;@     �A@     �O@      ;@      A@      P@      ^@     @^@      "@      7@      5@      @@      9@     �K@      6@     �S@      (@      6@      $@      9@      @@     �K@      1@      9@     �H@     �\@     �\@       @      0@      ,@      8@      6@      3@      $@      K@      @      "@              *@      $@      ?@      "@      2@      @@      G@     �L@       @      @      @      @              @      @      8@              �?              @      @      3@      �?       @      (@      &@      ;@              @      @                      .@      @      >@      @       @               @      @      (@       @      $@      4@     �A@      >@       @                      @              B@      (@      9@      @      *@      $@      (@      6@      8@       @      @      1@      Q@     �L@              *@      $@      3@      6@      A@      &@      1@      @      &@      $@      @      0@      7@       @      @      0@      M@      E@              &@      $@      2@      4@       @      �?       @               @              @      @      �?                      �?      $@      .@               @              �?       @       @       @      2@              @      @       @      @       @      $@      "@      .@      @      @      @      @      @       @      @      �?      �?      @              @      @       @      @      @       @      "@      "@      @      @      @      @      @      @      @      �?      �?      �?              @      @       @      @      �?      @      @      �?      �?      @              @      @      @      �?                      @              �?                               @      �?      @       @      @              @      @      �?       @       @      @      �?      (@                       @                      @       @              @       @      @                              �?              �?      �?      @                                              @      �?                                                                              @              @                       @                              �?              @       @      @                              �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ#,�ohG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKohnh4h7K ��h9��R�(KKo��hu�BH         >                     @�v=<���?�	           ��@                          �2@4?�Q�?�           |�@                           �?ڭ>Y��?�           �@                           �?e_�J�]�?�            �r@                          �1@:!��d�?.            �Q@                           �?�B!Ae�?            �G@������������������������       �B�f��?             ;@������������������������       �{�G�z�?             4@	       
                    �?��,d!�?             7@������������������������       �R���Q�?             $@������������������������       �������?
             *@                           �?�K:y�?�            �l@                          �0@�s3���?S            �`@������������������������       ����K��?             =@������������������������       �>ώ)��?B            �Z@                           @�HΌ���?<            �W@������������������������       �(46a���?1            �R@������������������������       �Ɓ�r�z�?             3@                            �?o�7�W�?!           �{@                           @0�� {�?�             u@                          �0@Rɿ{w��?�            �i@������������������������       ��|�l��?             A@������������������������       ��x9�O�?s            �e@                           �?ߝ�����?X            ``@������������������������       ��2���?/            �P@������������������������       �     ��?)             P@                           @j�n�s��?B            �Y@                           @�BpH��?;            �V@������������������������       �@��Z��?             7@������������������������       �ZP�Q���?,            �P@������������������������       �VUUUUU�?             (@        /                    �?������?�           l�@!       (                    @�ЋB�?&           ��@"       %                   �7@@%w��-�?�           h�@#       $                     �?7�S��Z�?�            �u@������������������������       ��'��4�?�            �q@������������������������       �
��d~�?$            @P@&       '                    �?�7���?�            0q@������������������������       ���<���?.            @Q@������������������������       ����5%��?~            �i@)       ,                    @0��{���?�            �m@*       +                     �?�eP*L��?             6@������������������������       �Y�����?             &@������������������������       ���!pc�?             &@-       .                   �6@����?�             k@������������������������       �ߜc���?T            @`@������������������������       �l�Ӑ���??            �U@0       7                   �6@���n�?�           ��@1       4                   �5@���jxx�?M           �@2       3                    �?tts�Q�?           `{@������������������������       ��q��X�?S             a@������������������������       �4�����?�            �r@5       6                     �?�}S<�[�?@            �Y@������������������������       ��+�@�?�?2            �T@������������������������       ��6��D�?             5@8       ;                   �<@zErMR�?t           �@9       :                     �?eS\���?           }@������������������������       ���QI�?v            �h@������������������������       �'�b�j�?�            �p@<       =                    �?�� �d��?^             b@������������������������       ��q�q�?             8@������������������������       �)9+��]�?M            @^@?       T                    �?�,Q
"�?�           ,�@@       G                   �1@9����U�?�            �@A       F                    @>
ףp}�?0             T@B       C                    �?8�e�?            �I@������������������������       �:/����?             ,@D       E                    �?,��c��?            �B@������������������������       �     ��?             0@������������������������       ������?
             5@������������������������       �&]^z���?             =@H       M                    �?�,V �i�?�           ��@I       J                    �?=��<���?r             e@������������������������       �o��x.�?"            �G@K       L                   �7@���G�q�?P            @^@������������������������       ��7V��?8            �V@������������������������       �,�2���?             ?@N       Q                    �?9�j��W�?            �|@O       P                    �?��4��{�?M             `@������������������������       ��9�Q�a�?&            �N@������������������������       �t�F���?'             Q@R       S                   �4@&�D�\\�?�            pt@������������������������       ��b)0��?=            �W@������������������������       ��e)����?�             m@U       d                   �7@)�M=��?"           �|@V       ]                    �?��%��
�?�            �v@W       Z                    @���*��?W            �a@X       Y                    �?��v���?E            �[@������������������������       ��p���?$             M@������������������������       �d���+��?!             J@[       \                    �?Ӏ����?            �@@������������������������       �ffffff�?             $@������������������������       ����Q��?             7@^       a                    @�s�V��?�            �k@_       `                    �?�Ra����?-            �P@������������������������       �����5�?             =@������������������������       ��e�ݥ��?            �B@b       c                    @�_��?^            �c@������������������������       �=;n,��?5             V@������������������������       � �����?)            @Q@e       j                    @��'�u�?@            @W@f       g                   �9@�N�?�0�?             A@������������������������       �B{	�%��?             "@h       i                    @���Mb�?             9@������������������������       ��|�j��?             .@������������������������       ����(\��?             $@k       l                    @������?%            �M@������������������������       �      �?             0@m       n                    �?#��,�?            �E@������������������������       ��q�q�?             (@������������������������       �V>�� =�?             ?@�t�bh�h4h7K ��h9��R�(KKoKK��h��B�A       �|@     �R@     �u@      <@      Q@      @@     �R@     ؁@     Ђ@     �T@     @S@     `c@     ��@     �y@      &@     �R@      M@     `c@      N@     �t@     �J@     �n@      .@     �B@      "@     �E@     �|@     �}@     �M@     �H@     �Y@     �x@     �p@      @      F@      ;@     �W@     �C@     �V@      @     �@@              @              @     �m@     �d@      @      @      1@     �[@      F@               @      @      ,@       @      C@              $@                              �?     �]@     �L@      �?              @     �H@      *@               @              @       @      3@               @                                      1@      .@                       @      &@       @                               @              ,@              �?                                      .@      @                      �?      @       @                                               @              �?                                      &@      @                               @       @                                              @                                                      @      @                      �?      @                                                      @              �?                                       @       @                      �?      @                                       @              @              �?                                       @      @                              �?                                                       @                                                              @                      �?      @                                       @              3@               @                              �?     @Y@      E@      �?               @      C@      &@               @               @       @      $@              @                                     �Q@      4@                      �?      9@      @                                              @               @                                      4@      �?                              @                                                      @              �?                                     �I@      3@                      �?      6@      @                                              "@              @                              �?      >@      6@      �?              �?      *@      @               @               @       @      @              �?                                      <@      5@      �?              �?      &@       @              �?                       @       @              @                              �?       @      �?                               @      @              �?               @              J@      @      7@              @              @     �]@      [@       @      @      *@      O@      ?@                      @      $@              G@      @      &@              @              @     �T@     �T@       @      @      "@     �K@      4@                      @      $@              9@      @      $@              @               @      E@     �N@       @      @      @      =@      ,@                      �?      @              �?              �?                                      @      8@                              �?      �?                                              8@      @      "@              @               @      B@     �B@       @      @      @      <@      *@                      �?      @              5@      @      �?                               @     �D@      6@                       @      :@      @                       @      @               @      �?      �?                                      9@      &@                      �?      1@      @                                              *@       @                                       @      0@      &@                      �?      "@      @                       @      @              @              (@                              �?      B@      9@                      @      @      &@                                              @              (@                              �?      A@      3@                      @      @      "@                                              @               @                              �?       @      �?                      @      �?       @                                                              @                                      @@      2@                              @      @                                               @                                                       @      @                                       @                                             @n@     �G@     �j@      .@      A@      "@     �B@     �k@     �s@      L@      G@     �U@     �q@      l@      @      E@      8@     @T@     �B@     @\@      4@     �R@      @      "@              $@     @^@     `e@      $@      ;@      3@      a@      W@              *@      @      5@      ,@     �V@      0@     �L@      @       @              $@      L@     �^@      @      3@      .@     @Y@     �P@              &@      @      2@      ,@      K@      �?      8@      @      @              @     �D@     �S@       @      $@      "@     �Q@      ;@               @       @      @      @     �B@      �?      5@      @      @              @      >@      P@       @      @      @     @P@      9@               @       @      @      @      1@              @                                      &@      .@              @      @      @       @                              @              B@      .@     �@@              @              @      .@      F@      @      "@      @      ?@      D@              "@      @      &@      &@      @      @      @                                      @      0@      �?      @      @      .@      @              @      �?      �?       @      =@      (@      =@              @              @      &@      <@      @      @      @      0@     �A@              @      @      $@      "@      7@      @      1@              �?                     @P@      H@      @       @      @     �A@      9@               @              @                              @                                      .@      �?                              �?      �?                                                              @                                      @      �?                                                                                                                                              "@                                      �?      �?                                              7@      @      *@              �?                      I@     �G@      @       @      @      A@      8@               @              @              ,@      �?      @                                     �A@      A@       @      �?      �?      ;@      @                               @              "@      @      @              �?                      .@      *@       @      @      @      @      2@               @              �?              `@      ;@     `a@      (@      9@      "@      ;@      Y@     �a@      G@      3@     �P@      b@     �`@      @      =@      1@      N@      7@     @R@      &@      P@      @      @      �?      $@     @R@     �U@      @       @      8@      J@      S@              $@      @      6@      "@      O@      @      J@       @      @      �?      $@      N@     �S@       @      @      5@      E@     �J@              @      @      2@      "@      4@      @      ;@                              @      @      ,@               @       @      &@      9@              @              $@      @      E@      @      9@       @      @      �?      @      K@     @P@       @      @      *@      ?@      <@              @      @       @      @      &@      @      (@       @      �?                      *@      @      @       @      @      $@      7@              @       @      @              "@      @      @      �?      �?                      *@      @      @       @      �?       @      2@              @       @       @               @              @      �?                                                               @       @      @              �?               @              L@      0@     �R@       @      3@       @      1@      ;@      L@      D@      &@     �E@     @W@      L@      @      3@      &@      C@      ,@     �H@      $@      O@      @       @      @      &@      ;@     �D@      @@      $@      <@     @T@     �E@       @      &@      @      5@      *@      ,@      @      ?@       @      @       @      @      @      "@      &@      "@      5@      ;@      ,@              "@      @      ,@      @     �A@      @      ?@      @      @      �?      @      4@      @@      5@      �?      @      K@      =@       @       @      @      @      @      @      @      *@       @      &@      @      @              .@       @      �?      .@      (@      *@      �?       @      @      1@      �?              @       @               @              �?              @              �?      @              �?              �?              �?              @      @      &@       @      @      @      @              (@       @              (@      (@      (@      �?      @      @      0@      �?      _@      5@     �Y@      *@      ?@      7@      ?@     @\@      _@      7@      <@      J@     �f@     `b@       @      >@      ?@      N@      5@     �Q@      *@      O@      "@      ;@      5@      6@      F@     �Q@      0@      8@      ?@     �Y@     �W@      @      0@      7@     �A@      2@      .@              @              @                      5@      @              �?       @      "@      0@                                              &@              �?              @                      0@      �?              �?      �?      @      (@                                              �?                                                      @                              �?      �?      @                                              $@              �?              @                      "@      �?              �?              @       @                                               @                              @                      @      �?              �?              @       @                                               @              �?                                      @                                              @                                              @              @                                      @      @                      �?      @      @                                             �K@      *@      L@      "@      8@      5@      6@      7@     �O@      0@      7@      =@     �W@     �S@      @      0@      7@     �A@      2@      4@       @      @               @       @      �?      1@      7@      "@      @      @      8@      5@              @      @      (@      @      @              �?              @                      @      @      @       @       @      �?      @              @       @      @       @      .@       @       @               @       @      �?      (@      0@      @       @      @      7@      1@                      @      "@      @      (@      �?       @              �?              �?      $@      ,@      @       @       @      4@      @                      @       @       @      @      �?                      �?       @               @       @                       @      @      $@                      �?      �?      @     �A@      &@     �J@      "@      0@      3@      5@      @      D@      @      3@      7@     �Q@      M@      @      *@      1@      7@      &@      3@       @      1@      @      "@      �?              �?      *@              @      @      9@      "@      �?      @      @      (@       @      *@      �?      @              @                      �?      @               @              *@      @      �?      �?              "@              @      �?      *@      @      @      �?                      @              �?      @      (@       @              @      @      @       @      0@      "@      B@      @      @      2@      5@      @      ;@      @      0@      4@     �F@     �H@      @       @      *@      &@      "@      @              1@                              �?      @      "@      �?      @       @      ;@      *@              �?              $@              (@      "@      3@      @      @      2@      4@      �?      2@      @      $@      2@      2@      B@      @      @      *@      �?      "@      K@       @     �D@      @      @       @      "@     @Q@      K@      @      @      5@     @S@      J@      @      ,@       @      9@      @     �F@       @      ?@      @      @       @      @      Q@     �H@      @      @      2@     �Q@      >@       @      &@      @      .@       @      7@              .@       @       @       @      �?      3@      4@                      @      <@      2@              @              @              0@              .@       @       @       @      �?      (@      2@                      @      5@      (@                              @              $@              $@                       @              $@      *@                               @      @                              �?              @              @       @       @              �?       @      @                      @      *@       @                              @              @                                                      @       @                              @      @              @                               @                                                      �?                                      @      @                                              @                                                      @       @                              @      @              @                              6@       @      0@      �?      �?              @     �H@      =@      @      @      *@      E@      (@       @      @      @      &@       @      @      �?      @                               @      &@       @               @      @      8@       @                               @              @                                                      @      @                       @      (@                                                      �?      �?      @                               @      @      @               @       @      (@       @                               @              2@      �?      $@      �?      �?              �?      C@      5@      @       @      "@      2@      $@       @      @      @      "@       @      ,@      �?      @      �?                              =@      &@                      @      @      @                      @      @       @      @              @              �?              �?      "@      $@      @       @      @      (@      @       @      @               @              "@      @      $@      �?      �?              @      �?      @      @              @      @      6@      �?      @      @      $@      �?      @              @      �?      �?                      �?       @      �?               @              ,@               @              @              @              �?      �?                              �?                                              @                                                               @              �?                               @      �?               @              &@               @              @                               @                                               @      �?               @              @              �?               @                                              �?                                                                      @              �?               @              @      @      @                              @              @       @              �?      @       @      �?      �?      @      @      �?      @      @                                      @              �?                               @                      �?                      �?       @       @      @                               @               @       @              �?      @       @      �?              @      @              �?      �?      �?                                               @       @                      �?      �?                              @              �?      �?      @                               @                                      �?      @      @      �?              @      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��2hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKuhnh4h7K ��h9��R�(KKu��hu�B�         :                   �2@� xţ��?�	           ��@       !                     @�xvC��?�           �@                           �?.9����?�           X�@                            �?�����q�?�             x@                           �?���bKv�?Y            @a@                           �?؉�؉��?            �C@������������������������       ��h$���?	             .@������������������������       ��q�q�?             8@	       
                   �1@�g��Q�??            �X@������������������������       �=�	�:�?%             O@������������������������       �-�R��?            �B@                           �?���`�E�?�            �n@                            �?����l+�?H            �[@������������������������       �������?+            �P@������������������������       ��o��%�?            �F@                           @�g���u�?[            �`@������������������������       �["i�m�?=            @V@������������������������       ��h�d0��?             G@                           @������?�            �t@                          �0@��7��=�?w            `f@                           �?�i��F�?             =@������������������������       �      �?             (@������������������������       ��������?             1@                          �1@JvNd��?c            �b@������������������������       �E�r*e�?2            �R@������������������������       �����p9�?1             S@                           @?�ƨ�?^             c@                           @�N贁�?K             ^@������������������������       �:J�����?              J@������������������������       �\��M��?+             Q@                             �?     ��?             @@������������������������       ��>4և��?
             ,@������������������������       �n�����?	             2@"       /                    �?����Ay�?�            ps@#       *                    @�$�#n�?Z             a@$       '                    @�mM`���??             W@%       &                    �?�[��Y��?0            @R@������������������������       �-C��6�?             9@������������������������       ���8����?             H@(       )                    �?~�Q���?             3@������������������������       ��T�x?r�?	             &@������������������������       �      �?              @+       ,                     @M�lRT�?            �F@������������������������       �������?             1@-       .                    @4և����?             <@������������������������       �ҳ�wY;�?             1@������������������������       �b���i��?             &@0       7                    @9B�-8��?r            �e@1       4                   �1@Y�BS��?Y            �a@2       3                    @�"?Uz��?3            �T@������������������������       �~X�<��?             B@������������������������       �dbOs�U�?            �G@5       6                    @��gS~Y�?&             M@������������������������       �<��b��?            �D@������������������������       �躍`3�?             1@8       9                    @���+	�?            �@@������������������������       ��ˠT�?             6@������������������������       ��x?r���?	             &@;       Z                    �?�ޟK���?�           ��@<       K                    �?����3�?(           x�@=       D                    �?H&<�6��?N           ��@>       A                   �3@�~ ��?v            �h@?       @                    �?�Ӫ�Ep�?             7@������������������������       ��<ݚ�?             "@������������������������       �������?	             ,@B       C                    @���h��?g            �e@������������������������       ��5�1	�?O            �a@������������������������       �Er����?             A@E       H                    @Qi�9��?�            u@F       G                     �?��1^��?�            �i@������������������������       �q�F�:�?=             W@������������������������       �*x9/g�?F             \@I       J                     @H�7C��?U            �`@������������������������       ���U�Ɓ�?)            �Q@������������������������       ����5��?,            �O@L       S                     �?~j60��?�           @�@M       P                    @^�q�VR�?           �{@N       O                   �6@�L�q`�?t            `g@������������������������       �CkR�W�?>            �X@������������������������       �
�g����?6            @V@Q       R                     �?��l(��?�            �o@������������������������       �Fs�e��?H            �`@������������������������       �}���k�?P            @^@T       W                    @z�FG[��?�            �t@U       V                   �4@�0�ͺ��?�            �h@������������������������       ���߭Q�?4            �T@������������������������       ���io�?N             ]@X       Y                    @ڤ�:�^�?L            �`@������������������������       �?��M��?:            �Y@������������������������       �     P�?             @@[       h                    �?���z�H�?�           ��@\       a                    �?d��\h�?�           ��@]       `                   �?@�����?�             o@^       _                    @v�w���?�            �m@������������������������       �ko��DE�?Z            �a@������������������������       �!�!���?8            @X@������������������������       �{�G�z�?             $@b       e                    �?��0��k�?@           �@c       d                   �;@ ����?R            �a@������������������������       ��������?H            @]@������������������������       �UUUUUU�?
             8@f       g                   �8@�����;�?�            �v@������������������������       �U=ޭ���?�            �h@������������������������       ���k�D��?h            @e@i       p                     �?˿K���?�           ��@j       m                     �?��u����?           p{@k       l                    @�<��%�?�            �j@������������������������       ���O�4A�?s            @g@������������������������       ��q-�T�?             :@n       o                   �9@��G���?�            `l@������������������������       ���-w�~�?            �h@������������������������       �/����?             <@q       t                   �?@o��ɹ�?�            �w@r       s                    @�'j�q��?�            w@������������������������       ��/�Bʊ�?�            �k@������������������������       �xCͯO�?V            �b@������������������������       ��8��8��?	             (@�t�bh�h4h7K ��h9��R�(KKuKK��h��BxE       �~@      R@     0t@      A@     �Q@      ?@     @U@     �@     Ȃ@      Q@     �R@     �e@     �@     {@      &@     �N@     �G@     @_@     �K@     �a@       @     �J@      �?       @              &@     0q@      h@      @      "@      5@     �g@      S@              "@      @      4@      @     @U@      @      6@              �?               @     �k@     �c@      @       @      ,@      _@     �G@              @      �?      "@       @     �D@      @       @                              @     `b@     @U@      �?      @      "@      N@      7@                              �?              ,@      @      �?                                     �G@      B@                      @      ;@      @                              �?              @       @                                              $@      @                      �?      ,@      @                                               @                                                      @      �?                              @      @                                              @       @                                              @      @                      �?      &@                                                      "@      �?      �?                                     �B@      @@                       @      *@      @                              �?              @                                                      ?@      4@                              @                                      �?              @      �?      �?                                      @      (@                       @      @      @                                              ;@              @                              @      Y@     �H@      �?      @      @     �@@      1@                                              (@              @                                     �K@      1@                       @      1@      @                                              @              �?                                     �C@      @                       @      $@      @                                              @               @                                      0@      (@                              @      �?                                              .@              @                              @     �F@      @@      �?      @      @      0@      (@                                              "@               @                              @      C@      2@              @       @      @       @                                              @               @                                      @      ,@      �?               @      $@      @                                              F@       @      ,@              �?              @      S@     �Q@      @      @      @      P@      8@              @      �?       @       @      <@      �?      $@              �?              @      ?@      ?@      @      @       @     �D@      ,@               @              @       @       @                                                       @      @                              @      �?                                              @                                                      @                                      �?      �?                                               @                                                      @      @                              @                                                      4@      �?      $@              �?              @      7@      8@      @      @       @      B@      *@               @              @       @       @      �?      @              �?              @      .@      &@              @       @      1@      @                                       @      (@              @                               @       @      *@      @                      3@      @               @              @              0@      �?      @                                     �F@      D@                      @      7@      $@              @      �?      @              ,@      �?      @                                      E@      A@                      @      ,@      @               @              �?              @              @                                      9@      *@                              @      �?                                               @      �?                                              1@      5@                      @      $@      @               @              �?               @              �?                                      @      @                              "@      @               @      �?      @              �?                                                       @      �?                               @      �?               @      �?      @              �?              �?                                      �?      @                              @      @                                              L@      @      ?@      �?      @              @      J@      B@      �?      �?      @     �P@      =@              @       @      &@      �?      :@       @      "@                              �?     �@@      &@      �?              @      A@      $@               @              @              .@       @      �?                              �?      1@       @      �?              @      ;@      $@               @              @              .@       @                                      �?      .@      �?                      @      6@      "@              �?               @              @       @                                              �?                              @      @      @              �?              �?               @                                              �?      ,@      �?                      �?      1@      @                              �?                              �?                                       @      @      �?                      @      �?              �?              �?                              �?                                       @      @                               @      �?              �?              �?                                                                              @      �?                      @                                                      &@               @                                      0@      @                              @                                                                      @                                      @       @                              @                                                      &@               @                                      (@      �?                               @                                                      @                                                      &@                                                                                              @               @                                      �?      �?                               @                                                      >@      �?      6@      �?      @               @      3@      9@              �?       @     �@@      3@              �?       @       @      �?      <@      �?      .@      �?      @                      @      6@              �?       @      <@      2@              �?       @      @      �?      2@      �?      $@              @                      @      *@                       @      $@      ,@              �?       @      �?              @      �?                      @                      @       @                       @      @      @                                              &@              $@              �?                      �?      @                              @      &@              �?       @      �?              $@              @      �?                              @      "@              �?              2@      @                              @      �?      @              @      �?                               @       @                              2@      �?                              �?              @                                                      �?      �?              �?                      @                              @      �?       @              @                               @      (@      @                              @      �?                              �?               @              @                               @      @                                      @      �?                                                                                                      @      @                               @                                      �?             �u@      P@     �p@     �@@      O@      ?@     �R@     �p@     �y@     �O@     �P@     @c@     0z@     Pv@      &@      J@      F@     @Z@      J@     �e@      1@     @\@      @      0@      @      5@     `d@     �n@      3@      :@      F@     `j@     �b@       @      1@      *@     �G@      7@      R@       @     �K@       @      "@      @      .@     �@@     @R@      @      (@      .@     �V@     �Q@       @      @      $@      =@      5@      8@      @      ,@              �?       @      �?      1@      B@      @      @       @      D@      A@              �?       @      @      @      @                                                      @      @                              �?      @                                               @                                                      �?      @                                       @                                              @                                                      @      �?                              �?      @                                              3@      @      ,@              �?       @      �?      (@      ?@      @      @       @     �C@      ;@              �?       @      @      @      0@      @      ,@              �?       @      �?       @      =@      @      @       @      7@      5@              �?       @      @      @      @                                                      @       @                              0@      @                               @      �?      H@      @     �D@       @       @       @      ,@      0@     �B@              "@      *@      I@     �B@       @      @       @      8@      0@     �C@       @      4@              @      �?      @      &@      .@              @      @     �@@      5@              @      @      5@       @      0@       @      $@              �?              @      @      @              @      @      1@      @               @              .@              7@              $@              @      �?              @      &@              �?      @      0@      ,@              @      @      @       @      "@       @      5@       @      @      �?      $@      @      6@              @      @      1@      0@       @              �?      @       @      @       @      0@               @              @       @      .@               @              @      $@                      �?       @      @      @              @       @      �?      �?      @      @      @               @      @      (@      @       @                      �?       @     �Y@      "@      M@       @      @      �?      @     @`@     `e@      *@      ,@      =@     @^@      T@              $@      @      2@       @     @P@      @      B@      �?                      @      M@     �[@       @       @      ,@      P@     �K@               @      �?      "@       @      9@      @      ,@                              @      4@     �N@      @              @      =@      0@                              @              (@              @                              @      "@     �D@      �?              @      2@      @                              �?              *@      @      $@                                      &@      4@      @                      &@      &@                              @              D@      �?      6@      �?                              C@     �H@      @       @      &@     �A@     �C@               @      �?       @       @      2@      �?      &@                                      0@      9@      @      �?       @      6@      9@               @              �?              6@              &@      �?                              6@      8@              @      @      *@      ,@                      �?      �?       @     �B@      @      6@      �?      @      �?       @      R@     �N@      @      @      .@     �L@      9@               @       @      "@             �A@       @      "@      �?       @      �?      �?      D@      I@       @      @      @      9@      2@              @              �?              1@              �?                      �?              7@      ,@      �?              @       @      &@               @              �?              2@       @       @      �?       @              �?      1@      B@      �?      @              1@      @              @                               @       @      *@              @              �?      @@      &@      @      @      &@      @@      @              @       @       @               @       @       @                                      <@       @      @      @      @      9@      @              @       @      @                              @              @              �?      @      @                      @      @                                      @              f@     �G@     �c@      =@      G@      :@     �J@     �Z@     �d@      F@      D@     �[@      j@     �i@      "@     �A@      ?@      M@      =@     �Q@      9@     �T@      ,@      :@      3@      ;@      9@      I@      8@      @@     @Q@     �T@     @]@      @      5@      4@      :@      5@      4@      @      8@              *@              @       @      1@      @      ,@      @@      G@      >@              @      @      $@      @      4@      @      8@              (@              @       @      1@      @      &@      ;@      G@      >@              @      @      "@      @      @      @      1@              "@              �?      @      .@              @      .@     �@@      0@              @      @      @       @      *@      @      @              @              @      �?       @      @      @      (@      *@      ,@              �?       @      @      @                                      �?                                              @      @                                              �?              I@      2@     �M@      ,@      *@      3@      4@      1@     �@@      4@      2@     �B@     �B@     �U@      @      1@      ,@      0@      ,@      6@      @      4@      @      @       @              $@      ,@      @              "@      (@      *@      �?      �?       @      @      @      4@      @      &@      @      @      @              $@      *@      @              "@      (@      *@      �?      �?      @      @      �?       @              "@              �?      @                      �?       @                                                      @               @      <@      .@     �C@      &@      "@      &@      4@      @      3@      ,@      2@      <@      9@     �R@      @      0@      @      (@      &@      4@       @      5@       @      @      @      "@      @      (@      @      "@      @      .@      L@              @              "@      @       @      @      2@      "@      @      @      &@              @      &@      "@      6@      $@      2@      @      (@      @      @      @     �Z@      6@     �R@      .@      4@      @      :@     �T@     �\@      4@       @     �D@     @_@     @V@      @      ,@      &@      @@       @     �L@      @      C@      $@      @      @       @      J@     @R@      .@       @      5@      I@      K@              @       @      1@      @      ;@      @      5@       @       @      @      @      ;@      8@       @      @      (@      :@      1@              @      @      *@      �?      0@      @      1@      @      �?      @      @      9@      7@       @      @      &@      6@      0@              @      @      *@      �?      &@              @      �?      �?                       @      �?                      �?      @      �?                                              >@       @      1@       @      @      �?      �?      9@     �H@      @      @      "@      8@     �B@               @      @      @      @      =@      �?      &@       @      �?              �?      7@     �H@      @      @      "@      6@      @@                      @      �?      @      �?      �?      @              @      �?               @              �?      �?               @      @               @              @              I@      0@      B@      @      ,@      @      2@      >@      E@      @              4@     �R@     �A@      @      @      @      .@      @     �H@      *@      ?@      @      ,@       @      2@      >@     �D@      @              4@     �R@     �A@      @      @      @      .@      @      7@      @      0@      @      $@       @      $@      7@      @@      @              2@     �E@      4@               @               @       @      :@      $@      .@              @               @      @      "@       @               @      @@      .@      @      @      @      @      �?      �?      @      @                      �?                      �?                                              �?                                �t�bub�r     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJՠ"QhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKqhnh4h7K ��h9��R�(KKq��hu�B�         @                     @�K�Cy��?�	           ��@       !                   �3@��~��C�?�           ʥ@                          �1@����*�?�           ��@                           @*�4���?           �{@                           @�L��Ա�?�             j@                           �? ��q�=�?n            �d@������������������������       ��v�,��?5            �S@������������������������       �ڦs@�?9            @U@	       
                    �?��aC��?            �F@������������������������       ��q�q�?	             (@������������������������       �`�[9��?            �@@                            �?x�	[��?�            �l@                           �?}�"��X�?b            �c@������������������������       �|�<�ւ�?7            �U@������������������������       �Е�܈I�?+            �Q@                           �?�u�C���?/            �R@������������������������       ��lev��?            �D@������������������������       ��x��6�?            �@@                           �?�,����?g           ��@                          �2@:ǖt��?c            �a@                           �?$����?:            �V@������������������������       ��(\����?             D@������������������������       �"6J^r��?"            �I@                           @;�;��?)             J@������������������������       �K~���?             >@������������������������       �L�9���?             6@                           @�(l��W�?            {@                           �?�Ć���?t            �f@������������������������       �+���{�??            �Y@������������������������       �_���D�?5            @T@                            @�9U�Fo�?�             o@������������������������       �A�� ;�?w            �i@������������������������       ������?             F@"       1                    �?<Ӿ�#��?o           ��@#       *                    �?�Z��5K�?�            �@$       '                   �<@ThSy$�?�            �o@%       &                     �?|��?y��?�            �j@������������������������       ����Sn�?|            �g@������������������������       ��A`��"�?             9@(       )                   �=@�j">���?            �D@������������������������       �Z�eY�e�?             5@������������������������       �)\���(�?             4@+       .                   �5@�d��6�?            z@,       -                    �?�]�`��?>             Z@������������������������       ���|���?             F@������������������������       ��h$���?#             N@/       0                    �?;�=�=�?�            �s@������������������������       �=<��\��?<            �U@������������������������       ���7+�?�            `l@2       9                   �:@�Y��Z�?�           8�@3       6                    @��g��?D           ��@4       5                    @|���t��?�             j@������������������������       �Z��:�r�?            `h@������������������������       �3�E��?             *@7       8                    @�M��?�           @�@������������������������       ����|��?%           �}@������������������������       �:�8�?z�?�            `m@:       =                    �?X����6�?u            �f@;       <                    �?�������?$            �M@������������������������       �x�"w���?             3@������������������������       ��p=
ף�?             D@>       ?                    �?�(w.6.�?Q            �^@������������������������       ��A�%���?!            �J@������������������������       �#���d��?0            �Q@A       `                   �6@�{dp��?�           ��@B       Q                    �?��.��N�?�            �@C       J                    @PR�/���?�            `v@D       G                    �?0�F�i}�?�            �k@E       F                    �?�cԧ���?J            @[@������������������������       �~4��?"            �J@������������������������       ��$I�$I�?(             L@H       I                    �?N;����?L            @\@������������������������       ��#Vn\1�?!             G@������������������������       ����-n��?+            �P@K       N                    @��¤��?Z             a@L       M                   �3@�����?            �G@������������������������       �~X�<��?             2@������������������������       ����;\I�?             =@O       P                    �?U��cV�?=            @V@������������������������       �F%u��?             9@������������������������       �     p�?*             P@R       Y                   �1@�P��?�            �u@S       V                    �?��+&�?>            �X@T       U                    @�;�;�?              J@������������������������       ��q-�T�?             :@������������������������       ��"AM��?             :@W       X                    �?�x���?             G@������������������������       �4%���?             1@������������������������       ��;N��?             =@Z       ]                    �?��η�?�             o@[       \                   �2@!�;^�/�?K            �_@������������������������       �1��D�\�?            �C@������������������������       ���U���?7            �U@^       _                    @� �0�?O            �^@������������������������       �i -�k��?4            �T@������������������������       ����|�l�?            �C@a       p                   �@@m'~WȌ�?           @z@b       i                   �9@<�xh�?�            �x@c       f                    @٩�/�?�            @i@d       e                    �?=C���?`            �a@������������������������       ����Q��?)             N@������������������������       �L�`D�?�?7            �T@g       h                   �7@���*�?#             N@������������������������       ���S�r
�?             <@������������������������       �     ��?             @@j       m                    �?��<��4�?t            �h@k       l                   �;@��`d���?2            �U@������������������������       �,r�|��?             C@������������������������       �UUUUU��?             H@n       o                   �>@�w#����?B            �[@������������������������       �UUUUUU�?9             X@������������������������       ��|�j��?	             .@������������������������       �u���?             5@�t�bh�h4h7K ��h9��R�(KKqKK��h��BC       p}@     @U@     �v@     �B@      S@      3@     �Q@     �@     x�@     �K@     �X@     �b@     ��@     py@      &@     �M@      D@     `c@     �M@      u@     �J@     �m@      6@      G@      @      I@     |@     �@     �D@     �P@     �X@     �y@     pp@      �?      D@      9@      Y@     �@@     @_@      $@     �J@       @       @              @     �q@     �m@      @      "@      3@      c@      T@              @       @      0@       @      K@      @      *@                              @     `a@     �]@              @      "@     �R@      0@                               @      �?      4@      @      "@                              @     �J@      O@              @      @      B@      $@                              �?      �?      3@      @       @                              @      G@     �A@              @      @      ?@      @                              �?      �?      .@       @      @                               @      6@      4@               @              $@                                              �?      @       @      @                              �?      8@      .@              @      @      5@      @                              �?              �?              �?                                      @      ;@                              @      @                                              �?                                                      @      @                               @      �?                                                              �?                                       @      8@                              @      @                                              A@      �?      @                                     �U@     �L@                      @      C@      @                              �?              ;@      �?      @                                     �J@     �B@                      @      ?@                                      �?              ,@              @                                      B@      ,@                      @      0@                                                      *@      �?                                              1@      7@                      �?      .@                                      �?              @              �?                                     �@@      4@                              @      @                                              �?                                                      6@      &@                               @      @                                              @              �?                                      &@      "@                              @      �?                                             �Q@      @      D@       @       @              @     �b@     �]@      @      @      $@     �S@      P@              @       @      ,@      �?      6@      @      1@                                      6@      9@      @       @      @      9@      0@              �?               @      �?      (@       @      *@                                      ,@      2@       @              @      4@      @                              �?               @              @                                      @      @                      �?      @      @                              �?              @       @      @                                       @      (@       @               @      *@       @                                              $@      �?      @                                       @      @      �?       @      �?      @      $@              �?              �?      �?      @      �?      @                                      @      @                              @      @              �?                              @                                                      @      �?      �?       @      �?      �?      @                              �?      �?     �H@       @      7@       @       @              @     �_@     �W@      @       @      @     �J@      H@              @       @      (@              *@              @                              @      I@      G@                      @      ;@      ?@              �?      �?                      @              @                                      <@     �A@                      @      .@      *@                                              "@              @                              @      6@      &@                      �?      (@      2@              �?      �?                      B@       @      0@       @       @              �?      S@      H@      @       @       @      :@      1@               @      �?      (@              ;@       @      *@       @                             �P@      D@      @       @      �?      0@      1@               @      �?      (@              "@              @               @              �?      $@       @                      �?      $@                                                     �j@     �E@     @g@      4@      F@      @     �E@     @d@     �p@      A@     �L@     �S@     @p@     �f@      �?      B@      7@      U@      ?@     @T@      8@     �V@      $@      5@      �?      7@      >@      O@      *@      >@     �A@     �T@     �R@              9@      &@     �B@      7@      =@      $@      9@      �?      @              $@      *@     �A@      @      *@      ,@     �E@      3@              @      @      &@      (@      <@      @      4@      �?      @               @      *@      ?@       @      &@      &@      E@      1@              @       @      $@      "@      ;@      @      .@      �?      @               @       @      :@      �?       @      $@      D@      .@              @       @      $@      "@      �?              @                                      @      @      �?      @      �?       @       @                                              �?      @      @              @               @              @       @       @      @      �?       @              �?      �?      �?      @      �?      @      �?                               @              @      �?                      �?                              �?               @              �?      @              @                              �?      �?       @      @               @              �?              �?      �?      J@      ,@     @P@      "@      ,@      �?      *@      1@      ;@      "@      1@      5@     �C@     �K@              4@       @      :@      &@      3@              $@              �?               @      (@      *@              �?      @      .@      .@               @               @       @      &@              @              �?                      @      �?              �?      �?      *@      @               @               @               @              @                               @      @      (@                      @       @      (@                              @       @     �@@      ,@     �K@      "@      *@      �?      &@      @      ,@      "@      0@      1@      8@      D@              2@       @      2@      "@      1@       @      (@      �?      @              @      �?      @      @      @      @      @      "@              @      �?      @              0@      (@     �E@       @       @      �?       @      @      @      @      &@      *@      1@      ?@              .@      @      &@      "@     �`@      3@      X@      $@      7@      @      4@     �`@      j@      5@      ;@      F@     @f@     @[@      �?      &@      (@     �G@       @     �\@      ,@     �R@       @      .@       @      0@     �]@     �h@      $@      8@      @@     �c@     �T@      �?      @      @      B@      @      5@      @      0@       @      �?       @      "@      (@     �J@      @      @      "@      A@      :@              @              @              4@      @      *@                       @       @      (@     �J@      @      @      "@      ?@      :@              @              @              �?              @       @      �?              �?                               @              @                                                     @W@      &@      M@      @      ,@              @     �Z@      b@      @      3@      7@     �^@      L@      �?      @      @      =@      @     �M@       @      A@      @      @              @     �S@     �Z@      @      ,@      .@     �U@     �A@      �?      @      @      .@      @      A@      @      8@      @      &@              @      <@      C@       @      @       @     �A@      5@              �?       @      ,@       @      2@      @      6@       @       @      �?      @      *@      (@      &@      @      (@      6@      ;@              @      @      &@       @               @      @       @      �?              �?       @       @      @      �?      �?      &@      *@                      @      �?                              @              �?              �?       @                              �?      @      �?                                                       @      @       @                                       @      @      �?              @      (@                      @      �?              2@      @      .@              @      �?      @      @      $@      @       @      &@      &@      ,@              @       @      $@       @      "@      �?      @              @                      @      �?      @       @      @      @      $@               @              @      �?      "@       @      &@              �?      �?      @              "@       @               @       @      @               @       @      @      �?     �`@      @@     �^@      .@      >@      .@      5@      W@     �\@      ,@      @@      I@      g@      b@      $@      3@      .@     �K@      :@     �X@      .@     �Q@      @      $@      @      @      T@     �T@      @      2@      6@      a@     @V@              (@      @      A@       @     �E@      &@     �C@      @      "@      @      �?      :@      B@      @      $@      .@     �O@     �H@              &@      @      ;@      @      <@      "@      1@      �?      @      �?      �?      7@      5@              "@      @      G@      ;@              @      �?      ,@      @      3@      @      @              @                       @      .@              @      @      0@      *@              @               @       @      $@      �?       @              @                      @      @                      �?      @      &@               @              @              "@      @      @              @                       @      $@              @       @      $@       @               @               @       @      "@      @      $@      �?      �?      �?      �?      .@      @              @      @      >@      ,@              @      �?      @      �?       @              �?                      �?      �?      (@      @                      @      *@      @                      �?      �?      �?      @      @      "@      �?      �?                      @       @              @      �?      1@       @              @              @              .@       @      6@       @       @       @              @      .@      @      �?       @      1@      6@              @      @      *@      �?      @              ,@                      �?                                              @      @      "@              @      @      @              �?              �?                                                                      �?       @      @              @       @      @              @              *@                      �?                                               @       @      @                      �?                      "@       @       @       @       @      �?              @      .@      @      �?      @      *@      *@                      �?      $@      �?      @               @                                              @       @                      @      �?                      �?      @      �?      @       @      @       @       @      �?              @      "@      �?      �?      @      "@      (@                              @              L@      @      ?@      @      �?              @      K@      G@      @       @      @     �R@      D@              �?      �?      @      @      .@              @                                      3@      ;@              �?      @      2@      "@                              �?              &@              @                                      &@      ,@                              &@       @                                              @               @                                       @      @                              @                                                       @              �?                                      @       @                              @       @                                              @               @                                       @      *@              �?      @      @      @                              �?              @               @                                              @                      @      @      �?                                              �?                                                       @      "@              �?              @      @                              �?             �D@      @      :@      @      �?              @     �A@      3@      @      @      @      L@      ?@              �?      �?      @      @      5@              .@                              �?      6@      $@      @      @      �?      =@      0@                      �?       @              (@              $@                                      $@      �?                              @      @                                              "@              @                              �?      (@      "@      @      @      �?      :@      *@                      �?       @              4@      @      &@      @      �?              @      *@      "@               @      @      ;@      .@              �?              @      @      $@      @      &@       @      �?              @      @      @               @       @      5@      *@                              @       @      $@                      �?                      �?      $@      @                      �?      @       @              �?              �?       @      A@      1@      J@      "@      4@      (@      ,@      (@      @@       @      ,@      <@      H@     �K@      $@      @      "@      5@      2@      A@      1@      J@      "@      0@      $@      ,@      (@      @@       @      ,@      8@      H@     �K@      @      @      "@      5@      .@      5@      @      =@       @      @      @       @      "@      9@      @      @      *@      ,@      >@      @              @      (@       @      .@       @      $@       @      @      @      @      @      9@      @      @      @      (@      7@       @              @      $@       @      @              @              �?      @              @      $@                               @      2@                      �?      @              $@       @      @       @      @              @       @      .@      @      @      @      @      @       @              @      @       @      @       @      3@              �?              @      @                       @      @       @      @       @              @       @               @              $@              �?                      @                       @       @       @      @       @                                      @       @      "@                              @                                      @              @                      @       @              *@      *@      7@      @      "@      @      @      @      @       @       @      &@      A@      9@              @       @      "@      *@      &@      @      "@      @      @                              @              @      @      8@      $@               @              �?      @      @      @      �?      @                                      @                      @      .@       @              �?              �?      @       @      �?       @              @                              �?              @       @      "@       @              �?                       @       @      "@      ,@      @      @      @      @      @      @       @      @      @      $@      .@              @       @       @       @       @      "@      ,@       @      @      @      @      @       @      �?      @      @      $@      &@              �?       @       @       @                               @              @                      �?      �?              �?              @               @                                                              @       @                                              @                      @       @                      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��|hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKihnh4h7K ��h9��R�(KKi��hu�B�         <                    �?Ћ2z���?�	           ��@       !                   �2@w6�c���?R           ��@                            @*��ԟR�?D           �@                           �?4FM0�'�?�            pw@                            �?6r3֛��?q            �f@                          �1@�E����?)             R@������������������������       ������?             F@������������������������       �����>�?             <@	       
                    @(�ŚR�?H            �[@������������������������       ���nk�?<             W@������������������������       �����p9�?             3@                           �?�q�e�?|             h@                           @�����?             7@������������������������       ���Q��?             $@������������������������       ��T�6|��?             *@                           @:?R��3�?o             e@������������������������       �~e�.y0�?$             J@������������������������       �4��f��?K            @]@                           @�����*�?W             `@                           �?���k(�?7             S@                          �1@�ٔ_���?)             M@������������������������       ��r
^N��?             <@������������������������       ��z�G��?             >@                          �1@��"e���?             2@������������������������       �Y�����?             &@������������������������       �������?             @                          �1@���U�?             �J@                            @|�j�Y��?             >@������������������������       ��1G����?             *@������������������������       �J,�ѳ�?
             1@                            @��+7��?             7@������������������������       ��(\����?             $@������������������������       �����W�?             *@"       1                     @�<ƍ(>�?           ��@#       *                    �?�0��}��?1           ��@$       '                   �7@6����?�            �r@%       &                   �6@�aS���?�            �j@������������������������       ��DIǽ��?t            `e@������������������������       ��N8���?             E@(       )                    �?��i�V��?;             V@������������������������       �4%���?             1@������������������������       �C�k��-�?-            �Q@+       .                    @��p8�?h           X�@,       -                   �4@�'�h�?�            `p@������������������������       ��5�u���?.            �S@������������������������       ���H�?r             g@/       0                    @(��3��?�            Pt@������������������������       �>vO5�?\            �c@������������������������       ��L�p�?l             e@2       9                    @zN ����?�            `w@3       6                   �6@^q���r�?�            u@4       5                    �?�v�x���?m            �f@������������������������       �$ ;�_��?;            �W@������������������������       �q"ԅ7��?2            @U@7       8                    �?^��P��?_            �c@������������������������       �lx5C��?&            �O@������������������������       �.���?9            �W@:       ;                    �?�����?            �B@������������������������       ���D���?
             5@������������������������       �     ��?             0@=       P                    �?���Q�?L           Ơ@>       G                    @n��5���?w           ��@?       @                   �0@�Þ����?           �{@������������������������       ���8��8�?             8@A       D                    @`e�Z#	�?
           pz@B       C                     �?�����?�            Pw@������������������������       ������?}            �h@������������������������       ��Ra��H�?m             f@E       F                   �7@-�����?              I@������������������������       �q-�lJ��?            �B@������������������������       �������?             *@H       K                   �2@�d���?`            �c@I       J                    @t�1s^1�?            �G@������������������������       ��V�߻�?             ;@������������������������       �q=
ףp�?             4@L       M                   �3@��꒸�?D            �[@������������������������       �9��8���?             (@N       O                   �4@;��/��?<            �X@������������������������       �V}��b�?             9@������������������������       ��MN�6�?,            @R@Q       \                   �5@�v��&�?�           �@R       Y                    @H��$�K�?�           ��@S       V                    @pt�]�=�?�           ��@T       U                     @B�N;�V�?E           �~@������������������������       ����Y��?�            q@������������������������       ����AM�?�             k@W       X                     �?b��?�            �p@������������������������       ���|��y�?a            �c@������������������������       ��*���?H            �[@Z       [                     �?8�Z$��?             :@������������������������       �      �?             0@������������������������       �ffffff�?             $@]       b                    �?�۸�w�?�           ��@^       a                     �?���v	��?.            @Q@_       `                     �?7��d��?             A@������������������������       ��t����?             1@������������������������       ��?�0�!�?             1@������������������������       �j]���~�?            �A@c       f                     @aw�����?�           ��@d       e                   �>@�l�Nr\�?!           }@������������������������       ����g6�?           @z@������������������������       ��o1�?             �F@g       h                    �?h�����?�             l@������������������������       �n��e'�?[             c@������������������������       �N������?/            �Q@�t�bh�h4h7K ��h9��R�(KKiKK��h��BX>       }@     �T@     `u@     �A@     �L@      >@     �W@     ��@     P�@     �P@      V@     `e@     0�@      {@      ,@     �L@     �F@     @b@     �K@     �m@      9@      `@      @      .@      $@     �B@     0t@     0t@      ,@     �A@     �K@     �r@     �d@              5@      *@     �G@      .@      O@      @      <@                              @      f@     �Z@      �?      @       @      R@      <@              �?              @              D@      @      (@                              @     �b@     �V@              @      @      H@      2@                                              3@              @                                     �V@      C@               @      @      0@      $@                                               @              @                                      =@      3@               @       @      @      @                                              @              @                                      6@      "@               @       @               @                                              @                                                      @      $@                              @      @                                              &@              �?                                      O@      3@                      �?      (@      @                                              @              �?                                     �K@      .@                      �?      (@       @                                              @                                                      @      @                                      @                                              5@      @       @                              @     �L@      J@              �?      @      @@       @                                                              �?                                      @      @              �?      �?      &@                                                                                                              @      @                      �?      �?                                                                      �?                                              �?              �?              $@                                                      5@      @      @                              @     �J@     �G@                       @      5@       @                                              "@      @      @                                      (@      4@                              @      �?                                              (@       @      @                              @     �D@      ;@                       @      1@      @                                              6@      �?      0@                              �?      <@      0@      �?               @      8@      $@              �?              @              0@      �?      @                              �?      &@       @      �?               @      2@      @              �?              @              (@      �?      @                              �?      $@      @      �?               @      &@      @              �?              @              &@              �?                                       @      �?      �?              �?      @       @                                              �?      �?      @                              �?       @       @                      �?       @      @              �?              @              @                                                      �?      @                              @      �?                                              �?                                                              @                              @                                                      @                                                      �?      �?                              �?      �?                                              @              (@                                      1@       @                              @      @                                              @              @                                      &@      @                              @       @                                                              �?                                      @      @                              @                                                      @              @                                       @                                               @                                               @               @                                      @       @                              @       @                                              �?               @                                      @       @                               @                                                      �?              @                                      @                                      �?       @                                              f@      3@     @Y@      @      .@      $@      ?@     `b@      k@      *@      @@     �G@      l@     @a@              4@      *@      D@      .@     �^@      *@     �R@       @      @              ,@      \@     �f@      "@      :@      ?@     �b@      V@              *@      @      @@       @     �B@      @      :@                              @     �@@     @V@      @      "@      2@      I@      5@               @              @      �?      4@      @      6@                              �?      7@     �O@      @      @      0@     �D@      .@                              �?              .@      @      2@                              �?      4@      M@              �?      $@      ?@      *@                              �?              @       @      @                                      @      @      @       @      @      $@       @                                              1@              @                              @      $@      :@              @       @      "@      @               @               @      �?      �?                                                      �?      @              @              @      �?                              �?      �?      0@              @                              @      "@      6@              �?       @      @      @               @              �?             �U@       @     �H@       @      @              $@     �S@     @W@      @      1@      *@     �X@     �P@              &@      @      =@      @      :@      @      ;@      �?      @              @      C@      F@       @      $@       @     �@@      B@              "@      �?      0@       @      &@      @              �?                              @      7@      �?       @       @      .@      @              @              @              .@              ;@              @              @      ?@      5@      �?       @      @      2@      ?@              @      �?      (@       @      N@      @      6@      �?      @              @     �D@     �H@      @      @      @     �P@      ?@               @      @      *@      @     �C@      @      "@               @              @      @      :@              @      �?     �@@      @               @      @      (@      @      5@      �?      *@      �?      �?              @      A@      7@      @      @      @     �@@      8@                              �?      �?     �J@      @      :@      �?      "@      $@      1@     �A@     �A@      @      @      0@      S@      I@              @       @       @      @      I@      @      :@      �?      @      $@      @      @@      A@      @      @      ,@      P@      I@              @      @      @      @      8@              @      �?      @      @              =@      ,@       @      @      @     �C@      @@              @      �?      @      @      $@              @      �?      @       @              "@      $@              @      @      5@      3@                      �?      �?      @      ,@              �?                      @              4@      @       @      �?       @      2@      *@              @              @              :@      @      4@              �?      @      @      @      4@       @       @      "@      9@      2@              @      @      �?      @      *@       @      "@                                      �?       @       @       @       @      2@      @              @                              *@      @      &@              �?      @      @       @      (@                      @      @      .@              �?      @      �?      @      @                               @              &@      @      �?                       @      (@                              �?       @              �?                               @              @       @      �?                              $@                              �?                       @                                              @      �?                               @       @                                       @             `l@     �L@     �j@      @@      E@      4@      M@     �m@     pp@     �J@     �J@      ]@     �q@     �p@      ,@      B@      @@     �X@      D@     @P@      .@      G@      @      "@      "@      *@      U@      X@      $@      ,@     �@@      R@     �S@      �?      ,@      (@      2@      &@      J@      &@     �D@      @      @      "@      "@     �@@     @Q@      $@      (@      ;@     �M@     �M@      �?      "@       @      2@      $@      @      �?                                              @      *@                              �?                                                     �G@      $@     �D@      @      @      "@      "@      =@      L@      $@      (@      ;@      M@     �M@      �?      "@       @      2@      $@      D@      "@      B@      @      @      "@      "@      ;@      G@      $@      @      ;@     �I@     �I@      �?      "@      @      0@      $@      5@              5@                      �?      @      1@      7@      @      @       @      <@      B@      �?      @      �?      (@      @      3@      "@      .@      @      @       @       @      $@      7@      @      @      3@      7@      .@              @      @      @      @      @      �?      @                                       @      $@              @              @       @                      @       @              @              @                                       @      $@                              @       @                                                      �?                                                                      @               @                              @       @              *@      @      @      �?       @              @     �I@      ;@               @      @      *@      3@              @      @              �?                      �?                                      7@      "@                      �?      @      @               @                                                                                      1@      @                      �?      �?      @                                                              �?                                      @      @                              @      @               @                              *@      @      @      �?       @              @      <@      2@               @      @       @      *@              @      @              �?       @                                                              @                                      @                      �?                      &@      @      @      �?       @              @      <@      (@               @      @       @      $@              @      @              �?       @               @      �?      �?                      @                                      @       @              �?                              @      @       @              �?              @      6@      (@               @      @      @       @               @      @              �?     @d@      E@     �d@      <@     �@@      &@     �F@     `c@     �d@     �E@     �C@     �T@     �j@     �g@      *@      6@      4@     @T@      =@     @Y@      ,@      R@      @      @              2@      `@      \@      (@      &@     �A@     ``@     �S@              $@      @     �C@      "@     �X@      ,@      R@      @      @              (@     @_@      \@      (@      &@     �A@     �_@     �Q@              $@      @      C@      @      Q@      (@     �I@      @      @              "@     �H@     �R@      $@      "@      8@     �T@     �O@               @      @      7@      @     �A@      @      <@                               @      C@     �I@      @      @      &@      E@      ?@              �?      �?      "@      @     �@@       @      7@      @      @              �?      &@      7@      @       @      *@      D@      @@              �?       @      ,@              ?@       @      5@      @      �?              @      S@      C@       @       @      &@     �F@      @               @      �?      .@      @      7@       @      @      @      �?              @      E@      1@               @      &@      9@       @              @      �?      &@      @       @              .@                                      A@      5@       @                      4@      @              �?              @      �?       @                                              @      @                                      @       @                              �?       @                                                      @      @                                              @                              �?       @       @                                              @                                              @      �?                                             �N@      <@     �W@      6@      <@      &@      ;@      ;@     �K@      ?@      <@      H@     �T@      \@      *@      (@      0@      E@      4@       @      �?      &@      @      @      �?                      @      @      �?              $@      1@      �?      �?      @      �?       @              �?      $@       @                                      �?      @      �?              @      @              �?      @              �?              �?      @                                              �?       @                      @       @                       @              �?                      @       @                                              �?      �?              @      �?              �?       @                       @              �?      �?      @      �?                      @      @                      @      ,@      �?                      �?      �?     �M@      ;@      U@      3@      9@      $@      ;@      ;@     �I@      8@      ;@      H@      R@     �W@      (@      &@      (@     �D@      2@      G@      3@     �I@      "@      6@      @      .@      6@     �@@      .@      0@     �A@     �M@      P@       @       @      @      >@      "@     �E@      2@     �F@      @      3@       @      *@      6@      @@      *@      ,@      7@     �M@      O@       @      @      @      ;@       @      @      �?      @      @      @      �?       @              �?       @       @      (@               @              �?       @      @      �?      *@       @     �@@      $@      @      @      (@      @      2@      "@      &@      *@      *@      ?@      $@      @      @      &@      "@      @      @      ?@      @       @      @      @       @      $@      @      &@      &@      @      3@      @       @      @      "@      @      @      @       @      @      �?               @      @       @      @               @      "@      (@      @      �?               @       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJS�&2hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKohnh4h7K ��h9��R�(KKo��hu�BH         4                   �2@����X��?�	           ��@                          �0@�&�<��?�           �@                            �?6������?�            `h@                           @���<,�?E             Y@                           �?�ݯ�f�?7             S@                           @�'�@݈�?             C@������������������������       �      �?             4@������������������������       ��8��8��?             2@	       
                    �?����U�?             C@������������������������       �J,�ѳ�?             1@������������������������       ����N8�?             5@������������������������       �VUUUUU�?             8@                           @���?=            �W@                           �?N��)x9�?             <@������������������������       �B{	�%��?             "@������������������������       �Dy�5��?             3@                           @@u8���?(            �P@                           �?�q�q�?             8@������������������������       ���(\���?             $@������������������������       �������?	             ,@                           �?Mtxj�-�?            �E@������������������������       �                     $@������������������������       �4 ��;��?            �@@       %                     @EjU�:0�?           �@                            @��Gx2b�?m           ��@                           @�U���`�?T           ��@                            �?`U(	:��?�            `u@������������������������       �Q��+Q�?k            �d@������������������������       ���L��?w            @f@                           @9��8���?r             h@������������������������       ��ZӼ��?             9@������������������������       �N�ư&�?d            �d@!       "                    @z3�Vf`�?            �D@������������������������       ��@�m�?             1@#       $                    @9��8���?             8@������������������������       ���(\���?             $@������������������������       ��X�C�?             ,@&       -                   �1@��8��?�             p@'       *                    �?f���.�?M            �]@(       )                    @�q�q�?             H@������������������������       ���(\���?             D@������������������������       �      �?              @+       ,                    @vzY���?.            �Q@������������������������       ��zv�X�?             F@������������������������       ��	j*D�?             :@.       1                    @�)񎴠�?\            �a@/       0                    �?w���??            �W@������������������������       �8��(y��?!            �I@������������������������       ���|���?             F@2       3                    �?f.i��n�?            �F@������������������������       ���8��8�?             8@������������������������       ����H��?             5@5       R                    �?hTT���?*           ��@6       C                    �?��7C��?�           ؎@7       <                    �?o����
�?           �y@8       ;                    �?�ܤ�?t             e@9       :                     �?��Kf��?h             c@������������������������       �䙢�c�?             G@������������������������       �1�Z�T�?K            �Z@������������������������       ���2Tv�?             .@=       @                    �?�%�J�?�            �n@>       ?                   �5@h�n��?0            @U@������������������������       �V>�� =�?             ?@������������������������       �Ix�5?�?              K@A       B                   �8@���(\?�?n             d@������������������������       �����	#�?H            �Y@������������������������       �N�e)���?&             M@D       K                   �;@��|���?q           ��@E       H                    @��^�?I           �@F       G                   �6@�UB���?�            �p@������������������������       ������H�?            �g@������������������������       ��Ԕ���?7            �T@I       J                   �8@>�s)�?�            �m@������������������������       �"��6%�?|            �h@������������������������       �Z�eY�e�?             E@L       O                   �=@�O��K��?(            @P@M       N                    �?�wC�Ҁ�?            �@@������������������������       ��T�6|��?             *@������������������������       ��Q����?
             4@P       Q                    �?     ��?             @@������������������������       �ףp=
�?             $@������������������������       �L�9���?             6@S       b                   �<@�C	�?�           ��@T       [                    �?L�{���?           ؙ@U       X                    @���tX�?�           8�@V       W                   �6@|X�/�?           �y@������������������������       �Q����?�            �m@������������������������       �K̠�?s            �e@Y       Z                    @?_��O�?�            �r@������������������������       �J���&0�?�            �p@������������������������       ����X�?             <@\       _                   �3@>|�����?J           x�@]       ^                    �?]����?X             b@������������������������       �O�ݥu�?!            �J@������������������������       �wj�s�?7             W@`       a                   �:@Eju��?�           ��@������������������������       �*b���?�           ��@������������������������       ��,x4T�?C            �[@c       j                    @jcèS@�?�            �n@d       g                    �?H��S�?]            �c@e       f                    @5��g�?            �A@������������������������       ��u]�u]�?	             5@������������������������       �s
^N���?
             ,@h       i                     @KfMP�?J            �^@������������������������       ���H!]�?+            @Q@������������������������       �&<���/�?            �J@k       n                    @�>��=��?<            �U@l       m                   �@@F>n���?6            �S@������������������������       � �$D4�?#            �G@������������������������       �]"?ӧ
�?             ?@������������������������       �|	�%���?             "@�t�bh�h4h7K ��h9��R�(KKoKK��h��B�A       �y@     �T@     �u@     �A@     @R@      ;@     �T@     ��@     ��@     @R@     @V@      e@     P�@     �{@      $@     @P@      O@     �_@      F@     @Z@      2@      P@       @       @              "@     �q@     �j@      "@       @      =@     �c@     �V@               @      @      7@      @      9@               @                                      S@     �G@                              ;@      &@                              �?              1@              @                                      <@      A@                              ,@       @                              �?              .@              @                                      9@      3@                              (@                                      �?              @              @                                      .@      $@                              @                                                      �?              @                                      @      @                              @                                                      @              �?                                      $@      @                                                                                      $@                                                      $@      "@                               @                                      �?               @                                                      @      @                               @                                                       @                                                      @       @                              @                                      �?               @                                                      @      .@                               @       @                                               @              @                                      H@      *@                              *@      "@                                              @               @                                      @      �?                              @       @                                              �?              �?                                      �?      �?                              @      �?                                              @              �?                                      @                                       @      @                                              @               @                                      E@      (@                              @      �?                                              �?                                                      3@      �?                               @      �?                                                                                                       @      �?                              �?                                                      �?                                                      &@                                      �?      �?                                               @               @                                      7@      &@                              @                                                                                                              $@                                                                                               @               @                                      *@      &@                              @                                                      T@      2@      L@       @       @              "@     �i@     �d@      "@       @      =@     @`@     �S@               @      @      6@      @     �G@      @      ;@                              "@     �e@     �_@      "@      @      ;@      R@      L@              @      @       @       @     �F@      @      7@                               @      c@     @_@      @      @      8@      R@     �J@              @      @      @      �?     �B@      @      ,@                              @      V@     �P@      @      @      3@      L@      @@              �?       @      @      �?      5@              @                               @      <@     �@@      @      @      "@      A@      1@              �?              @      �?      0@      @      @                              @      N@      A@      �?              $@      6@      .@                       @      �?               @       @      "@                              �?      P@      M@       @              @      0@      5@              @      �?      �?                                                                      2@       @                               @      @                                               @       @      "@                              �?      G@      L@       @              @      ,@      2@              @      �?      �?               @              @                              �?      4@       @       @      �?      @              @                               @      �?      �?              @                              �?      @      �?       @      �?                       @                                      �?      �?                                                      0@      �?                      @              �?                               @              �?                                                       @                                              �?                                                                                                       @      �?                      @                                               @             �@@      &@      =@       @       @                      A@      C@              @       @      M@      7@              @       @      ,@      @      6@               @               @                      2@      8@              �?       @      7@      "@              @       @      @              ,@              @                                      @      .@                              "@      �?                                              *@              �?                                      @      (@                              "@      �?                                              �?              @                                              @                                                                                       @              @               @                      ,@      "@              �?       @      ,@       @              @       @      @              @               @               @                      *@       @              �?      �?      @      @                                              @              �?                                      �?      �?                      �?      @      @              @       @      @              &@      &@      5@       @                              0@      ,@              @             �A@      ,@                              $@      @      @      "@      4@       @                              $@       @              �?             �@@      @                              @               @      "@      0@                                       @      @              �?              &@       @                              @               @              @       @                               @      @                              6@      �?                                              @       @      �?                                      @      @               @               @      &@                              @      @      @                                                               @                              �?      "@                              @       @       @       @      �?                                      @      @               @              �?       @                                      �?     s@      P@     �q@     �@@     �Q@      ;@     @R@     �q@     �w@      P@     @T@     `a@     �|@     0v@      $@     �L@     �L@      Z@     �C@     �\@      0@      P@      (@      =@      "@      (@     �W@     @e@      7@      9@     �A@      d@     `a@      @      *@      6@      ?@      ,@      N@       @      A@      @      4@      @      @      3@     �G@      (@      3@      (@     �K@     �M@      @      @      *@      5@      "@      ?@      �?      1@              @               @       @      >@       @      @      @      <@      0@               @       @      *@       @      ?@      �?      .@              @              �?      @      ;@      �?      @      @      ;@      $@               @       @      *@       @      *@              @                                              "@              �?      �?      $@       @                       @      @              2@      �?      &@              @              �?      @      2@      �?      @      @      1@       @               @              "@       @                       @                              �?      �?      @      �?                      �?      @                                              =@      @      1@      @      0@      @      @      &@      1@      $@      *@       @      ;@     �E@      @      @      &@       @      @      "@              @              @              @      @      "@      @      &@      �?      &@      .@               @      @       @      @       @                              �?              @      @      @              "@               @      @              �?      @                      @              @              @              �?              @      @       @      �?      "@      &@              �?      �?       @      @      4@      @      ,@      @      (@      @      �?       @       @      @       @      @      0@      <@      @       @      @      @      @      0@      @      @              "@      @               @      @      �?       @      @      (@      8@              �?      @       @              @      @      "@      @      @      �?      �?              @      @               @      @      @      @      �?       @      @      @     �K@       @      >@      @      "@      @      @      S@     �^@      &@      @      7@     @Z@      T@              @      "@      $@      @     �K@      @      =@      @       @      @      @     @R@     �]@      @      @      1@     @W@     �Q@              @      @      @      @      8@      @      2@      @      @      @      @      5@     �Q@      �?      �?      ,@     �I@     �F@              @              @       @      *@       @      @               @       @       @      2@      M@              �?      &@      ?@      B@                              @       @      &@      �?      &@      @       @      �?      �?      @      *@      �?              @      4@      "@              @                              ?@       @      &@       @      @              �?      J@      H@       @       @      @      E@      9@              @      @      @      @      >@       @      &@       @       @              �?      C@      D@                      @     �@@      9@              @              @      @      �?                               @                      ,@       @       @       @              "@                      �?      @                              @      �?      �?      �?       @      �?      @      @       @      @      @      (@      $@                      @      @                       @                                      �?      @      @      @      @      @      �?      @                      @      @                                                              �?      @      �?                      @      �?      @                                                       @                                                      @      @      @                                              @      @                      �?      �?      �?      �?       @                               @               @      &@      @                      @      �?                                              �?                                                              "@                                                              �?      �?      �?               @                               @               @       @      @                      @      �?             �g@      H@     `k@      5@      E@      2@     �N@     `g@     @j@     �D@      L@      Z@     �r@      k@      @      F@     �A@     @R@      9@     `f@     �F@     �e@      1@      :@      @      J@     �f@     �i@      <@     �G@      S@     �q@      h@              <@      ?@     �O@      2@     @S@      (@     �P@      @      *@       @      4@      [@     �X@      "@      2@      4@     ``@     �T@              (@      0@      2@      @      F@      @     �D@      �?       @       @      (@     �R@     �P@       @      &@      $@     �P@     �D@              "@      "@      "@      @      C@      �?      <@              @              @      N@     �A@      �?      @              B@      1@              @              @              @      @      *@      �?      @       @       @      .@      ?@      �?      @      $@      >@      8@              @      "@      @      @     �@@       @      9@       @      @               @     �@@      @@      @      @      $@     @P@     �D@              @      @      "@      @      @@       @      6@       @      @              @      ?@      >@      @      @      $@     �L@     �D@               @       @      "@      @      �?              @               @               @       @       @       @                       @                      �?      @                     �Y@     �@@     �Z@      ,@      *@      @      @@     @R@     �Z@      3@      =@      L@     �c@     �[@              0@      .@     �F@      (@      3@       @      $@      @      �?                      4@      @@       @       @      @      9@      $@                       @      &@      �?      @      �?      @      @                              �?      @       @       @      @      @      "@                       @      $@      �?      *@      �?      @              �?                      3@      <@                       @      3@      �?                              �?             �T@      ?@      X@      &@      (@      @      @@     �J@     �R@      1@      ;@     �I@     ``@     @Y@              0@      *@      A@      &@     �S@      8@      V@       @      $@      �?      :@     �I@      O@      (@      :@      F@     @^@     @T@              &@      @      >@      @      @      @       @      @       @      @      @       @      (@      @      �?      @      $@      4@              @      @      @      @      &@      @     �G@      @      0@      &@      "@      @      @      *@      "@      <@      ,@      7@      @      0@      @      $@      @      @      @      6@      @       @      @       @      @       @      $@       @      :@      "@      *@      @      *@      @      @       @              �?      "@              @               @      �?      �?      @              @      @                                       @                      �?      "@               @                      �?              @              @                                                                                              @               @              �?                       @      @                                       @              @       @      *@      @       @      @      @      @      �?      @       @      4@      @      *@      @      *@      @      �?       @      @       @      (@      �?       @      @              �?              @      @      .@      @       @       @      @      �?      �?      �?       @              �?      @              @      @       @      �?      @      @      @       @      @      @      "@       @              �?      @              9@               @      @      �?       @      @      @      �?       @      @      $@       @      @      �?      @      @      @              3@               @      @      �?       @      @      @      �?       @      @      "@       @      @      �?      @      @      @              @              @      @      �?       @      @              �?      �?      @      @              @      �?      @      @      �?              ,@              �?                              �?      @              �?              @       @                      @      �?                      @                                                                                      �?                              �?      �?�t�bub�,     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJI#hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmK}hnh4h7K ��h9��R�(KK}��hu�BX         >                   �4@FD���?�	           ��@       !                    �?P逩�@�?]           ��@                          �1@��G,8�?           ؊@                           @с�?�            `s@                           �?Jm_!'1�?}            �h@                            �?M��E"|�?Y            �a@������������������������       �\���(��?2             T@������������������������       ��r����?'             N@	       
                     �?^N��)x�?$             L@������������������������       �     ��?
             0@������������������������       �333333�?             D@                            �?p�� ��?@            �\@                           @��Y��O�?             ?@������������������������       ��s����?             5@������������������������       ����(\��?             $@                            �?���I��?.            �T@������������������������       ��������?             1@������������������������       ��袋.��?#            �P@                            �?�����?a           (�@                           @�Z����?�            @r@                           �?�q���?x             h@������������������������       �YL�Q��?Q            @_@������������������������       ����c��?'            �P@                           �?-����?C             Y@������������������������       �9��8���?             B@������������������������       �     ��?-             P@                          �3@,�� "�?�            p@                           �?7��G�?p            `f@������������������������       �~Ց�X��?&            �M@������������������������       �/�?�P��?J             ^@                            @��]���?6            �S@������������������������       ����*�?            �E@������������������������       �F�&�;K�?            �A@"       1                    @��Pr���??           P�@#       *                     @��wH��?�           p�@$       '                    @rl�f�(�?           �{@%       &                   �3@I��I��?w            @g@������������������������       ��*��=��?`            �b@������������������������       ��D�ϣ1�?             C@(       )                     �?    �C�?�             p@������������������������       �F�w>�
�?k            �d@������������������������       �^M<+	�?5            �V@+       .                    @��C�S�?�            �j@,       -                    @�S3��'�?q            �f@������������������������       ���ҥ��?e            `d@������������������������       ��P�n#�?             1@/       0                   �2@     @�?             @@������������������������       ���.���?             6@������������������������       �
ףp=
�?             $@2       7                    @�?�����?�            �o@3       4                   �0@��,j�?r            �f@������������������������       ��X�C�?
             ,@5       6                    @�t��*�?h             e@������������������������       �!���u��?M            �_@������������������������       �h�T�B�?            �D@8       ;                    �?��o!`��?1            �Q@9       :                     �?:/����?             <@������������������������       ��s�n_�?             *@������������������������       �
ףp=
�?             .@<       =                   �2@D�����?             E@������������������������       �/k��\�?             1@������������������������       �$������?             9@?       ^                    �?܈��(�?4           Ƞ@@       O                   �<@��=�_|�?q           �@A       H                   �7@�q��r�?�           8�@B       E                    �?:05V��?�             y@C       D                   �6@�{��7��?e            �d@������������������������       ��5��?E             Z@������������������������       ��8։'�?             �O@F       G                    �?��
�4�?�            `m@������������������������       �������?<            �Y@������������������������       ���HJ�}�?U            �`@I       L                    �?mpI�?�            Py@J       K                    �?���iO�?U            �a@������������������������       ����s��?!            �K@������������������������       ����lQ6�?4            @U@M       N                    �? xJ��4�?�            �p@������������������������       �Pdl<)�?1            �S@������������������������       ��k��ƕ�?x            `g@P       W                   �?@�	�1���?}            @k@Q       T                    @�p��[u�?I            @_@R       S                    �?p����?;            @Y@������������������������       �t��:��?             C@������������������������       �W�7�L�?$            �O@U       V                   �=@�q�q�?             8@������������������������       �     ��?             0@������������������������       �      �?              @X       [                     @�s����?4            @W@Y       Z                    �?\�\��?            �I@������������������������       �ƵHPS!�?             *@������������������������       �g�˹�?             C@\       ]                    �?�^�:�?             E@������������������������       ��.�?�P�?             .@������������������������       ��T'"7�?             ;@_       n                    �?Ш�さ�?�           ��@`       g                     �?�pi���?�            @s@a       d                     �?�����?s            @f@b       c                   �7@a���i��?8             V@������������������������       �8^s]e�?!             M@������������������������       ���O��O�?             >@e       f                   �5@����<�?;            �V@������������������������       �n�1�^�?             A@������������������������       �����>4�?)             L@h       k                    �?��oOa��?[            @`@i       j                     @�`�`�?+             N@������������������������       �G ��h�?            �E@������������������������       �P�|�@�?             1@l       m                   �<@�������?0            �Q@������������������������       �-�����?$             I@������������������������       ��G�z��?             4@o       v                   �<@Z{L��?�           x�@p       s                   �;@s�K�i^�?�           �@q       r                    @O;�O�?�           Є@������������������������       �R)�Ǝ&�?h           ��@������������������������       ��ƺ�W�?3            @R@t       u                     �?��Q��?             D@������������������������       ��K~���?             .@������������������������       �������?             9@w       z                   �?@F4�����?C            @[@x       y                    @�U�����?)            �P@������������������������       �Ό��i�?            �G@������������������������       �ffffff�?             4@{       |                    @�^�:�?             E@������������������������       ������?             7@������������������������       ����Դ�?             3@�t�bh�h4h7K ��h9��R�(KK}KK��h��B8J       0}@     �S@     �r@     �E@      T@      =@     �T@     �@     ��@      P@     @R@      d@     ��@     �{@       @     �N@     �J@      `@     �P@     �n@      1@     @\@      @      ,@      �?      2@     0z@     ps@      @      8@     �J@     �q@     �e@              3@      @     �G@      &@     �^@      @      C@      �?      @      �?      $@      p@     �d@              "@      4@     �`@     �P@              @              3@       @     �J@      @      ,@                              @      _@     �M@                      �?     �D@      &@                              �?              <@      @       @                              �?     @V@      <@                      �?      ?@      @                                              3@      @       @                                     @Q@      4@                      �?      ,@      @                                              "@              @                                     �H@      $@                      �?      @       @                                              $@      @      @                                      4@      $@                              "@      @                                              "@                                              �?      4@       @                              1@      �?                                              �?                                                      @       @                              $@                                                       @                                              �?      1@      @                              @      �?                                              9@              @                               @     �A@      ?@                              $@      @                              �?              @                                               @      "@      0@                                                                      �?               @                                               @      @      (@                                                                      �?              �?                                                      @      @                                                                                      6@              @                                      :@      .@                              $@      @                                               @               @                                      @       @                               @                                                      ,@              @                                      7@      *@                               @      @                                             �Q@       @      8@      �?      @      �?      @     �`@     �Z@              "@      3@     �V@      L@              @              2@       @      E@              (@      �?      �?               @      O@     �Q@              @      "@     �L@      5@               @              @              2@              @      �?                       @      D@     �L@              @      @      D@      0@               @              @              *@              @                                      4@     �B@               @      @      =@      ,@                              @              @              �?      �?                       @      4@      4@               @              &@       @               @              �?              8@               @              �?                      6@      ,@              @      @      1@      @                              �?              $@               @              �?                      (@      �?               @      @      @                                                      ,@              @                                      $@      *@              �?       @      (@      @                              �?              <@       @      (@               @      �?      @      R@     �A@               @      $@      A@     �A@              @              *@       @      5@      �?      "@                              @      J@      <@              �?       @      4@      1@              @              &@       @       @      �?      @                                      "@      &@                       @      @       @              @               @              *@              @                              @     �E@      1@              �?      @      1@      "@                              @       @      @      �?      @               @      �?              4@      @              �?       @      ,@      2@                               @              @              @               @      �?              .@      @              �?      �?      @      @                              �?              @      �?                                              @      �?                      �?      "@      *@                              �?             �^@      (@     �R@      @      &@               @      d@     @b@      @      .@     �@@     �b@     �Z@              *@      @      <@      "@     �W@      (@     �G@      @      "@              @     @`@      W@      @      .@      2@      ]@     @T@               @       @       @       @     �P@      @      7@              @              @     @Z@     @Q@      @      "@      &@     �R@      K@              @              @      @      9@       @      1@              �?              @      <@      A@      @      @       @      >@      ;@              @               @      @      9@       @      &@              �?              @      3@      ?@      @      @       @      6@      3@              @                       @                      @                                      "@      @                               @       @                               @       @     �D@       @      @              @              �?     @S@     �A@      �?      @      "@     �F@      ;@               @              �?       @      :@       @      @              @              �?      E@      2@              @      "@      =@      7@               @              �?       @      .@               @                                     �A@      1@      �?                      0@      @                                              <@       @      8@      @      @              @      9@      7@              @      @     �D@      ;@              @       @      @       @      :@      @      5@      @      @              @      3@      6@              @      @      B@      6@              �?      �?      @      �?      9@      @      4@      @      @               @      (@      5@              @      @     �A@      2@                      �?      @      �?      �?              �?                              �?      @      �?                              �?      @              �?                               @       @      @                                      @      �?                      @      @      @               @      �?      �?      �?       @      �?                                              @      �?                      @       @       @               @      �?      �?      �?              �?      @                                                                              @      @                                              <@              <@       @       @              �?      ?@      K@                      .@     �A@      9@              @      @      4@      �?      $@              5@       @       @                      6@      C@                      *@      :@      4@              @      @      1@      �?                                       @                      @      @                                                                                      $@              5@       @                              1@      ?@                      *@      :@      4@              @      @      1@      �?       @              3@       @                              @      8@                      "@      3@      0@               @      @      0@      �?       @               @                                      $@      @                      @      @      @              @      �?      �?              2@              @                              �?      "@      0@                       @      "@      @                              @              &@              @                                      �?       @                       @      �?      @                              @              @              @                                      �?                               @               @                              �?              @               @                                               @                              �?      �?                               @              @               @                              �?       @      ,@                               @       @                                              �?              �?                              �?      @      @                               @      �?                                              @              �?                                       @      "@                              @      �?                                             �k@     �N@     �g@     �B@     �P@      <@     @P@      d@     �q@      N@     �H@     �Z@     �s@     q@       @      E@      G@     �T@      L@     �Z@      ;@     �X@      9@      F@      6@      A@     �A@     �W@      <@     �@@     @Q@     �_@     @a@      @      9@     �A@     �C@      E@      W@      7@     @S@      0@      4@      *@      9@     �A@      S@      6@      4@     �J@     �^@     �^@      �?      1@      5@      9@      :@     �I@       @     �D@       @      @      @      @      8@     �H@      *@      (@      5@      O@     �K@              $@       @      .@      @      <@              *@       @      @      �?       @      .@      2@       @       @      @     �B@      6@              @      @      @      �?       @              "@       @       @      �?       @      $@      &@                       @      >@      3@              @      �?      �?      �?      4@              @              �?                      @      @       @       @      @      @      @              �?      @      @              7@       @      <@      @      @      @      @      "@      ?@      &@      $@      ,@      9@     �@@              @      @      &@      @      0@      �?      .@      @      �?              @      @      6@       @       @      @      *@      &@              �?      �?      @              @      @      *@      @      @      @       @      @      "@      "@       @       @      (@      6@              @      @       @      @     �D@      .@      B@       @      *@      @      2@      &@      ;@      "@       @      @@      N@      Q@      �?      @      *@      $@      5@      8@       @      $@              @       @       @      @      "@      �?      @       @      <@      4@              �?      �?      @      &@      @      @      @                      �?       @      �?      @              @      @      (@      @                      �?      @      @      5@       @      @              @      �?              @      @      �?              @      0@      0@              �?               @      @      1@      @      :@       @      $@      @      0@      @      2@       @      @      8@      @@      H@      �?      @      (@      @      $@      $@      �?      $@      @       @              �?               @      �?              @      ,@      5@              �?              @       @      @      @      0@      @       @      @      .@      @      0@      @      @      1@      2@      ;@      �?      @      (@       @       @      ,@      @      5@      "@      8@      "@      "@              2@      @      *@      0@      @      .@      @       @      ,@      ,@      0@      (@      @      0@       @      "@      @      @              1@      @      @      @      @      @              @      @      (@      "@      &@      @      ,@       @      @      @      @              1@      @      @      @       @       @              @      @      &@      @      "@      @      @               @              �?              @       @       @       @               @               @              @      @       @      �?      $@       @      �?      @      @              ,@      @      �?       @       @                      �?      @       @      @      �?               @              @                                              �?               @      @              �?      @      �?      @      �?               @              @                                                               @      @                                      @                                      �?                                              �?                      �?              �?      @      �?               @              @      @      .@      @       @              �?      �?      "@      (@              "@      @      @       @       @      @       @              @      @      @      �?                      �?      �?      @      (@              @              �?      @       @               @              @               @                                               @                      @                      �?                                      �?      @      @      �?                      �?      �?      @      (@              �?              �?      @       @                              �?       @       @      @       @                              @                      @      @      @       @              @                                      @               @                                                      @      �?       @       @                                      �?       @      @      @                                      @                       @      @      �?                      @      ]@      A@     �V@      (@      6@      @      ?@     @_@     �g@      @@      0@      C@     `g@     �`@      @      1@      &@     �E@      ,@      =@      1@      6@      @      @      @      @      ?@     @R@      (@      @      "@      B@     �F@               @       @      "@              (@      �?      1@              �?      �?      @      7@     �I@      $@       @      @      6@      <@              �?               @              @              @                      �?      @      @      2@       @       @      @      *@      2@              �?               @              @              @                      �?       @      @      *@               @       @      $@      &@                               @              @                                              �?      �?      @       @              �?      @      @              �?                              @      �?      &@              �?                      1@     �@@       @              �?      "@      $@                                              �?      �?      @                                      @      2@                              @       @                                              @              @              �?                      ,@      .@       @              �?      @       @                                              1@      0@      @      @       @       @      @       @      6@       @      @      @      ,@      1@              �?       @      @              (@      @      @                               @      @      *@               @      �?      $@      @              �?                              $@      @      @                               @      @      (@               @              @                      �?                               @      �?                                                      �?                      �?      @      @                                              @      (@       @      @       @       @      �?       @      "@       @       @      @      @      &@                       @      @              @      &@       @               @              �?       @      @       @               @      @      $@                      �?       @                      �?              @               @                       @               @       @      �?      �?                      �?      @             �U@      1@     @Q@      "@      3@      @      9@     �W@     @]@      4@      $@      =@     �b@     �V@      @      .@      "@      A@      ,@     �S@      0@     �L@      "@       @      �?      8@     �V@     @\@      &@      $@      4@     �`@     @R@      �?      &@      "@      9@      ,@      S@      *@     �L@       @       @      �?      8@     @V@      [@      "@      $@      3@     �^@      R@      �?      &@      @      8@      "@     �P@      &@     �H@      @      @      �?      1@      S@     �Z@       @       @      1@     �[@      Q@              $@      @      7@      "@      $@       @       @      @      @              @      *@      �?      �?       @       @      *@      @      �?      �?              �?               @      @              �?                               @      @       @              �?      (@      �?                      @      �?      @               @                                                                              �?      �?      �?                      @              @       @      �?              �?                               @      @       @                      &@                                      �?              "@      �?      (@              &@       @      �?      @      @      "@              "@      0@      1@       @      @              "@              @              @              &@                      @              @              @      ,@      (@      �?       @               @              @              �?              &@                      �?              @               @      "@      "@      �?      �?              @              �?               @                                       @                              �?      @      @              �?              @              @      �?      "@                       @      �?              @      @              @       @      @      �?       @              �?              �?      �?      @                       @                              @              @       @       @      �?       @                               @              @                              �?              @       @                              @                              �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��xyhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKyhnh4h7K ��h9��R�(KKy��hu�Bx         :                   �2@�Qb�g{�?�	           ��@                           @�#,��?�           ��@                           �?���7�??            �@                          �1@��7F�?�             v@                            �?
�GILH�?y            `i@                           �?�X� �(�?:            �X@������������������������       �B�0�~��?             F@������������������������       �2��ޥ�?"            �K@	       
                    @M�h���??             Z@������������������������       �L�r*��?4            @U@������������������������       ����,�?             3@                           �?���.��?d            �b@                            @F���\��?+            �O@������������������������       �6YE�?            �@@������������������������       �t�@�t�?             >@                           @���y��?9            �U@������������������������       �     �?*             P@������������������������       ������?             6@                            @�6��,�?b            �d@                           @=�>���?G            �]@                           �?36����?9            �X@������������������������       �c��gS~�?"             M@������������������������       ��b����?            �D@                            �?�(\����?             4@������������������������       ���(\���?             $@������������������������       �{�G�z�?             $@                           @��Sڙ��?            �F@������������������������       ���x��?             7@������������������������       ��ˠT�?             6@       -                     @:�_ra�?h           �@       &                    @�c�����?           P{@        #                   �1@��&��?�            Pt@!       "                    @��>��G�?�            �j@������������������������       ����RP��?�            `i@������������������������       ��q�q�?	             (@$       %                     �?��D!Z�?M            �[@������������������������       ���0�*�?             9@������������������������       ��������?<            @U@'       *                    �?����>4�?E             \@(       )                    �?�&1��?             I@������������������������       ��(ݾ�z�?             :@������������������������       ���8��8�?             8@+       ,                     �?�� =�	�?&             O@������������������������       ��]K�=�?             I@������������������������       �9��8���?             (@.       5                   �1@��}��?I             [@/       2                    @��9Z�?+            �M@0       1                    @T����?             C@������������������������       �<5rԹ��?             7@������������������������       ��h$���?	             .@3       4                    �?4և����?             5@������������������������       �9��8���?	             (@������������������������       �X�<ݚ�?             "@6       7                    �?�R�����?            �H@������������������������       �Cu��?             5@8       9                    @c}h���?             <@������������������������       �*�c{��?             3@������������������������       �0�����?             "@;       Z                    �?��ړ��?�           H�@<       K                    �?�	���3�?3           0�@=       D                    �?�3��0��?            z@>       A                     �?�#t�K��?Y            �`@?       @                    �?w�M��:�?             ;@������������������������       ��1G����?
             *@������������������������       ��Cc}�?
             ,@B       C                    �?�GLS^��?E            �Z@������������������������       �	j*D>�?#             J@������������������������       ��,騷}�?"             K@E       H                   �<@E�(��?�            �q@F       G                    �?^M<+��?�             n@������������������������       ����Y��?9            �S@������������������������       �v@A�W�?f             d@I       J                    �?�o1�?            �F@������������������������       ��o^M<+�?
             .@������������������������       �>
ףp=�?             >@L       S                    �?��x�G�?           P�@M       P                   �=@    �l�?�             p@N       O                   �;@�r���V�?�            `m@������������������������       ��9�mR�?�            �j@������������������������       �q=
ףp�?             4@Q       R                   �>@lv�"��?             5@������������������������       �VUUUUU�?             "@������������������������       �UUUUUU�?             (@T       W                    �?O�Ï�a�?|           P�@U       V                    @ ������?�            �o@������������������������       �[$��m�?             J@������������������������       ����O���?{            @i@X       Y                     �?�:�z!M�?�            �v@������������������������       �ss���?K            �`@������������������������       �w�T�|�?�            �l@[       j                    �?OQ{H�?�           `�@\       c                    @�v�|S��?.           @]       `                   �9@ ?R�N��?�            �q@^       _                    �?%�4�X��?�            �l@������������������������       � �C5�?M            �\@������������������������       ���ʅ���?A            �\@a       b                   �;@P�����?            �M@������������������������       ��zv��?
             6@������������������������       ��,b+���?            �B@d       g                    �?��D�x�?�            @j@e       f                    @�d��?:            �X@������������������������       ��̿0�=�?             ?@������������������������       �y�rك8�?#            �P@h       i                    ;@Y�Cc�?I             \@������������������������       ��P�)�?B            @Y@������������������������       ��ˠT�?             &@k       r                   �:@`.�e`�?�           ��@l       o                   �7@��g9*�?4           �@m       n                    �?�&GI���?�           `�@������������������������       �ڪ�&�?�            Ps@������������������������       �a��'9�?�            pw@p       q                    �?�l�37�?�             j@������������������������       � �~s��?;            @W@������������������������       ��f>���?J             ]@s       v                     @f�b�_��?h            @e@t       u                    @�V����?R            �`@������������������������       �H�4����?4            �T@������������������������       ��\m����?             I@w       x                    @]��N��?             C@������������������������       ��5;j��?             5@������������������������       �J,�ѳ�?
             1@�t�bh�h4h7K ��h9��R�(KKyKK��h��B�G       �{@     �Q@     �u@      =@     �N@      7@      U@     ��@     ��@     @P@     �W@     �a@      �@     }@      .@     �O@     �G@      _@      H@     �`@      *@     @T@      �?      @              $@     r@      j@      @      $@      1@     �f@     @S@              @       @      3@      @     �T@      @      H@      �?      @               @     �W@     �Y@      @       @      "@     �W@      E@              @      �?      (@      @     �O@      @     �@@      �?      @              �?      Q@     �I@      �?      @       @      R@      8@              @      �?      &@      @     �F@              .@              @                      J@      6@      �?       @      @      E@      &@              �?      �?       @       @      3@              @              �?                     �A@      (@      �?       @      �?      2@       @                              �?       @      &@              @                                      *@      "@                              @      �?                                               @               @              �?                      6@      @      �?       @      �?      &@      �?                              �?       @      :@              $@               @                      1@      $@                      @      8@      "@              �?      �?      �?              6@              @               @                      1@       @                      @      6@      @              �?      �?                      @              @                                               @                               @      @                              �?              2@      @      2@      �?                      �?      0@      =@               @      @      >@      *@              @              "@      �?      "@       @       @                                      *@      @              �?      �?      1@      @              @              @              @               @                                      $@      @              �?      �?       @      �?                                               @       @                                              @       @                              "@      @              @              @              "@       @      0@      �?                      �?      @      8@              �?      @      *@      "@                              @      �?      @       @      $@      �?                      �?      �?      6@              �?      @      "@      @                              @              @              @                                       @       @                              @       @                                      �?      3@      �?      .@                              �?      ;@      J@       @      @      �?      7@      2@                              �?              0@              *@                              �?      7@      D@      �?      @      �?       @      &@                              �?              .@              (@                              �?      3@      ;@      �?      @      �?      @      &@                              �?              @              @                                      *@      4@              @      �?      @      @                              �?               @               @                              �?      @      @      �?                      @      @                                              �?              �?                                      @      *@                              �?                                                                                                              �?       @                              �?                                                      �?              �?                                      @      @                                                                                      @      �?       @                                      @      (@      �?                      .@      @                                              @               @                                      �?      @                              $@      @                                                      �?                                              @       @      �?                      @      @                                             �I@       @     �@@                               @     @h@     �Z@       @       @       @     �U@     �A@               @      �?      @       @     �C@       @      &@                              @     �d@      W@       @      �?      @     �P@      ?@               @      �?      @              5@      @      "@                              @      a@     @Q@      �?      �?      @     �K@      6@                              �?              0@      @      @                               @     @V@      M@              �?       @      ?@      @                              �?              ,@      @      @                               @     @U@      M@              �?       @      =@      @                              �?               @                                                      @                                       @      @                                              @              @                              �?      H@      &@      �?              �?      8@      .@                                              @                                                       @      @                      �?      @      "@                                               @              @                              �?      G@       @      �?                      1@      @                                              2@      @       @                              @      ;@      7@      �?              @      &@      "@               @      �?      @              @               @                              @      1@       @                       @      @      @              �?              �?              @              �?                                      &@      @                       @              @                                              @              �?                              @      @       @                              @      @              �?              �?              (@      @                                              $@      .@      �?              �?       @      @              �?      �?      @              @      @                                              $@      (@      �?              �?      @      @              �?      �?      @              @                                                              @                              @                                                      (@              6@                              �?      >@      ,@              �?       @      4@      @                                       @       @              @                                      4@      "@              �?      �?      (@      @                                               @              @                                      0@      @              �?              @      @                                               @              �?                                      &@      @              �?              �?       @                                                               @                                      @      �?                              @       @                                              @              �?                                      @      @                      �?      @                                                      @              �?                                       @      @                                                                                                                                               @                              �?      @                                                      @              2@                              �?      $@      @                      �?       @                                               @      �?              "@                                       @       @                              �?                                                      @              "@                              �?       @      @                      �?      @                                               @       @              "@                                              �?                              @                                                      �?                                              �?       @       @                      �?                                                       @     ps@     �L@     pp@      <@      M@      7@     �R@     �p@     �y@      N@      U@      _@     �z@     @x@      .@     �L@     �F@     @Z@     �E@      a@      :@     @b@      .@      C@      1@      B@      Q@      a@      ;@      J@     �P@     @e@     `g@      &@     �@@      @@      N@      A@      A@      @     �A@      �?      .@      �?      &@      :@     �L@       @      7@      3@     �S@     �M@              "@      "@      2@      $@      $@       @      @               @              @       @      ?@      �?      &@       @      6@      7@              @      @       @      @      @               @              �?              �?              &@              �?              @                               @                       @                                                              @                              @                              �?                      �?               @              �?              �?              @              �?              �?                              �?                      @       @      @              �?               @       @      4@      �?      $@       @      0@      7@              @      @       @      @      @       @      @                                      @      ,@      �?      @      �?      $@      @                               @      �?      @                              �?               @      @      @              @      �?      @      3@              @      @               @      8@      @      >@      �?      *@      �?       @      2@      :@      @      (@      1@      L@      B@              @      @      0@      @      7@      @      5@      �?      $@      �?      @      1@      8@      @      $@       @     �J@      ?@              @      @      0@      @      @       @      @              �?      �?       @      *@      &@       @      @       @      3@      @              �?      �?      �?       @      3@      �?      .@      �?      "@               @      @      *@      @      @      @      A@      9@              @       @      .@      @      �?              "@              @              @      �?       @       @       @      "@      @      @              �?      �?               @                      �?                                      �?       @       @              �?       @      @                                      �?      �?               @              @              @                               @       @      �?                      �?      �?              �?     �Y@      5@     �[@      ,@      7@      0@      9@      E@     �S@      3@      =@      H@      W@      `@      &@      8@      7@      E@      8@     �J@       @      8@      �?      $@              @      1@      ?@       @       @      $@      =@     �A@      @      @      @      1@       @      G@       @      7@      �?      @              @      1@      >@      @       @      $@      =@     �A@      @      @      @      ,@       @      E@       @      7@      �?      @              @      1@      :@      @       @      $@      =@      =@      @      @      @      ,@              @                              @              �?              @                                      @                                       @      @              �?              @                              �?      @                                              �?      �?      @              @                                                                      �?                                              �?              @              @              �?              @                              �?      @                                                      �?                      I@      3@     �U@      *@      *@      0@      5@      9@      H@      &@      ;@      C@     �O@     @W@       @      4@      3@      9@      6@     �A@      @      @@      @      @      @      ,@      ,@      >@              @      "@      @@      @@              @      (@      @      $@      @              &@                              �?      @      @              �?       @      @      @              @       @       @      @      =@      @      5@      @      @      @      *@      "@      8@              @      @      =@      <@              �?      $@      @      @      .@      .@     �K@      "@      "@      &@      @      &@      2@      &@      5@      =@      ?@     �N@       @      0@      @      2@      (@      @      @      8@      @      @      @       @      @      @       @      $@      @      (@      ;@              &@       @      @       @      $@       @      ?@      @      @      @      @       @      &@      "@      &@      7@      3@      A@       @      @      @      .@      $@     �e@      ?@     @]@      *@      4@      @      C@     `i@     pq@     �@@      @@     �L@     Pp@      i@      @      8@      *@     �F@      "@      G@      *@      ?@      @      @      @      &@     �K@     �\@      "@       @      6@     �R@     �S@              (@      �?      @      @      6@      @      3@       @      �?      @      @      6@     @P@      @       @      3@     �I@     �E@              "@              @      �?      5@      @      *@              �?       @      @      4@     @P@              �?      *@     �E@      A@               @              �?      �?      "@      @      @              �?      �?              @     �@@              �?       @      =@      .@                              �?              (@              "@                      �?      @      ,@      @@                      @      ,@      3@               @                      �?      �?              @       @              �?      �?       @              @      @      @       @      "@              @               @              �?               @                                      �?              @               @               @              @                                              @       @              �?      �?      �?              @      @      @       @      �?               @               @              8@      @      (@      �?      @              @     �@@      I@       @              @      8@     �A@              @      �?       @      @      $@      @      @                                      0@     �@@                       @      ,@      .@                                              @              �?                                      "@      "@                       @       @      @                                              @      @      @                                      @      8@                              (@      &@                                              ,@      @      @      �?      @              @      1@      1@       @              �?      $@      4@              @      �?       @      @      ,@      �?      @      �?      @              @      1@      0@       @              �?      "@      1@              @      �?       @      �?              @                                                      �?                              �?      @                                      @      `@      2@     �U@      $@      .@      @      ;@     �b@     �d@      8@      8@     �A@     @g@     �^@      @      (@      (@      D@      @     @Z@      *@      R@      "@      @              3@     �a@     �c@      *@      5@      <@     `d@     �V@      @      "@      @      @@      @     �V@      (@      J@      @      @              *@      ^@      _@      (@      ,@      7@      ^@     �M@              @      @      5@       @      B@      @      0@      �?                      @     @P@     �Q@      @       @       @      J@      ;@              �?      @      .@              K@      "@      B@      @      @              "@     �K@      K@      @      @      5@      Q@      @@              @       @      @       @      .@      �?      4@      @      �?              @      6@     �@@      �?      @      @     �E@      @@      @      @              &@      �?      @      �?      @       @                      �?      ,@      .@      �?      @      @      1@      3@              @              @      �?      $@              0@       @      �?              @       @      2@              @       @      :@      *@      @                      @              7@      @      ,@      �?       @      @       @      @      @      &@      @      @      7@      @@              @      @       @      �?      7@      @      &@      �?      @      �?      @      @      @      "@      @      @      ,@      7@               @      @       @      �?      $@      @      @              @      �?      �?      @      @       @               @      "@      1@               @      @      @              *@      �?       @      �?                       @       @              �?      @       @      @      @                      @      �?      �?              �?      @              �?       @      @               @       @              @      "@      "@              �?                                               @              �?              @               @       @              �?              "@                                                      �?      �?                       @      �?                                       @      "@                      �?                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�EcmhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKuhnh4h7K ��h9��R�(KKu��hu�B�         8                    �?�/�s��?�	           ��@                           �?"o��P�?            p�@                           �?���q��?h           @�@                          �6@��K���?�            `p@                            �?;�lO�?a             c@                          �1@h�����?              L@������������������������       �������?             .@������������������������       ����.}*�?            �D@	       
                     �?9��8�c�?A             X@������������������������       ���ӭ�a�?             B@������������������������       ���Wϊ�?&             N@                          �7@=�@�Nk�?D            �[@������������������������       �h���I�?             7@                           @X#��^�?8            �U@������������������������       ��g���j�?(            @P@������������������������       ��7�A�?             6@                          �1@��*1��?�             r@������������������������       ��m۶m��?             <@                          �<@�ɒ���?�            `p@                           �?�����?�             m@������������������������       ����O_[�?,            @P@������������������������       �¡�ZJ�?s            �d@                          �?@hE#߼�?             >@������������������������       �窷uJ��?             3@������������������������       �*L�9��?             &@       )                    @*b�z9�?�           А@       "                   �<@�<�]a �?�           0�@                           �?d]!��?e           ��@                            @[C:�{H�?�            @k@������������������������       ��:�
�7�?F            �]@������������������������       �k+��ݓ�?E             Y@        !                    @B������?�            �u@������������������������       ���O~��?�            �o@������������������������       �9�M���?>            �W@#       &                   �=@��v��?1            �S@$       %                    �?�!pc��?             6@������������������������       �      �?              @������������������������       ��m۶m��?             ,@'       (                     �?�X�C�?"             L@������������������������       ��� Ce��?             >@������������������������       ���c����?             :@*       1                   �3@HĮ��:�?           �z@+       .                    @(vb'vb�?;             Z@,       -                     �?���З�?            �C@������������������������       �     ��?             0@������������������������       �`������?             7@/       0                    @�K���?$            @P@������������������������       �W��_��?            �K@������������������������       ��(\����?             $@2       5                     �?[��g!�?�            `t@3       4                   �:@�0���.�?=            @Z@������������������������       �[�6z���?%            @P@������������������������       ��p=
ף�?             D@6       7                    �?����W�?�            �k@������������������������       �N����?8            �T@������������������������       �h��O�?R            @a@9       V                    �?�:Xʺ��?�           ڡ@:       I                    @*���?�           <�@;       B                    @~v@����?�           ��@<       ?                    @�p��b��?'            }@=       >                     @ )O7�?�             r@������������������������       �d�*����?�            �j@������������������������       ���
���?1            �R@@       A                   �7@g�aA�;�?v            @f@������������������������       ��N(i�?`            @b@������������������������       �     `�?             @@C       F                     �?��b���?d            �c@D       E                    @n�'�*��?4            �T@������������������������       ���*�?-            �Q@������������������������       �b���i��?             &@G       H                   �2@A�F<��?0             S@������������������������       �jW�v%j�?            �D@������������������������       �5��g�?            �A@J       O                    @�q{��?'           �}@K       L                    �?`�����?            �D@������������������������       �؇���X�?             ,@M       N                    @ن��s��?             ;@������������������������       ��h$���?
             .@������������������������       ��q�q�?             (@P       S                   �1@/G(�S>�?           `{@Q       R                   �0@�V�����?1            @R@������������������������       �θ	j*�?             :@������������������������       ������w�?             �G@T       U                   �8@�:r:���?�            �v@������������������������       ���\o�1�?�            0r@������������������������       �3�B��?/            �R@W       f                   �5@w}�����?�           x�@X       _                   �1@6�D]��?�           ��@Y       \                     @��kv��?             j@Z       [                   �0@�ՙ�?g             e@������������������������       ��k|���?"            �O@������������������������       ����D��?E            @Z@]       ^                    @��RQJ�?            �D@������������������������       �������?             .@������������������������       �5��?�?             :@`       c                     @�i� �?<           8�@a       b                   �2@�%ˏ��?�            �y@������������������������       �y�*3��?.            �S@������������������������       ����
֊�?�            �t@d       e                   �2@`��((�?F            �Z@������������������������       ��m(�9W�?            �E@������������������������       �     ��?,             P@g       n                   �9@�u�?�?1           `|@h       k                     �?���;�?�             q@i       j                    @�p=
�c�?3             T@������������������������       �Ę}�V`�?            �A@������������������������       �ڤ�:�^�?            �F@l       m                    @jJ�$���?�            @h@������������������������       �Weׇ�n�?Z            �`@������������������������       �S��d�?)             N@o       r                   �;@��*̉�?{            �f@p       q                    @��xJ���?.            @Q@������������������������       �fP*L��?             6@������������������������       �Y�� ��?             �G@s       t                    @�>�6�?M            �[@������������������������       ������*�?"             H@������������������������       �l|��Y�?+            �O@�t�bh�h4h7K ��h9��R�(KKuKK��h��BxE       p~@     �R@     `t@      C@     �V@      7@     �Y@     p�@     �@      H@      U@     `e@     �@     �y@      ,@     @S@      G@      `@     �H@     �k@     �A@      e@      ,@     �K@      1@      I@     �_@     �h@      6@      I@     �V@     `h@      i@      @     �F@      ;@      R@     �A@     �T@       @      E@      �?      2@      �?      (@      N@     @U@      "@      ,@      ?@     �Q@     �O@              *@      @      3@      0@      B@      @      5@              @      �?      @      B@      L@      @       @      "@      B@      8@              @      �?      @       @      6@              *@               @               @      A@     �@@              @      @      6@      $@                              @              (@              @                                      @      *@                      @      $@      @                                              @              @                                      @      �?                              �?       @                                              "@              �?                                              (@                      @      "@      @                                              $@              "@               @               @      =@      4@              @      �?      (@      @                              @              @               @               @               @      &@      $@              �?              @                                                      @              @                                      2@      $@              @      �?      "@      @                              @              ,@      @       @              �?      �?      �?       @      7@      @      @       @      ,@      ,@              @      �?       @       @       @               @                                               @      @      �?       @              @                                              @      @      @              �?      �?      �?       @      5@       @      @              ,@      "@              @      �?       @       @      @      @      @              �?      �?              �?      4@       @      @              @      @              @      �?      �?      @       @       @                                      �?      �?      �?                              "@       @              �?              �?       @      G@       @      5@      �?      .@              "@      8@      =@      @      @      6@     �A@     �C@              "@      @      ,@       @       @                                                      &@      @                      �?      "@      �?                                              F@       @      5@      �?      .@              "@      *@      9@      @      @      5@      :@      C@              "@      @      ,@       @      F@       @      4@      �?       @               @      *@      9@      @      @      1@      9@     �B@               @      @      "@       @      "@              �?              @              �?       @      @       @      �?      @      @      ,@              @      @      �?      �?     �A@       @      3@      �?      @              �?      @      3@       @      @      &@      5@      7@              @       @       @      @                      �?              @              @                               @      @      �?      �?              �?      �?      @                              �?              @              @                                      �?      �?      �?                      �?      @                                              @                                               @      @                              �?              �?             `a@      ;@     �_@      *@     �B@      0@      C@     �P@     @\@      *@      B@     �M@      _@     @a@      @      @@      4@     �J@      3@     @Z@      2@     �N@       @      9@       @      2@     �D@     @P@      $@      0@      <@     �P@     @X@      @      5@      *@     �B@      @     �X@      1@     �J@      @      8@       @      $@     �D@      O@      "@      *@      3@     @P@      W@      @      $@      &@      :@      @     �E@      @      (@              @       @      @      ;@      5@              @      @      >@      A@       @       @      @       @      �?      5@      �?      $@               @               @      6@      @              @      @      .@      .@              @      @      @              6@      @       @              �?       @       @      @      .@              �?      �?      .@      3@       @      �?      @      @      �?     �K@      *@     �D@      @      5@      @      @      ,@     �D@      "@       @      (@     �A@      M@      �?       @      @      2@       @      >@      "@      @@      @      .@      �?      @      @      A@      @      @       @      ?@     �E@      �?       @      @      2@      �?      9@      @      "@      �?      @      @              @      @      @      @      @      @      .@                                      �?      @      �?       @      @      �?               @              @      �?      @      "@       @      @              &@       @      &@       @       @      �?      @              �?              @                                      @       @      �?                                      �?      �?      �?                      �?               @                                              �?      �?                                      �?      �?              @                              @                                      @      �?                                                      @              @      @                      @              @      �?      @      @              @              &@       @      &@      �?      @              �?      �?                      @               @                      �?               @              @              &@              �?              @      @                                      �?      �?      @       @               @              @       @              �?      A@      "@     @P@      @      (@       @      4@      :@      H@      @      4@      ?@     �L@     �D@      @      &@      @      0@      ,@      4@              @                                      4@      2@              @      @      0@      "@               @              @              @              @                                              @              @      @      (@      @              �?               @              @               @                                                              @              @      �?                                              @              �?                                              @                      @      @      @              �?               @              *@               @                                      4@      .@                       @      @      @              �?              @              *@              �?                                      1@      .@                      �?      @       @                              @                              �?                                      @                              �?      �?      @              �?                              ,@      "@      N@      @      (@       @      4@      @      >@      @      1@      9@     �D@      @@      @      "@      @      &@      ,@      @              9@      �?      �?       @       @      �?      (@               @      @      .@      "@              @       @      @      @       @              9@              �?              @      �?      @              @      �?       @      @              @      �?      �?              �?                      �?               @      @              @              @       @      @      @              @      �?       @      @      &@      "@     �A@      @      &@      @      (@      @      2@      @      "@      6@      :@      7@      @       @      @       @      "@      $@      @      &@       @      "@      �?      @       @      $@                      @      "@       @                      @       @      @      �?      @      8@       @       @      @       @      @       @      @      "@      2@      1@      .@      @       @       @      @      @     �p@     �C@     �c@      8@     �A@      @      J@     �x@     �{@      :@      A@     @T@     �w@     �j@       @      @@      3@     �L@      ,@     `a@      3@      O@      �?      (@       @      0@     �l@     �n@      (@      ,@      <@     �h@     �V@              @      @      1@      @     �T@      &@     �F@              &@       @      &@     �[@     �c@      @      @      2@     �]@      @@              @              "@       @     @P@      &@      :@               @       @      $@     �R@      _@      @       @      .@     @U@      ;@              @               @       @      E@      @      2@              @       @      @      C@     �Q@      @              &@     �L@      5@              @              @              7@      @      *@              @              @      =@      O@       @              @      C@      .@              �?              @              3@              @                       @              "@       @      �?              @      3@      @               @                              7@      @       @              �?              @      B@      K@      �?       @      @      <@      @                              @       @      ,@      @       @              �?              @      A@      J@                       @      6@      @                               @              "@       @                                      �?       @       @      �?       @       @      @       @                              �?       @      1@              3@              @              �?     �B@     �@@      �?      @      @     �@@      @              �?              �?              @              *@                              �?      (@      3@                      @      7@       @              �?              �?              @              *@                              �?      "@      0@                      @      3@       @              �?              �?              �?                                                      @      @                              @                                                      $@              @              @                      9@      ,@      �?      @              $@      @                                              "@              @                                      1@      @                              @                                                      �?               @              @                       @      @      �?      @              @      @                                             �L@       @      1@      �?      �?              @      ^@     �V@      @       @      $@     �S@      M@              @      @       @      @      @              �?                                      9@      @                              @      @                                                                                                      (@       @                                                                                      @              �?                                      *@      @                              @      @                                                                                                      @      @                              @      @                                              @              �?                                       @                                                                                              K@       @      0@      �?      �?              @     �W@     @U@      @       @      $@      S@      K@              @      @       @      @       @              �?                                      ;@      ,@                       @      4@      �?                                              @                                                      ,@      @                               @                                                      @              �?                                      *@      "@                       @      2@      �?                                              G@       @      .@      �?      �?              @      Q@     �Q@      @       @       @      L@     �J@              @      @       @      @     �B@       @      *@                              @     �M@     �N@      @      @       @     �C@      H@               @      @      @      @      "@      @       @      �?      �?                      "@      $@       @      @      @      1@      @              �?              �?             �_@      4@      X@      7@      7@      @      B@      e@     �h@      ,@      4@     �J@     �f@      _@       @      9@      .@      D@      "@     @T@      "@      J@      $@      @              0@      a@      d@      �?      0@      5@      \@     �O@              ,@      @      5@      @      .@      �?      (@                              �?      L@      N@              @      "@      @@      *@                              @              *@      �?      "@                              �?      I@      E@              �?      @      ?@      &@                              @              @              @                                      6@      *@                      �?      (@      @                              �?              "@      �?      @                              �?      <@      =@              �?      @      3@      @                               @               @              @                                      @      2@              @      @      �?       @                              @              �?                                                       @      @                      @              �?                              @              �?              @                                      @      *@              @              �?      �?                                             �P@       @      D@      $@      @              .@     @T@      Y@      �?      (@      (@      T@      I@              ,@      @      .@      @     �J@      @      :@      @      @              (@     �R@     �V@      �?      $@       @      K@      E@              &@      @       @      @      @       @       @                              @      2@      &@      �?              �?      (@      @               @      �?      @              H@      @      8@      @      @              @      L@     �S@              $@      @      E@     �A@              @       @      @      @      *@       @      ,@      @      �?              @      @      $@               @      @      :@       @              @              @       @      @              @                              @      @       @               @      �?      .@       @                              @      �?       @       @       @      @      �?                      @       @                      @      &@      @              @              @      �?      G@      &@      F@      *@      2@      @      4@      ?@      B@      *@      @      @@     @Q@     �N@       @      &@      (@      3@       @      ?@       @      <@      &@       @      �?      ,@      7@      >@      @      @      ,@     �G@      <@      @      @      @      @      �?       @              *@      @                      $@      @      @               @      @      .@      @              @               @              @               @       @                      @              @              �?              @      @              @                              �?              @      @                      @      @                      �?      @      (@       @               @               @              7@       @      .@      @       @      �?      @      0@      :@      @      �?      $@      @@      7@      @      �?      @      @      �?      0@      @      "@      @              �?       @      &@      ,@      @      �?      @      :@      6@      �?      �?      @      �?              @      �?      @               @               @      @      (@                      @      @      �?      @                       @      �?      .@      @      0@       @      $@      @      @       @      @      @      �?      2@      6@     �@@       @      @      "@      ,@      �?      @              @              @      �?      @      @       @      �?              @      @      3@              @              @      �?       @                                      �?       @                                      �?               @               @              @      �?      �?              @              @              �?      @       @      �?              @      @      &@              @              �?              (@      @      "@       @      @       @      @      �?      @      @      �?      ,@      1@      ,@       @              "@       @               @      @      �?       @              �?                       @      @      �?      $@      @      "@      �?              @      @              $@               @              @      �?      @      �?       @       @              @      *@      @      �?              @      @        �t�bub�r     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��30hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         4                   �2@\��
 ��?�	           ��@                            @�Q���?�           ��@                           �?8�Va���?�           ��@                          �1@7a��?�?�            px@                            �?���ٺ�?�            �j@                            @)\���h�?4             T@������������������������       �ɶ���?            �C@������������������������       �`�I\�(�?            �D@	       
                    @�`���@�?[            �`@������������������������       �d;�O���?E             Y@������������������������       ��1�O�c�?            �@@                           @Y@�}�U�?i            @f@                            �?l�Z±g�?G            �]@������������������������       ��*:��?1            �S@������������������������       �����[�?            �D@                           @�:���?"            �M@������������������������       �)\���(�?             D@������������������������       ��:�lO�?             3@                            �?�9m��?�            �v@                           @�m #�C�?�            q@                           @z�a���?l            �f@������������������������       �a��V�?H            �]@������������������������       �ėO.2��?$            �O@                            �?"3>�T�?>            �V@������������������������       ��ۘ9��?"            �G@������������������������       �Ra���i�?             F@                           @W�{w�?:            @V@                          �1@>��>��?3            @S@������������������������       �N=��� �?            �G@������������������������       ��|�j�?             >@������������������������       ��q�q�?             (@        %                   �0@�F�����?�            �r@!       "                    �?@dO�%f�?            �F@������������������������       �F]t�E�?	             &@#       $                    @�P�n#�?             A@������������������������       �h�����?             ,@������������������������       �{�G�z�?             4@&       -                    @�~�$�?�             p@'       *                    @t�/���?R            ``@(       )                    �?�l����?C            �Z@������������������������       ��;N��?             =@������������������������       ����
2��?3            @S@+       ,                    �?�&S��?             9@������������������������       �p=
ףp�?             $@������������������������       ���A���?	             .@.       1                    �?��i�$��?W            �_@/       0                    @Ӈ<��?$            �I@������������������������       �ƵHPS!�?             :@������������������������       ��D���J�?             9@2       3                    �?���=A�?3             S@������������������������       ���WV��?!             J@������������������������       �UUUUUU�?             8@5       T                    �?������?�           R�@6       E                    �?c�)�:Q�?.           ,�@7       >                    �?�oz��?F            @8       ;                     �?��MY��?o            �d@9       :                     �?���g�?C            �X@������������������������       ��Zn���?#            �H@������������������������       � A�c�]�?              I@<       =                     @o#،A��?,             Q@������������������������       ��d�����?             3@������������������������       ���Z��?            �H@?       B                     �?{S"�?�            �t@@       A                    >@F�_���?2             U@������������������������       ��j U��?,            �Q@������������������������       �s
^N���?             ,@C       D                    �?������?�            �n@������������������������       ��l����?;            �S@������������������������       ��1�&�?j             e@F       M                    �?���5h�?�           Ȉ@G       J                    @�]K޽��?�            �p@H       I                   �>@��:����?r             g@������������������������       ���$�H�?j            �d@������������������������       �����K�?             2@K       L                   �;@���Q8�?.             T@������������������������       �Ԁ�C`(�?'            �P@������������������������       ��T�6|��?             *@N       Q                   @@@�Xǰy�?H           ��@O       P                     @�j)�V�?1           �~@������������������������       ��|B���?�            �p@������������������������       ��S�~�@�?�            �k@R       S                     @      �?             D@������������������������       ��������?             4@������������������������       �R���Q�?             4@U       d                   �:@7��:�d�?�           x�@V       ]                     @}���?&           ��@W       Z                    �?ȡ@��?�           p�@X       Y                    �?��A�?�            `v@������������������������       �U�|��Q�?z            �h@������������������������       �3p�ZAJ�?g            �c@[       \                   �8@��1���?�           ��@������������������������       �)q�v9��?m           Ђ@������������������������       �Vn\1�K�?:             W@^       a                    @e�i~���?�            @q@_       `                    @L�eL��?Q            �a@������������������������       ���K����?J            �_@������������������������       �0��b�/�?             .@b       c                    @"\1&1e�?M            �`@������������������������       ��N�?�0�?             A@������������������������       ���� ��?5            @Y@e       l                    �?�,�d�S�?�            �m@f       i                    �?���,�?2            �P@g       h                   �<@�~j�t��?             9@������������������������       ��s�n_�?             *@������������������������       �9��8���?             (@j       k                   �<@/�����?"             E@������������������������       �t�@�t�?             .@������������������������       �I��D�?             ;@m       p                   �;@�Y�X\,�?g            `e@n       o                     @�|�j��?            �F@������������������������       �`Y�K�?             :@������������������������       �X�3�R�?	             3@q       r                     �?��q�5A�?L            �_@������������������������       �[������?!            �J@������������������������       �K�(N��?+            @R@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       �|@     @S@     `v@      ?@     �Q@      :@      T@     ��@     H�@     @R@     @V@     �c@     x�@     �z@      3@     @Q@      K@     �_@      L@     �^@      @     �Q@      �?      @              ,@     �q@     �j@      (@      $@      ;@     �f@     �S@               @      @      2@      @      S@      �?     �B@              �?              (@      m@      e@      $@      @      .@     �`@     �H@              @      �?       @      �?      D@      �?      (@                               @     �b@      W@               @      @      P@      6@                              �?              6@              @                               @     �X@      E@                      @     �A@      @                              �?              @              @                                     �D@      &@                              0@      �?                              �?              @              @                                      8@      @                              @      �?                                              @                                                      1@      @                              *@                                      �?              .@              �?                               @     �L@      ?@                      @      3@      @                                              "@              �?                               @      G@      8@                      @      (@      @                                              @                                                      &@      @                              @       @                                              2@      �?       @                                     �I@      I@               @      @      =@      0@                                              @      �?      @                                     �@@     �D@                              3@      (@                                              @      �?      �?                                      3@      7@                              2@      &@                                              �?              @                                      ,@      2@                              �?      �?                                              (@              �?                                      2@      "@               @      @      $@      @                                              $@                                                      @       @               @      @      "@      @                                               @              �?                                      *@      �?                              �?      �?                                              B@              9@              �?              $@     �T@     @S@      $@      @      "@      Q@      ;@              @      �?      @      �?      =@              7@              �?              @     �G@      P@       @      @       @     �J@      1@              @      �?      @      �?      *@              7@              �?              @      7@      F@       @      @      @     �D@      $@              �?      �?      @      �?      $@              &@              �?                      1@      1@      @      @      @     �@@      "@              �?      �?      @      �?      @              (@                              @      @      ;@       @              �?       @      �?                                              0@                                              @      8@      4@                      �?      (@      @              @              @              @                                               @      0@      *@                      �?      @      @                              �?              *@                                               @       @      @                              @      @              @              @              @               @                              @      B@      *@       @              �?      .@      $@                                              @               @                              @     �A@      $@       @              �?      &@       @                                              @                                              �?      0@       @                      �?      "@       @                                              �?               @                               @      3@       @       @                       @                                                       @                                                      �?      @                              @       @                                              G@      @      A@      �?      @               @     �I@      G@       @      @      (@      H@      >@              @      @      $@       @      ,@      �?      @                                      .@      @                              @      @                                              @                                                      @       @                               @                                                      $@      �?      @                                      (@       @                              �?      @                                              "@      �?                                              �?                                      �?       @                                              �?              @                                      &@       @                                      @                                              @@      @      ?@      �?      @               @      B@      E@       @      @      (@     �F@      9@              @      @      $@       @      (@       @      4@              @               @      .@      0@       @      @      @      @@      (@                              @              (@       @      @              @              �?      (@      .@       @      @      @      ;@      (@                              @              @      �?                                              @      �?       @              @      (@                                      @              "@      �?      @              @              �?       @      ,@              @       @      .@      (@                              @                              .@                              �?      @      �?                              @                                                                      @                                       @      �?                                                                                                       @                              �?      �?                                      @                                                      4@      �?      &@      �?                              5@      :@               @      @      *@      *@              @      @      @       @      @              @                                      (@      *@                       @      @      @               @               @              @               @                                       @      @                       @      �?      @                              �?              @              �?                                      @       @                              @                       @              �?              ,@      �?       @      �?                              "@      *@               @      @      @      "@               @      @      �?       @      *@              @      �?                              @       @              �?      @       @       @                      @      �?       @      �?      �?      @                                      @      @              �?      �?      @      �?               @                             u@      R@     �q@      >@     �P@      :@     �P@     `o@      w@     �N@     �S@     @`@     �{@     �u@      3@     �N@      I@      [@     �J@     �`@      B@      b@      (@      B@      5@      E@     �L@     �]@      :@     �M@     �P@     �e@     �f@      ,@     �A@      C@      L@     �E@     �P@      "@     �I@       @       @      @      2@      >@      P@      @      6@      9@     �U@     �I@      @      "@      0@      (@      2@      3@      @      .@                       @              .@      @@      @       @      @     �D@      *@               @      �?       @      @      2@      @       @                                      @      3@      �?      @      @      6@      "@              �?               @      �?      @       @      @                                       @      $@               @       @      ,@       @              �?               @      �?      &@       @      @                                      @      "@      �?      @      �?       @      @                                              �?              @                       @              $@      *@       @       @      @      3@      @              �?      �?              @      �?              @                                      @      �?      �?      �?              @                                                                      @                       @              @      (@      �?      �?      @      ,@      @              �?      �?              @      H@      @      B@       @       @      �?      2@      .@      @@              ,@      3@      G@      C@      @      @      .@      $@      ,@      &@      �?      $@               @              "@      @      "@              @      �?      "@      @              �?      @      @      @      &@      �?      $@               @               @      @      @              @      �?      "@      @              �?               @      @                                                      �?               @               @                      @                      @       @             �B@      @      :@       @      @      �?      "@      &@      7@              "@      2@     �B@      ?@      @      @      &@      @      @      ,@      �?      ,@              �?                      @       @               @      �?      ,@      $@               @              @      �?      7@      @      (@       @      @      �?      "@      @      .@              @      1@      7@      5@      @      @      &@      �?      @     �P@      ;@     @W@      $@      <@      2@      8@      ;@      K@      7@     �B@      E@     �U@     @`@      &@      :@      6@      F@      9@     �B@       @      >@              "@      �?      @      ,@      1@      @      (@      ,@      G@     �B@               @      @      $@       @      6@       @      ,@              @      �?      @      $@      ,@      �?      "@      (@     �A@      =@              @      �?      "@      @      6@       @      (@              @      �?      @      $@      ,@      �?      @      @     �A@      =@              @      �?      @      @                       @              @                                              @      @                                               @              .@              0@               @              @      @      @      @      @       @      &@       @              @       @      �?      @      &@              ,@                                      @      @      @      @       @      "@       @              @       @      �?      @      @               @               @              @                                               @                                                      =@      3@     �O@      $@      3@      1@      2@      *@     �B@      2@      9@      <@      D@     @W@      &@      2@      3@      A@      1@      =@      3@     �J@       @      3@      0@      2@      *@      B@      1@      8@      4@      D@     @W@      @      2@      ,@     �@@      *@      0@      @      9@      @      @      �?      @      *@      6@      .@      ,@      "@      4@      L@      @      .@      *@      2@      @      *@      *@      <@      @      (@      .@      ,@              ,@       @      $@      &@      4@     �B@      �?      @      �?      .@       @                      $@       @              �?                      �?      �?      �?       @                      @              @      �?      @                      @                                              �?      �?              @                                      @      �?       @                      @       @              �?                                      �?      �?                      @                               @     �i@      B@     �a@      2@      >@      @      8@     @h@     �o@     �A@      4@     �O@     �p@     �d@      @      :@      (@      J@      $@     �g@      :@     @\@      .@      9@      �?      2@      g@     @m@      .@      (@      F@     �m@     `a@      @      6@      @     �C@      @     @d@      (@     �W@      "@      ,@              &@     �b@     `j@      &@      (@      >@     @g@     �Z@              &@      @      >@       @      G@      @      ?@               @              @     �F@     @Y@      @              2@     �K@     �A@              @      �?       @      �?      <@      @      .@                                      5@     �M@      �?              (@      E@      (@              @                              2@              0@               @              @      8@      E@       @              @      *@      7@               @      �?       @      �?      ]@      @     �O@      "@      (@              @     �Y@     �[@       @      (@      (@     ``@     �Q@              @       @      <@      �?     @Z@      @      J@      "@      $@              @     @W@     �Y@       @      $@      &@     �Z@      N@              @       @      3@      �?      &@              &@               @              �?      $@       @               @      �?      9@      &@              �?              "@              ;@      ,@      3@      @      &@      �?      @     �B@      7@      @              ,@      I@     �@@      @      &@       @      "@      @      ,@      $@      *@      @       @      �?       @      .@      (@                      (@      9@      (@              @      �?      @      @      @      $@      (@      @       @      �?       @      .@      &@                       @      9@      &@              @      �?      @      @      @              �?                                              �?                      @              �?                              �?              *@      @      @      �?      @              @      6@      &@      @               @      9@      5@      @       @      �?      @              @                      �?                      �?      "@      @                              @      &@                              �?              "@      @      @              @              @      *@      @      @               @      6@      $@      @       @      �?      @              .@      $@      >@      @      @      @      @      "@      2@      4@       @      3@      A@      <@      �?      @      @      *@      @       @       @      @      �?       @              �?      @      @      @      @      @      1@      @              @              �?              �?      �?                                      �?      @      @                       @      $@                       @                              �?                                              �?      @       @                       @      @                                                              �?                                                      @                              @                       @                              @      �?      @      �?       @                      @       @      @      @       @      @      @              �?              �?               @      �?              �?      �?                      �?              �?       @              @                                      �?              @              @              �?                      @       @       @      �?       @       @      @              �?                              @       @      :@       @      @      @      @       @      &@      1@      @      .@      1@      8@      �?      �?      @      (@      @      �?      �?      (@                      �?      @       @       @      �?               @       @      ,@              �?                      �?      �?      �?      (@                      �?      �?       @              �?              �?       @      @              �?                                                                              @               @                      �?              &@                                      �?      @      @      ,@       @      @      @                      "@      0@      @      *@      .@      $@      �?              @      (@      @               @      $@              @      �?                      �?      &@      @       @      $@      @                      @       @      �?      @      @      @       @               @                       @      @       @      &@      @      @      �?              @      $@       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ=�(hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKmhnh4h7K ��h9��R�(KKm��hu�B�         4                   �2@��>��?�	           ��@                            @݇	I��?�           (�@                           �?�V��	
�?�           �@                           �?#��k�4�?�            `q@                            �?�١A���?g             f@                           @��hJ,�?M             a@������������������������       ���9�-��?             G@������������������������       ��:�^���?2            �V@	       
                   �0@`�I\�(�?            �D@������������������������       �X�<ݚ�?             "@������������������������       �     ��?             @@                          �0@쁟�Y�?@            @Y@������������������������       ���Q���?             4@                            �?,�D���?5            @T@������������������������       �E�T���?'            �M@������������������������       �HN�zv�?             6@                          �0@*�����?           �z@                           @خ�u��?3            �R@                           @r�qG�?              H@������������������������       �Z0Rb�?             =@������������������������       �ԍx�V�?             3@                           �?���+�w�?             :@������������������������       �x9/���?
             ,@������������������������       ��������?	             (@                           �?�P~^T�?�             v@                            �?���>4��?             <@������������������������       �0��b�/�?             .@������������������������       �"���c��?             *@                           @1j۬�8�?�            `t@������������������������       ��%���?N            �_@������������������������       ��@���=�?            �h@        '                   �0@���|��?�            �t@!       $                    �?�IF�E��?&            �P@"       #                    �?�>�\��?             ?@������������������������       �r�q��?             (@������������������������       ����.�?
             3@%       &                    @4և����?            �A@������������������������       �d}h���?
             ,@������������������������       ���{�~�?             5@(       /                    @;�O�?�            `p@)       ,                    �?] ܢm��?�            �j@*       +                    @��Jr�?A            �X@������������������������       ��sly47�?3            �R@������������������������       �9��8���?             8@-       .                    �?��}���?I            @\@������������������������       ���|��?             >@������������������������       �K�m_8�?8            �T@0       1                   �1@a��+e�?             I@������������������������       ��8��8��?             (@2       3                    �?��	"P�?             C@������������������������       ��eP*L��?             6@������������������������       �      �?	             0@5       T                   �:@`�9���?"           ~�@6       E                     @�*�mn{�?�           �@7       >                   �5@a���8�?           h�@8       ;                    �?��:�Ļ�?            �@9       :                    @H�H�Κ�?�             q@������������������������       �     ��?P             `@������������������������       ����I��?d            @b@<       =                     �?FJJՃ��?N           ��@������������������������       �ά�wc7�?           �y@������������������������       �T	<�v�?L            �]@?       B                    �?k�p�:|�?           ��@@       A                   �6@L�_U���?�            Px@������������������������       ���J��z�?B            �Z@������������������������       �H)Ꟶ�?�            �q@C       D                    @���N��?           {@������������������������       ����Bo�?t            @e@������������������������       ��wG2��?�            pp@F       M                    @R������?�           ��@G       J                   �6@�{ǃ}��?           �z@H       I                    �?u����?�             q@������������������������       ��ݟ�ߦ�?Y            �a@������������������������       ����*���?U            @`@K       L                   �9@���m�?]             c@������������������������       �\HC��!�?S            `a@������������������������       �^N��)x�?
             ,@N       Q                    �?Lݿ��!�?�            �p@O       P                    @�������?E            �Y@������������������������       �9��8���?             8@������������������������       ����Y� �?3            �S@R       S                    �?Ns�g �?l            �d@������������������������       �|>�+78�?            �A@������������������������       ��IJ6��?S            @`@U       d                   @@@ĦE���?a           ��@V       ]                    �?���4}�?$           p}@W       Z                    �?~�-����?s            �f@X       Y                     @�����?$            �L@������������������������       �3�E��?            �C@������������������������       �)O���?
             2@[       \                    �? AR�A�?O             _@������������������������       ��5�����?(            @P@������������������������       ���˰���?'            �M@^       a                    @M�%�k�?�             r@_       `                     �?�O��Oz�?�             n@������������������������       �6�9�?O            �_@������������������������       �n��jE?�?H            �\@b       c                     �?W�/�'�?             I@������������������������       ��8	���?
             3@������������������������       �E���|,�?             ?@e       j                    �?�cp��?=            �V@f       g                    �?bΊx��?'             M@������������������������       ��������?             $@h       i                     @�8��8��?!             H@������������������������       ��L-���?             ;@������������������������       �lv�"��?             5@k       l                   @A@     ��?             @@������������������������       ��|�j��?             .@������������������������       �ZZZZZZ�?             1@�t�bh�h4h7K ��h9��R�(KKmKK��h��B�@       P|@     �R@     �u@      =@      U@      3@     �V@     �@     ��@     @T@      Q@     �e@     ��@     �{@      *@      H@      J@      `@      M@     @]@      @      Q@              @              ,@     �p@      l@      @      "@     �A@     `c@     �T@              "@      @      :@      @     �Q@      @      @@                               @     `j@      e@      @      @      :@     @Y@      I@              @      @      &@      �?      ?@              @                                      [@      Q@       @       @      $@      B@      (@              �?              @      �?      .@                                                     �U@      D@              �?      @      4@       @                                               @                                                     @R@      8@              �?      @      0@       @                                              @                                                      :@      @              �?      @      @      @                                               @                                                     �G@      5@                       @      *@      @                                              @                                                      ,@      0@                              @                                                       @                                                      @                                      �?                                                      @                                                       @      0@                              @                                                      0@              @                                      5@      <@       @      �?      @      0@      @              �?              @      �?      @              �?                                      @      &@                                                                                      &@              @                                      2@      1@       @      �?      @      0@      @              �?              @      �?      "@               @                                      "@      *@              �?      @      ,@       @              �?              @      �?       @              �?                                      "@      @       @                       @       @                                              D@      @      <@                               @     �Y@     @Y@      @      @      0@     @P@      C@              @      @       @              @              �?                                      4@     �@@                       @      "@       @                               @              @              �?                                      &@      =@                              @                                                      @              �?                                       @      ,@                              @                                                                                                              @      .@                              �?                                                       @                                                      "@      @                       @      @       @                               @              �?                                                      @      @                              @                                                      �?                                                      @      �?                       @      �?       @                               @             �A@      @      ;@                               @     �T@      Q@      @      @      ,@      L@      B@              @      @      @              @              @                              �?      �?      &@                      �?      �?      �?                                              @              @                              �?              @                                      �?                                               @                                                      �?       @                      �?      �?                                                      >@      @      4@                              @     �T@     �L@      @      @      *@     �K@     �A@              @      @      @              @      @      $@                              @      <@      =@      �?      �?       @      <@      $@                              @              7@              $@                              @      K@      <@       @       @      &@      ;@      9@              @      @      @              G@              B@              @              @      L@      L@              @      "@      K@     �@@              @      �?      .@       @      ,@              @               @                      8@      $@                               @      @                                              @               @                                      (@       @                              @      �?                                               @               @                                      @                                      �?      �?                                              @                                                      @       @                              @                                                      @              @               @                      (@       @                              �?       @                                              @                                                      @       @                              �?      �?                                                              @               @                      "@      @                                      �?                                              @@              ?@              @              @      @@      G@              @      "@      G@      >@              @      �?      .@       @      ;@              .@              @              @      6@     �D@              @      "@      B@      >@              @      �?      .@       @      *@              @                              @      1@      3@                      @      4@       @              @              @              (@              @                              @      0@      @                      @      1@       @               @              @              �?              @                                      �?      ,@                              @                      �?              �?              ,@               @              @                      @      6@              @      @      0@      6@                      �?      "@       @      @               @                                      �?      @               @               @       @                              @       @       @              @              @                      @      0@               @      @      ,@      4@                      �?       @              @              0@                              @      $@      @                              $@                      �?                              @                                                      �?       @                              @                      �?                              �?              0@                              @      "@      @                              @                                                                      .@                              @      @                                      �?                                                      �?              �?                                      @      @                              @                                                      u@     �Q@     pq@      =@     �S@      3@      S@     �n@     Py@      S@     �M@     �a@     |@     �v@      *@     �C@     �F@     �Y@     �K@     �q@      D@     �k@      4@     �H@      &@     �K@     `l@     w@     �F@      G@     �Z@     @x@      s@      @      <@      9@     �P@      :@      j@      0@      d@      @      =@      @      @@     �f@     �q@      ;@      A@     �P@     pq@     �h@      @      4@      *@     �H@      ,@     �[@      @     �Q@       @      (@               @     �^@     �d@      @      &@      >@     �`@     �T@               @      @      <@      "@      :@      �?      .@              @               @      C@     @T@              @      (@      G@      C@               @      �?       @      @      .@               @                                      @      G@               @      @      1@      7@               @               @              &@      �?      @              @               @      ?@     �A@               @      @      =@      .@                      �?              @     @U@      @     �K@       @      "@              @      U@     @U@      @      @      2@     �U@     �F@              @       @      :@      @     @Q@       @      G@       @      @              @      J@      N@      @      @      1@     �P@      B@              @       @      6@      @      0@      �?      "@               @                      @@      9@      �?              �?      3@      "@                              @             �X@      (@     �V@      @      1@      @      8@     �N@     �]@      6@      7@      B@     `b@     @\@      @      (@      $@      5@      @     �G@      @      G@      �?      @              @     �@@      U@      @      @      0@      N@     �L@               @      @      @      �?       @      �?      2@              @              �?       @      ?@              �?      �?      4@      (@                       @      �?             �C@      @      <@      �?      �?              @      9@     �J@      @      @      .@      D@     �F@               @      �?      @      �?     �I@      @     �F@      @      *@      @      1@      <@     �A@      1@      3@      4@     �U@      L@      @      @      @      ,@      @      ;@      @      3@      �?                      @      7@      2@      @      @      @      :@      5@      �?       @       @      @      �?      8@       @      :@       @      *@      @      ,@      @      1@      *@      *@      ,@     �N@     �A@      @       @      @       @      @      S@      8@     �N@      ,@      4@       @      7@      F@      U@      2@      (@      D@     @[@      [@      �?       @      (@      2@      (@     �I@      ,@      <@      (@      .@      @      @      @@      O@       @      @      2@      R@     �Q@              @      @      &@      @      C@      &@      0@      @      $@       @       @      ;@      =@      @      @      @     �K@      H@              @               @      @      1@              @               @      �?              6@      1@               @              A@     �@@               @              @      @      5@      &@      (@      @       @      �?       @      @      (@      @       @      @      5@      .@              @              @       @      *@      @      (@       @      @      @      �?      @     �@@      @              *@      1@      7@              �?      @      @              "@      @      (@       @      @      @      �?      @      @@      @              "@      1@      7@                      @      @              @                               @      �?                      �?                      @                              �?      �?                      9@      $@     �@@       @      @       @      4@      (@      6@      $@       @      6@     �B@     �B@      �?       @      @      @      @      @       @      $@       @       @      �?       @      "@      &@              @      &@      6@      $@              �?      �?      @              �?               @      �?                      @       @      @              �?      �?       @                                                      @       @       @      �?       @      �?      @      @      @              @      $@      4@      $@              �?      �?      @              4@       @      7@              @      �?      (@      @      &@      $@      @      &@      .@      ;@      �?      �?      @      @      @      "@      �?       @                              �?      �?              @       @              @      �?                      @              @      &@      @      5@              @      �?      &@       @      &@      @       @      &@      (@      :@      �?      �?              @      @     �I@      >@     �L@      "@      =@       @      5@      1@      B@      ?@      *@      A@     �N@      N@       @      &@      4@      B@      =@     �F@      <@     �I@      @      9@      @      2@      1@      A@      3@      "@      6@      L@      N@      �?      @      .@      A@      6@      ;@      &@      &@              "@              @      *@      0@      @      @      @      ?@      3@              �?      @      $@      "@      ,@      @      �?              �?              �?              &@              �?      �?      (@      @                       @                       @      @                      �?              �?              &@              �?      �?      @      @                       @                      @       @      �?                                                                               @      �?                                              *@      @      $@               @              @      *@      @      @      @      @      3@      (@              �?      @      $@      "@      "@       @      @               @              @              @       @      �?      @      @      @                      @       @      "@      @      @      @              @                      *@      �?      �?      @              (@      @              �?               @              2@      1@      D@      @      0@      @      *@      @      2@      0@       @      2@      9@     �D@      �?      @      $@      8@      *@      *@      ,@      :@      @      0@      @      *@      @      2@      *@       @      0@      6@     �B@      �?      @      @      ,@      *@      "@      @      5@      @      @      �?      @      @      @      @      �?      $@      0@      2@              @      �?       @       @      @      @      @              "@      @      @              &@      @      �?      @      @      3@      �?              @      (@      &@      @      @      ,@      �?                              �?              @               @      @      @                      @      $@                               @                                      �?              �?               @              �?                      @       @              @      @      (@      �?                                               @                      @      @                               @              @       @      @      @      @      @      @               @      (@      @      (@      @              @      @      @       @      @      @              @      @      @               @              �?      @      @      $@                      @      @      @       @      @                      �?       @       @                                      @      �?                                              �?                      @               @       @       @               @              �?      �?      @      $@                      @      @      @       @      @      �?               @      �?       @                              �?      �?      @      @                              �?      @       @      @       @                      �?                       @                                      @                      @      @                       @      @       @      @                      @      �?              �?       @               @      @                      �?      �?               @      �?      �?                                                              @              �?      @                      �?      �?               @       @      �?      @                      @      �?              �?      @              �?                                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�a�KhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKyhnh4h7K ��h9��R�(KKy��hu�Bx         :                   �4@V�e4Ħ�?�	           ��@                          �0@���>Y�?�           4�@                            �?�
��P�?�             l@                           @��e�?R            ``@                           @�|WB�p�?<            �V@                           �?Vx�����?+            @Q@������������������������       �J��LQ�?             7@������������������������       ��z�l/��?             G@	       
                     �?�0�~�4�?             6@������������������������       ��8��8��?	             (@������������������������       ���(\���?             $@                           �?�G�z�?             D@������������������������       �X�Cc�?	             ,@                           @�]�`��?             :@������������������������       �r�q��?             (@������������������������       �*x9/��?             ,@                           �?Ҫ~�Z��?7            �W@                           �?��X��?             <@������������������������       ���!pc�?             &@������������������������       ��l� {�?
             1@                            @IJ�}�o�?&            �P@                           �?��Hx��?             B@������������������������       ���?�v��?             =@������������������������       ��$I�$I�?             @                           �?�K~���?             >@������������������������       ���>4և�?             ,@������������������������       �     ��?	             0@       +                     @�'����?�           ��@       $                    �?[6L5��?�           �@       !                   �3@X������?�            �q@                           �1@��gL�?�            �k@������������������������       ��z�� �?-            �P@������������������������       �zW&Hѩ�?d            @c@"       #                    �?�$ğӯ�?&            �O@������������������������       �;U��j�?             =@������������������������       �7��d��?             A@%       (                    @J��$B��?
           X�@&       '                    @��3����?�           ��@������������������������       �5yy8,�?l            `c@������������������������       �t��'���?*           P}@)       *                   �3@������?t            `g@������������������������       �vQ���
�?Y            `b@������������������������       �q=
ףp�?             D@,       3                    @|��~F�?;           P~@-       0                    @���y�?�            �v@.       /                    @Ý�y�?�            pr@������������������������       �"K�� 2�?�            �k@������������������������       ��W#����?3            �R@1       2                   �3@G���U�?'             Q@������������������������       �D̏S�?            �I@������������������������       �v�f��?
             1@4       7                   �3@���7�H�?M            �^@5       6                    @fP*L��?7             V@������������������������       �h�2�q�?1            �S@������������������������       ���Q��?             $@8       9                    �?{�/��>�?             A@������������������������       �'�%����?             7@������������������������       �F]t�E�?             &@;       Z                    @�#���@�?2           x�@<       K                    �?sѪ�]e�?W           ̔@=       D                   �9@�������?a            �@>       A                   �7@�6��3��?�            @u@?       @                   �6@2(��F�?�            �l@������������������������       �C]���?j             d@������������������������       �$،A���?-             Q@B       C                    @��c��-�?N            �[@������������������������       ��*F4���?H            @Y@������������������������       �p=
ףp�?             $@E       H                   �=@[��K���?|            �i@F       G                   �;@T(�b�2�?U            @a@������������������������       ���֢���?,            �R@������������������������       ��ܤ��?)            �O@I       J                    @]t�E�?'            �P@������������������������       ��j�=F?�?             E@������������������������       �9��8���?             8@L       S                   �>@�B,��?�           ��@M       P                    �?�D�Y/e�?�           �@N       O                   �7@X9��v��?�             i@������������������������       ��p.gR �?A            @W@������������������������       �|U����?A            �Z@Q       R                    �?U���=s�?C           �@������������������������       ���w�m�?�            `v@������������������������       �,<���?b            `b@T       W                    �?Y�3�a�?1            �T@U       V                     �?<�:�k+�?$             O@������������������������       ��	"P7��?	             3@������������������������       �J1|w���?            �E@X       Y                     �?�(\����?             4@������������������������       ���"e���?             "@������������������������       ��ˠT�?             &@[       j                    �?p�>���?�           H�@\       c                    �?d!Y��?�             w@]       `                    @����B�?J             \@^       _                   �6@��(\���?             D@������������������������       ��q�q�?	             (@������������������������       �^N��)x�?             <@a       b                    @X�<ݚ�?1             R@������������������������       ��#��Z=�?             6@������������������������       ��*��	�?"             I@d       g                    @    @!�?�             p@e       f                   �=@�Y�Y�?^            �e@������������������������       ����}4��?X             d@������������������������       �r�q��?             (@h       i                   �5@��� ���?4            �T@������������������������       �+7����?             7@������������������������       �������?'             N@k       r                    @M����?�            �y@l       o                    @YqG9�{�?�            `n@m       n                   �6@���2�?Q            `a@������������������������       ��0`�Ī�?             M@������������������������       ���oo�5�?2            @T@p       q                    @؉�؉��?>             Z@������������������������       ��X�A��?            �D@������������������������       �u���?'            �O@s       v                     @Z ����?p            �d@t       u                    �?i��b�I�?Q            �]@������������������������       ����D=�?             ?@������������������������       ��A�0�~�?>             V@w       x                   �8@��L��z�?            �G@������������������������       �����S��?             <@������������������������       ������?             3@�t�bh�h4h7K ��h9��R�(KKyKK��h��B�G        }@     �W@     �w@     �A@     �U@      ?@      R@     ��@     ��@      M@     �S@      d@     ��@     �y@      0@     @P@     �B@      `@      S@     @n@      ,@     �`@      "@      4@              (@     �w@     �v@      ,@      9@      N@     �r@     �b@              2@      @      D@      0@     �A@       @      &@               @                     @T@      M@                              =@      @                              �?              6@              "@                                     �B@     �E@                              1@       @                              �?              $@              @                                      5@     �B@                              0@                                                      $@              @                                      3@      2@                              .@                                                      @              @                                      @      @                              �?                                                      @              �?                                      (@      *@                              ,@                                                                                                               @      3@                              �?                                                                                                              �?      &@                                                                                                                                              �?       @                              �?                                                      (@               @                                      0@      @                              �?       @                              �?              �?               @                                      $@      �?                                                                                      &@                                                      @      @                              �?       @                              �?               @                                                      @      @                              �?       @                              �?              "@                                                      @       @                                                                                      *@       @       @               @                      F@      .@                              (@      @                                               @       @                                              $@      �?                              @       @                                                                                                      @                                      @       @                                               @       @                                              @      �?                              �?                                                      @               @               @                      A@      ,@                              @       @                                               @                                                      7@      @                              @       @                                              �?                                                      3@      @                              @                                                      �?                                                      @                                               @                                              @               @               @                      &@      "@                              @                                                       @                                                      @      @                              @                                                      �?               @               @                       @      @                                                                                     �i@      (@      _@      "@      2@              (@     pr@     @s@      ,@      9@      N@     q@      b@              2@      @     �C@      0@      a@      @     �P@      @      @              $@     �m@     @n@      $@      ,@      D@     �g@     �V@              *@      @      0@      $@      G@      �?      9@       @      @              �?      E@     �H@      @      @      .@     �G@      7@              @              $@      @     �A@      �?      6@       @      @              �?     �B@      D@      @      @      *@      =@      ,@              �?               @      @      "@              @              @                      &@      @       @       @      @      ,@      @                              �?      @      :@      �?      2@       @                      �?      :@     �@@      @      @      @      .@      $@              �?              @      �?      &@              @                                      @      "@                       @      2@      "@              @               @      �?      @              �?                                      @      @                              "@      @                                      �?      @               @                                      �?       @                       @      "@      @              @               @             �V@      @     �D@      @      @              "@     �h@      h@      @      "@      9@     �a@      Q@              "@      @      @      @     �O@      �?      <@      �?      �?              @     `e@      d@       @      "@      0@     @Y@      K@              @       @      @      @      9@              @      �?      �?              @     �B@     �E@                      @      *@      1@              �?      �?      �?      �?      C@      �?      6@                              �?     �`@     @]@       @      "@      (@      V@     �B@               @      �?       @      @      ;@      @      *@       @       @              @      :@     �@@      @              "@      D@      ,@              @       @      @              7@      @      "@       @                      @      5@      <@      @               @      7@      *@              @       @      @              @              @               @                      @      @                      �?      1@      �?              �?                             �Q@      @      M@      @      (@               @      L@     �P@      @      &@      4@     @U@      K@              @      �?      7@      @      K@      @      G@      @      (@               @      H@     �G@               @      &@      P@     �E@              @      �?      "@      @     �D@      @      B@      @      (@               @      A@      E@               @      "@     �M@      ?@               @              @      @     �B@      @      ;@       @      (@               @      3@      >@               @      @      D@      7@               @              @      @      @       @      "@      �?                              .@      (@                      @      3@       @                                              *@       @      $@                                      ,@      @                       @      @      (@              �?      �?       @      �?      &@       @      @                                      (@       @                       @      @      "@              �?      �?       @      �?       @              @                                       @      @                                      @                                              1@              (@      �?                               @      3@      @      @      "@      5@      &@               @              ,@      �?      ,@               @      �?                              @      3@       @      @      @       @      @               @              $@      �?      ,@               @      �?                              @      0@       @      @      @      @      @               @              $@      �?                                                                      @                      @      @                                                      @              @                                      �?               @               @      *@      @                              @              @              @                                      �?               @                      &@       @                                                                                                                                       @       @      @                              @             �k@      T@     �n@      :@     �P@      ?@      N@     �c@      n@      F@      K@     @Y@     q@     @p@      0@     �G@      @@     @V@      N@     @`@     �J@      e@      7@      I@      =@      D@      I@     �`@      @@     �E@      R@     `b@     �f@       @      B@      8@      P@     �H@     @Q@      5@     �Q@      @      *@      @      2@      ;@     �R@      @      2@      6@      S@      Q@              .@      "@      (@      2@      D@      &@     �G@      @       @      @      $@      4@      O@              @      2@     �F@      D@              "@      @      @      @     �B@      @      C@      @      @      @      @      ,@     �A@              @      &@      @@      7@              @      �?       @      �?      4@      @      >@      @      @      @      @      "@      9@               @      @      8@      5@              @               @      �?      1@       @       @                              �?      @      $@              @      @       @       @              @      �?                      @      @      "@               @       @      @      @      ;@              �?      @      *@      1@              @      @      @      @      @      @      @               @       @      @      @      ;@              �?      @      @      1@              @      @      @      @                       @                                                                      �?      @                                                      =@      $@      8@      �?      @               @      @      *@      @      &@      @      ?@      <@              @      @      @      ,@      2@      $@      2@      �?      �?              @      @       @               @      �?      <@      6@              @      @      @      $@      (@      @      &@      �?                       @              @                      �?      3@      @              @      @      @      @      @      @      @              �?               @      @      @               @              "@      0@                                      @      &@              @              @              @       @      @      @      "@      @      @      @              @              @      @      &@                                                       @       @      @      "@       @       @      @              @              �?      @                      @              @              @              @                      �?      �?      @                               @             �N@      @@     �X@      3@     �B@      8@      6@      7@     �L@      =@      9@      I@     �Q@      \@       @      5@      .@      J@      ?@     �M@      @@     @V@      $@     �@@      3@      6@      6@     �I@      2@      5@     �D@     �Q@     @[@       @      3@      (@      I@      :@      8@      @      9@              "@      @       @      $@      $@      @      @      "@     �B@      ;@              @      @      0@      @      ,@      �?      2@              �?              �?      @      @       @      @      @      1@      "@              �?      �?      @      @      $@      @      @               @      @      �?      @      @      @              @      4@      2@              @       @      "@       @     �A@      :@      P@      $@      8@      0@      4@      (@     �D@      *@      2@      @@     �@@     �T@       @      ,@      "@      A@      4@      5@      5@     �F@      "@      5@      $@      .@       @      5@      $@      ,@      9@      2@     �O@       @      (@      "@      4@      ,@      ,@      @      3@      �?      @      @      @      @      4@      @      @      @      .@      3@               @              ,@      @       @              "@      "@      @      @              �?      @      &@      @      "@      �?      @      @       @      @       @      @       @               @      @      @      @                      @      @      @       @                      @       @       @      �?      @                      @      @               @                                              @                              �?              �?       @       @              @      �?      @      @                      @      @      @      @                      @      �?       @              @                      �?      @                              �?               @              �?      �?      @                      �?      �?                                                                                      @                      �?       @                      �?      �?                              �?      @                              �?              @              �?              �?                                              W@      ;@     @S@      @      1@       @      4@     @[@     @[@      (@      &@      =@     �_@      T@       @      &@       @      9@      &@      B@      $@      8@              $@              "@     �O@     �Q@      @      @      1@      P@      B@              @      �?      "@      @      3@       @      @               @              @      "@     �A@      �?      @       @      5@      "@                                              &@      �?                       @              @              $@      �?               @       @      �?                                               @      �?                                       @              @                              @                                                      "@                               @               @              @      �?               @      @      �?                                               @      �?      @                                      "@      9@              @              *@       @                                               @              @                                      @      @              @              @      @                                              @      �?      �?                                      @      5@              �?              "@      @                                              1@       @      4@               @              @      K@     �A@      @       @      .@     �E@      ;@              @      �?      "@      @      $@      @      (@              @              @     �D@      :@              �?      @      B@      2@              @      �?      @      �?      $@      @      (@               @              @     �D@      8@              �?      @      B@      *@               @      �?      @      �?                                      @                               @                                      @              �?                              @      @       @               @                      *@      "@      @      �?      $@      @      "@              @              @       @                      @               @                      @      @                      @      �?                                      �?              @      @      @                                      @      @      @      �?      @      @      "@              @              @       @      L@      1@     �J@      @      @       @      &@      G@     �C@       @      @      (@      O@      F@       @      @      @      0@       @      ?@      *@      8@       @      @      �?      @      A@     �@@      @      @      @      E@      8@      @      @      �?      @              3@      &@      3@                      �?      @      <@      *@      @      �?      @      .@      .@      �?       @      �?      @              *@              @                               @      9@      @                      @      �?      @                                              @      &@      .@                      �?      �?      @      "@      @      �?      �?      ,@      "@      �?       @      �?      @              (@       @      @       @      @               @      @      4@      @      @       @      ;@      "@       @       @              @              $@               @       @                              @      @              @       @      @      @               @              �?               @       @      @              @               @       @      1@      @                      4@      @       @                       @              9@      @      =@      �?      @      �?      @      (@      @       @              @      4@      4@      @      �?      @      $@       @      1@              :@      �?      @              @      &@      @       @              @      (@      .@              �?      @      @       @      @              �?                               @      $@      �?      �?                      @      @                                      @      (@              9@      �?      @               @      �?      @      �?              @      "@      &@              �?      @      @      @       @      @      @              �?      �?       @      �?       @                       @       @      @      @                      @               @       @       @              �?                      �?      �?                              @       @      @                       @                       @      �?                      �?       @              �?                       @      @      @                              @        �t�bub�2     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ| '"hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKkhnh4h7K ��h9��R�(KKk��hu�Bh         :                     @��%��?�	           ��@                           �?����G�?�           ��@                          �4@	����?c            �@                           @N<4����?�            �t@                          �3@a����?�             r@                            �?z%�u���?�             m@������������������������       �UZP�Q��?Q            �`@������������������������       ���D���?C            �X@	       
                    @����X�?%            �L@������������������������       �Ɲ N&��?            �F@������������������������       ���8��8�?
             (@                          �2@�F<�A+�?             C@������������������������       �Ɓ�r�z�?
             3@������������������������       �Dy�5��?	             3@                          �<@z}-�_�?�           ��@                          �5@�M?���?N           0�@                           �?)?�E�?8            �W@������������������������       ����[���?             B@������������������������       �~D'�$H�?#             M@                           �?�U��?           �z@������������������������       ��9��?o            �d@������������������������       �ib$�[�?�             p@                           @Vo����?I            �\@                            �?p��%��?            �F@������������������������       �      �?	             0@������������������������       �K�]l���?             =@                          �?@*�c����?.            @Q@������������������������       ��q�q�?             B@������������������������       �f��S�?            �@@       +                    @�#�%ܕ�?~           |�@       &                   �4@�8a$M��?           �z@        #                   �1@,Źo��?y            �h@!       "                    @S��-fe�?.            �S@������������������������       ��~_� �?%            �N@������������������������       ������H�?	             2@$       %                    @贁N��?K             ^@������������������������       � ����v�?'            @P@������������������������       �����n��?$            �K@'       *                    @�/�v�?�            �l@(       )                   �6@/sxQ�X�?�             k@������������������������       ��Fc58��?(            �N@������������������������       �KE���?d            `c@������������������������       ��	j*D�?             *@,       3                    �?�9m9Vh�?n           ̕@-       0                   �2@PI$K�?�           p�@.       /                    @� /XR��?�            �m@������������������������       �pp�zSy�?}            @f@������������������������       �|�j�Y�?%             N@1       2                   �:@I�$I��?            |@������������������������       ��Qڛ�?�             y@������������������������       ���8��x�?             H@4       7                   �3@�3:�@�?�           (�@5       6                     �?'έ���?�            �p@������������������������       �>��CZ�?l            �f@������������������������       ���}�?=            �V@8       9                   �5@�f�_.��?           `{@������������������������       ���w���?c            �c@������������������������       �e�� ���?�            �q@;       T                    @���+��?�           ��@<       I                   �7@bT�����?&           ��@=       D                   �6@�(
���?w           ��@>       A                    �?��$�x��?T           �@?       @                    �?��bNP�?�            �p@������������������������       �"��/g�?P            �_@������������������������       �3��|-��?P            `a@B       C                    �?�VR�s&�?�            �q@������������������������       ��)x9o�?C             \@������������������������       �������?q             e@E       H                    �?$���~��?#             I@F       G                    @A��?�?             ;@������������������������       �     ��?             0@������������������������       ����k���?             &@������������������������       ��^|�!�?             7@J       O                    @��yrkd�?�            �o@K       N                   @@@��'�s?�?�            `j@L       M                    �?i@nkw�?�            �h@������������������������       ��%7)��?o             e@������������������������       ��q�q�?             >@������������������������       �3�E��?
             *@P       S                   �;@�J����?             F@Q       R                    @j*D>�?             :@������������������������       ����X�?             ,@������������������������       �9��8���?	             (@������������������������       �n�����?             2@U       `                    @�C��K�?�            pq@V       [                    �?�����?             g@W       Z                    �?��v'���?7            �T@X       Y                   �8@Vx>y���?,            @P@������������������������       �p�j���?            �C@������������������������       �D>�Q�?             :@������������������������       ����Hx�?             2@\       ]                   �3@�Y�b�?H            @Y@������������������������       �Z�eY�e�?             5@^       _                   �9@���(\��?8             T@������������������������       ������?)            �L@������������������������       �/�6�G��?             7@a       f                    @����k��?8            �W@b       c                   �1@��7��d�?             I@������������������������       ��]�`��?	             *@d       e                    @��
6���?            �B@������������������������       �؉�؉��?             :@������������������������       ��x?r���?             &@g       j                    @c�� �?            �F@h       i                   �5@B�9(���?             ?@������������������������       ��q�q�?             (@������������������������       �"P7��?             3@������������������������       �����X�?	             ,@�t�bh�h4h7K ��h9��R�(KKkKK��h��B�?       �{@     �U@     �s@     �D@     �S@      ;@     �T@     @�@     X�@      N@      T@     �c@     ��@     �z@      .@     @P@      G@     �_@     �K@     �t@     �I@     �k@      ;@      G@      @     �L@     p|@      ~@      G@      O@      Z@     `{@     �q@       @     �B@      ;@     �V@      9@     �^@      0@     �Y@      $@      9@      @     �@@     @S@      ^@      1@      C@      H@     @a@     �Z@      �?      4@      0@      G@      4@      H@       @      :@               @              @     �C@     �N@      @      $@      5@     �O@     �@@              @              $@       @     �B@       @      9@                              @      C@     �K@      �?      @      3@     �N@      >@              @              $@              A@       @      6@                              @      @@      J@      �?      @      0@     �B@      3@              �?               @              5@       @       @                               @      0@      9@      �?      @       @      ;@      (@                              @              *@              ,@                               @      0@      ;@                       @      $@      @              �?              �?              @              @                                      @      @                      @      8@      &@               @               @               @              �?                                      @      @                      @      6@       @                               @              �?               @                                       @                                       @      @               @                              &@              �?               @                      �?      @      @      @       @       @      @                                       @      @              �?                                                      @      @       @       @       @                                       @      @                               @                      �?      @               @                      �?                                             �R@      ,@      S@      $@      7@      @      =@      C@     �M@      *@      <@      ;@     �R@     �R@      �?      1@      0@      B@      2@     �Q@      "@     @P@      @      &@              6@     �B@      F@      "@      8@      3@     �Q@     �P@      �?      *@      (@      =@      "@      ,@              ,@                              @      ,@      (@              @       @      @      &@                              @      �?      �?              "@                               @      �?      @              @      �?      @      @                              �?              *@              @                              @      *@      @                      �?      @      @                              @      �?      L@      "@     �I@      @      &@              .@      7@      @@      "@      1@      1@      P@      L@      �?      *@      (@      8@       @      =@      @      2@      @      @                      "@      1@      �?      "@      @      A@      6@               @      @      @       @      ;@      @     �@@      @       @              .@      ,@      .@       @       @      *@      >@      A@      �?      &@      @      3@      @      @      @      &@      @      (@      @      @      �?      .@      @      @       @      @      @              @      @      @      "@      @      @      @              @              �?              (@      @       @       @       @      �?               @      �?      �?              @              �?                                               @      �?       @                                      �?                                      @      @              @              �?              @       @               @       @      �?              �?      �?      �?              �?      �?      @      @      @      @      @      �?      @      �?       @      @       @      @               @      @      @      "@      �?      �?       @                              @      �?      �?               @      �?       @      @              �?       @      @      @                      @      @      @      @      �?               @      �?              @              �?              �?      �?              @     �i@     �A@     �]@      1@      5@      @      8@     �w@     �v@      =@      8@      L@     �r@     �e@      �?      1@      &@      F@      @     @P@      $@     �@@       @      @       @      @      M@     �Y@      $@       @      "@      J@     �G@              @      @      "@              B@              "@      �?      �?               @      E@     �P@      �?      @       @      *@      0@                      �?      @              "@              @                              �?      6@      =@              @              @      @                              �?              "@               @                              �?      6@      *@              @              @      @                              �?                               @                                              0@                                                                                      ;@              @      �?      �?              �?      4@     �B@      �?               @       @      &@                      �?      @              &@              @                              �?      .@      5@                       @      @      @                              �?              0@               @      �?      �?                      @      0@      �?                       @      @                      �?      @              =@      $@      8@      �?      @       @      @      0@      B@      "@      @      @     �C@      ?@              @      @      @              ;@      $@      7@              @       @      @      0@      B@      "@       @      @     �B@      =@              @      @      @              @      �?      $@               @      �?              �?      .@                      @      &@      (@                                              7@      "@      *@               @      �?      @      .@      5@      "@       @      @      :@      1@              @      @      @               @              �?      �?      �?                                              @               @       @              �?                             �a@      9@     �U@      .@      .@      �?      1@      t@      p@      3@      0@     �G@      o@     �_@      �?      *@      @     �A@      @      M@      (@      3@      @      @              @     `g@     �d@      "@      &@      5@     �]@     �M@               @       @       @      @      *@       @                                      �?      Y@      K@       @              &@     �@@      6@                                              @       @                                      �?     @U@     �B@                      $@      5@      0@                                              @                                                      .@      1@       @              �?      (@      @                                             �F@      $@      3@      @      @              @     �U@     �[@      @      &@      $@     @U@     �B@               @       @       @      @     �D@       @      2@      @      @              @     @U@     @[@      @      "@      @     @Q@      <@               @       @       @       @      @       @      �?               @              �?       @      �?      @       @      @      0@      "@                                      �?     �T@      *@     �P@      (@      $@      �?      (@     �`@     �W@      $@      @      :@     @`@     �P@      �?      &@      @      ;@       @     �@@      @       @      �?                      @      V@      H@       @      �?      @      F@      ;@              �?      �?      @              5@      @      @      �?                      @      J@      >@              �?      @      B@      1@              �?      �?      @              (@              @                                      B@      2@       @              �?       @      $@                              �?              I@      $@     �M@      &@      $@      �?      "@     �F@      G@       @      @      5@     �U@      D@      �?      $@      @      5@       @      <@              2@              @               @      :@      3@               @       @      =@       @              @      �?      @       @      6@      $@     �D@      &@      @      �?      @      3@      ;@       @       @      *@     �L@      @@      �?      @      @      1@             �]@     �A@     �X@      ,@     �@@      4@      :@     @X@     `a@      ,@      2@     �J@     `g@     �b@      *@      <@      3@     �B@      >@     �W@      :@     �Q@      $@      5@      0@      &@     �S@     @^@      &@      $@     �B@      a@     @_@      @      5@      ,@      4@      8@     �R@      "@     �G@      @      (@      @       @     �R@     �Y@       @      @      7@     �[@     @T@      �?      (@      @      ,@      @     �P@       @     �F@      @      &@       @       @     �Q@     �U@      @      @      3@      [@      T@              (@      @      *@      @      >@      �?      4@      �?      @                      K@     �E@              @      @      I@     �D@              @      @      @       @      (@      �?      @      �?      @                      6@      4@                      @      3@      =@               @      @      @       @      2@              1@                                      @@      7@              @              ?@      (@              �?               @              B@      @      9@       @       @       @       @      1@     �E@      @      @      ,@      M@     �C@              "@              @      @      ,@       @      $@       @      @      �?      �?       @      7@      @      �?      @      0@      &@              @              �?      �?      6@      @      .@              �?      �?      �?      "@      4@       @      @       @      E@      <@              @              @       @       @      �?       @              �?      @              @      0@      @              @       @      �?      �?              @      �?              @               @              �?                      �?       @      �?               @      �?      �?      �?               @                      @               @              �?                      �?      �?      �?                      �?      �?      �?                                                                                                      @                       @                                       @                      �?      �?                              @               @       @       @               @      �?                              �?      �?              4@      1@      7@      @      "@      $@      "@      @      3@      @      @      ,@      :@      F@      @      "@       @      @      3@      .@       @      5@      @      @      "@       @      @      (@       @      @      ,@      2@     �D@      @       @      @      @      2@      .@       @      4@      @      @      "@       @      @      (@       @       @      ,@      2@     �D@              @      @      @      1@      ,@       @      1@      @      @      "@      @       @      $@              �?      &@      0@      A@              @      @      @      1@      �?              @       @                       @      �?       @       @      �?      @       @      @              @              �?                              �?       @      �?                                              �?                              @       @      �?              �?      @      "@       @               @      �?      �?      �?      @      �?                       @      @      �?      �?      �?              �?      @       @      �?               @              �?      �?      @      �?                      @      @      �?              �?              �?      �?       @      �?               @              �?              @      �?                      �?                              �?                      @                                                      �?                                       @      @      �?                              �?              @      �?                      �?                      @                              @                      �?                              9@      "@      <@      @      (@      @      .@      3@      2@      @       @      0@     �I@      9@      @      @      @      1@      @      2@      @      7@      @      "@      @       @      "@      $@      @      @      *@      9@      ,@      @      @      @      *@      @       @      @      @              @       @       @      @      "@      �?      @      @      3@      @      @       @       @       @       @      @      @       @              @       @       @      @      @              @      @      0@      @      @       @       @       @       @      @               @              �?       @              @      @              @      @      @      @               @               @               @      @                       @               @                                              "@      �?      @               @               @      @              �?                                      @      @      �?               @      @                                                      $@       @      4@      @      @       @      @       @      �?       @      @       @      @      @      @      �?       @      &@      @      @              �?                                                               @      �?      �?      @                      �?       @      �?      @       @      3@      @      @       @      @       @      �?       @       @      @      @      @      @      �?      �?      @      @      @      �?      1@       @       @      �?      @       @      �?       @       @      @      @       @                      �?      �?      �?      �?      �?       @      �?      @      �?      �?                                      �?               @      @      �?               @       @      @      @      @      �?      @              @      $@       @              �?      @      :@      &@              @      �?      @              @      �?      @      �?      �?              �?       @      @              �?      @      1@      @                      �?                      @                              �?                      @                               @      �?                                                       @      �?      @      �?                      �?      @      @              �?      �?      0@      @                      �?                       @      �?              �?                              �?      @              �?      �?      &@      @                      �?                                      @                              �?       @                                      @                                                      �?      @       @               @              @       @      @                              "@      @              @              @              �?      �?      �?                               @       @       @                              "@      @              @              @                                                                       @       @                              @                                      �?              �?      �?      �?                               @                                               @      @              @               @                       @      �?               @              @              @                                      �?                              �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJm�PhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKahnh4h7K ��h9��R�(KKa��hu�B8         :                     @:�����?�	           ��@                          �2@��(�Q�?�           @�@                          �0@�Q��1��?�           ��@       	                    @�GL{"�?_            �a@                            �?     �?2             P@                           �?���c���?(             J@������������������������       ���D���?             5@������������������������       ���Y��O�?             ?@������������������������       �9��8���?
             (@
                           @� u#��?-             S@������������������������       �zv�X�?
             6@                           �?p�<�R�?#             K@������������������������       ���G���?            �B@������������������������       ��&5D�?             1@                           �?�O�n�?d           H�@                            �?���G���?�            s@                           �?E�2�AV�?�            �l@������������������������       ��3�E���?             :@������������������������       �Y�I�:��?w            �i@                           @t���`��?.            �R@������������������������       �     L�?'             P@������������������������       ���ˠ�?             &@                          �1@��bSi�?�            �q@                           @KL���?Q            `a@������������������������       ������?A            �\@������������������������       �9��8���?             8@                           �?Q�oa��?^            �a@������������������������       ��8��8��?              H@������������������������       ��η���?>            @W@       -                    �?�������?�           ,�@       &                   �<@����w!�?�           ��@        #                   �3@3o6r&��?�           �@!       "                    �?1��k���?4            �U@������������������������       ����H��?             E@������������������������       �6�h$��?            �F@$       %                    �?�GN��?X           P�@������������������������       ��9w�(��?�            �i@������������������������       ��}����?�            �s@'       *                     �?R�����?O            �\@(       )                   �@@������?B            @W@������������������������       �߂��w�?8            @S@������������������������       �     ��?
             0@+       ,                    @.�袋.�?             6@������������������������       ��8��8��?             (@������������������������       �R���Q�?             $@.       3                    �?`+��E�?           ܓ@/       2                    @@��^�l�?           0{@0       1                     �?|(��N�?�            0z@������������������������       �9�vW���?�            Pp@������������������������       �k'�ؿ��?V            �c@������������������������       �     ��?             0@4       7                    @��3�m��?            �@5       6                    �?����?{            �h@������������������������       �9��8���?             8@������������������������       ���-fX�?m            �e@8       9                    �?q=
ףS�?�            �@������������������������       �I��mk��?            �G@������������������������       ��f<��4�?z           ��@;       V                    @��1ݪ��?�           ��@<       K                   �6@���(��?�           H�@=       D                   �2@G�ї�/�?�           ��@>       A                    @��?ӟ�?�            Pr@?       @                    @����ۚ�?s             g@������������������������       ���Z�s�?\            �a@������������������������       �0,Tg��?             E@B       C                    �?�Je+���?E            @[@������������������������       �?N]l{��?            �I@������������������������       �� B�~�?&             M@E       H                    �?�m��D\�?�            y@F       G                    �?r�᮹��?m             e@������������������������       �\4仓�?>            �Y@������������������������       ���1��!�?/            �P@I       J                    �?�:Gf0Y�?�             m@������������������������       �r�qG�?U             b@������������������������       ��x?r���?4             V@L       S                   �@@��]��y�?            �y@M       P                   �7@��M�S�?�            px@N       O                    �?Q����?2            �U@������������������������       ���%����?            �@@������������������������       ��7���`�?$             K@Q       R                    @�s��:�?�             s@������������������������       �8T�r��?�            @j@������������������������       �2����*�?<            �W@T       U                    @�fG-B��?             5@������������������������       �����W�?             *@������������������������       �      �?              @W       Z                    �?�o�_,��?6            �U@X       Y                    7@*L�9��?             6@������������������������       ��T�x?r�?
             &@������������������������       �Y�����?             &@[       `                    @�A?�E~�?&            @P@\       _                   �9@��e�S�?             �L@]       ^                    �?!����?            �F@������������������������       �      �?	             0@������������������������       ����Kϟ�?             =@������������������������       ��8��8��?             (@������������������������       �      �?              @�t�bh�h4h7K ��h9��R�(KKaKK��h��B�9        |@      U@     v@      G@      W@      =@     @U@     ��@     (�@     �L@     �V@     `b@     X�@     �z@      "@     �P@     �E@     �`@     �E@     �s@      L@      m@      <@      J@      @     @P@     Pz@     �}@      D@     @P@     @W@     �{@     p@      @     �G@      8@     @T@      3@     @S@      @     �C@                              0@     @l@      d@      @      @      3@     @\@      F@              @              "@      @      0@              @                                      K@      F@                      �?      1@      @                                              @              @                                      0@      ;@                              $@      �?                                              @              @                                      $@      :@                              @      �?                                               @               @                                      @      "@                              �?      �?                                              @              �?                                      @      1@                              @                                                       @                                                      @      �?                              @                                                      "@              �?                                      C@      1@                      �?      @      @                                              @                                                      $@      �?                              @                                                       @              �?                                      <@      0@                      �?      @      @                                               @              �?                                      2@      ,@                               @                                                                                                              $@       @                      �?      �?      @                                             �N@      @     �A@                              0@     �e@      ]@      @      @      2@      X@      D@              @              "@      @      @@       @      *@                              @      ]@     @P@      �?              $@      B@      8@                                              9@       @       @                              @     @W@      I@      �?              @      6@      0@                                              @              @                                      @      @                      �?      @      @                                              4@       @      @                              @     �U@     �G@      �?              @      3@      *@                                              @              @                                      7@      .@                      @      ,@       @                                              @              @                                      6@      "@                      @      ,@      @                                              �?              �?                                      �?      @                                       @                                              =@      @      6@                              $@      L@     �I@      @      @       @      N@      0@              @              "@      @      0@      @      @                              @      =@      :@      �?      @      @      @@      @                               @      @      .@      @      @                              @      5@      5@              @      @      >@      @                                      @      �?              �?                                       @      @      �?              @       @      �?                               @              *@              .@                              @      ;@      9@      @               @      <@      &@              @              @              $@              �?                                      (@      @                      �?      @      @              @              @              @              ,@                              @      .@      3@      @              �?      5@       @                               @             �m@     �I@      h@      <@      J@      @     �H@     `h@     �s@     �A@     �M@     �R@     �t@     �j@      @      F@      8@      R@      0@      V@      1@     �V@       @      ;@      @      4@     �D@     @S@      .@      @@      ?@      [@     �R@      @      9@      *@      C@      &@      T@      ,@      U@      @      (@      �?      (@      D@     @P@      @      9@      6@     �Z@      Q@      @      7@      @      >@      @      *@       @      $@                                      $@      (@       @      @      @      $@      1@               @              �?               @              @                                      @       @       @                       @      @                                              @       @      @                                      @      @              @      @       @      &@               @              �?             �P@      (@     �R@      @      (@      �?      (@      >@     �J@      @      6@      1@     @X@     �I@      @      5@      @      =@      @     �@@      @      4@       @      @      �?      @      $@      6@      �?      *@       @     �I@      1@              @       @      @      @      A@      @      K@      @       @              "@      4@      ?@      @      "@      .@      G@      A@      @      ,@      @      6@       @       @      @      @      @      .@      @       @      �?      (@      "@      @      "@      �?      @               @       @       @      @      @      @      @      @      "@      @       @      �?      (@       @      @       @      �?      @               @       @      @       @      @      @      @       @      @      @       @      �?      &@      @      @      @      �?      @              �?       @      @       @                              �?       @                              �?      @              @                              �?              �?              �?                              @                                      �?       @      �?               @                      @      �?       @                                      @                                      �?       @                       @                       @                      �?                              �?                                                      �?                                      @      �?       @     �b@      A@     �Y@      4@      9@      @      =@     @c@     �m@      4@      ;@     �E@     �k@     @a@              3@      &@      A@      @     �D@      0@      9@      @      @      �?      @     �M@     �[@      @      &@      *@     �Q@      N@              @      �?      @      @     �D@      0@      9@      @      @              @     �M@     �[@      @      &@      *@     �P@      J@              @                      @      0@      �?      0@              @              @      B@     @R@      @       @      "@      G@      E@               @                       @      9@      .@      "@      @                       @      7@     �B@      �?      @      @      5@      $@              @                      �?                                              �?                                                      @       @                      �?      @             �Z@      2@     @S@      1@      6@       @      8@     �W@     �_@      .@      0@      >@      c@     �S@              *@      $@      ?@       @      9@      @      0@       @      *@       @      "@      0@      7@      @      @      �?      >@     �@@              @      @      @      �?      �?              @              @              @      @       @                              @                              @      �?              8@      @      *@       @      $@       @      @      (@      5@      @      @      �?      ;@     �@@              @              @      �?     �T@      ,@     �N@      .@      "@              .@     �S@     �Y@      (@      (@      =@     �^@     �F@              $@      @      8@      �?      $@              �?      @                       @      @       @      @                      @       @               @              �?              R@      ,@      N@      $@      "@              *@      R@     @Y@       @      (@      =@     �]@     �B@               @      @      7@      �?     �`@      <@     @^@      2@      D@      6@      4@      [@     �a@      1@      9@      K@     �e@     @e@      @      4@      3@     �I@      8@      _@      ;@     @Z@      1@      B@      2@      ,@     �Y@     �`@      .@      5@     �G@     @e@     �c@      @      4@      2@     �H@      8@     @S@      0@      P@      @      *@      @      @     �V@     �V@      @       @      7@      a@     �X@              @      @     �B@      @     �B@      @     �A@      �?       @              �?     �K@     �D@              @      @     �K@      A@              @       @      *@              ;@      @      *@      �?       @              �?      5@      9@               @      �?      E@      ;@              @       @      (@              ;@      @      &@      �?       @              �?      2@      (@               @      �?     �A@      .@              @       @      @                               @                                      @      *@                              @      (@                              @              $@              6@                                      A@      0@              �?      @      *@      @                              �?              @              1@                                      @      $@              �?      @       @       @                                              @              @                                      ;@      @                       @      @      @                              �?              D@      &@      =@       @      &@      @      @     �A@      I@      @      @      1@     �T@      P@              @      @      8@      @      2@              *@      �?      �?      @              9@      7@      �?      @       @      <@      A@               @       @      "@       @      (@              $@      �?      �?      @              &@      .@              �?      �?      &@      :@              �?      �?      @       @      @              @                      �?              ,@       @      �?       @      �?      1@       @              �?      �?      @              6@      &@      0@      �?      $@              @      $@      ;@      @       @      .@      K@      >@               @      @      .@      @      (@      @       @              "@              @      �?      $@      @       @      *@     �A@      4@               @      @      &@      @      $@      @       @      �?      �?              �?      "@      1@                       @      3@      $@                              @      �?     �G@      &@     �D@      ,@      7@      *@      "@      (@     �E@       @      *@      8@     �@@     �N@      @      *@      &@      (@      2@     �G@      &@     �C@      ,@      6@      $@       @      (@     �E@       @      &@      7@     �@@     �N@      @      @      &@      (@      .@      .@       @      @       @       @      @              @      1@      @      @       @      @      @                      @      �?       @      "@       @                      @      @              �?      @       @                       @       @                      �?                      @              @       @      �?      �?              @      *@       @      @       @      @      @                       @      �?       @      @@      "@     �@@      (@      ,@      @       @      @      :@      @       @      5@      :@     �K@      @      @       @      &@      *@      :@      @      5@      &@      &@      @       @      �?      3@      @      @      (@      0@      D@              @      @      &@       @      @      @      (@      �?      @      �?      @      @      @              @      "@      $@      .@      @       @      �?              @                       @              �?      @      �?                               @      �?                       @      @                      @                                      �?      @                                                                      �?      @                       @                       @                              �?                               @      �?                      �?                              �?      &@      �?      0@      �?      @      @      @      @      @       @      @      @      @      &@                      �?       @              $@              �?                              �?       @       @                      �?      @       @                                              @              �?                                      �?       @                      �?       @      �?                                              @                                              �?      �?                                      �?      �?                                              �?      �?      .@      �?      @      @      @      @      @       @      @      @       @      "@                      �?       @              �?              ,@      �?      @      @      @      @       @       @      @      @       @      @                      �?      �?              �?              ,@      �?                      @      @       @       @      @      @       @      @                      �?                                      @                                       @              �?              @      �?                              �?                      �?              @      �?                      @       @       @      �?      @       @      �?      @                                                                              @      @       @                                                      �?                              �?                      �?      �?                                               @                                      @                              �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�� ihG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKyhnh4h7K ��h9��R�(KKy��hu�Bx         >                   �2@:�N�{�?�	           ��@                           �?��l o�?�           0�@                           @�'�ם�?S           x�@                           �?@���*��?�            �l@                           @��[�?\            �b@                          �1@���<4�?-            �P@������������������������       ������w�?            �B@������������������������       �K~���?             >@	       
                     @�¾����?/            @T@������������������������       ��g:b߱�?            �F@������������������������       ��E��ӭ�?             B@                           @jU����?/            @T@                           �?����#8�?            �J@������������������������       �*L�9��?            �@@������������������������       ��Q����?             4@                          �0@      �?             <@������������������������       ��g���e�?             &@������������������������       ��?	             1@                           @1��P"`�?�            �r@                           @1�έ��?�            @m@                            �?!����?|            �g@������������������������       �@�0�!��?             A@������������������������       ��sy���?e            �c@                          �1@��&!�?            �E@������������������������       �ܶm۶m�?             <@������������������������       �l�l��?             .@                            @     ��?-             P@                           @��C�2E�?%            �H@������������������������       �xC�Ҁ��?            �@@������������������������       �     ��?             0@������������������������       �ƒ_,���?             .@        /                   �1@��®��?G           �@!       (                    �?¡g�\B�?�            �q@"       %                    �?ȥ�I M�?E            �X@#       $                   �0@v��`��?             =@������������������������       ��q�q�?             @������������������������       ��^|�!�?             7@&       '                    �?�=,E��?/            �Q@������������������������       �	�c��?             9@������������������������       �`���V�?            �F@)       ,                     �?��e�;M�?r            `g@*       +                    @=�U����?<             Y@������������������������       �r�?�b�?4            @V@������������������������       �*L�9��?             &@-       .                    @9�vW���?6            �U@������������������������       �;�yz7�?'            �P@������������������������       �lv�"��?             5@0       7                    @jxa�?��?�            �k@1       4                    @�hly+��?l            �e@2       3                    �?]Wن��?K             ]@������������������������       �5h0zF�?=            �X@������������������������       ��E��ӭ�?             2@5       6                    �?T�r
^N�?!             L@������������������������       �ֳC��2�?             F@������������������������       �VUUUUU�?
             (@8       ;                     �?�K����?$            �I@9       :                     �?�X�g�?             A@������������������������       ��Q����?             4@������������������������       ����S�r�?	             ,@<       =                    @/k��\�?             1@������������������������       ����(\��?             $@������������������������       �������?             @?       ^                   �7@��B}���?           z�@@       O                   �5@��j�N�?.           ��@A       H                    �?����&�?�           ؑ@B       E                    �?�L�����?           p}@C       D                     �?rm�< �?�            �l@������������������������       �S��d��?O             ^@������������������������       �Lh/����?A             [@F       G                    �?2.��V�?�            `n@������������������������       �����KT�?}            `j@������������������������       �     ��?             @@I       L                     @���z �?�           ��@J       K                    �?#'B�M��?'           �|@������������������������       �T�e~���?|            �g@������������������������       �M?q�?�            �p@M       N                   �4@Rf�M�K�?�             j@������������������������       ���y�b��?T             a@������������������������       ��2�tk~�?0             R@P       W                    @�m��Z�?d           ��@Q       T                     @������?�            �u@R       S                     �?</?��?�            �j@������������������������       ���B��B�?p            �f@������������������������       �     @�?             @@U       V                    @��7��?O             `@������������������������       ��������?'             Q@������������������������       ��9�pJ�?(            �N@X       [                    �?*-+��&�?�            `k@Y       Z                     �?��{a�?I             ]@������������������������       �<ݚ)�?*             R@������������������������       ��k����?             F@\       ]                    @W�A�_�?J            �Y@������������������������       �GE|A���?A            �V@������������������������       �ƵHPS!�?	             *@_       n                    �?%\,�<J�?�           P�@`       g                   �<@}��K
��?�           ��@a       d                    @�}��?           �y@b       c                     �?�H����?�            �r@������������������������       �ٝ�����?:            �V@������������������������       ��v��t�?�            @j@e       f                    @nh�)r��?G            �[@������������������������       ��!��u��?A             Y@������������������������       �{�G�z�?             $@h       k                    �?8�;���?v            �f@i       j                    �?��Eac��?%             K@������������������������       �ffffff�?             $@������������������������       ��Z=;n�?             F@l       m                   @A@     ��?Q             `@������������������������       ��*;L�?A            @Z@������������������������       ��x�W�?             7@o       v                   @A@��Uc��?e           �@p       s                    @R�+(���?X           X�@q       r                    �?�e
�S��?�            �o@������������������������       �c����?@            @Z@������������������������       ������W�?Z            �b@t       u                    @xS]$)�?�            �r@������������������������       �;Ocw���?            �i@������������������������       ������:�??             X@w       x                    @r�q��?             8@������������������������       �����X�?             ,@������������������������       ��G�z��?             $@�t�bh�h4h7K ��h9��R�(KKyKK��h��B�G       }@     @S@     �v@      @@     @T@      2@     �R@     ��@     `�@      Q@     �S@     �c@     H�@     0z@      @      P@      @@     �^@     �L@     �^@      @      R@      �?      @              @     �q@     �k@      @      @      8@     �d@     @S@              @      @      1@       @      L@      @      5@                              �?      h@     �`@       @              $@     �Q@      @@              �?              @             �@@       @      @                              �?      O@     @P@      �?              @     �@@      0@              �?              @              2@       @      @                              �?      F@     �A@                      @      2@      ,@              �?              @              "@      �?                                      �?      6@      "@                       @      @      &@              �?              @              @                                                      0@      @                       @       @      @                                              @      �?                                      �?      @       @                              @      @              �?              @              "@      �?      @                                      6@      :@                      @      *@      @                                               @      �?       @                                      $@      $@                      @      &@                                                      �?               @                                      (@      0@                               @      @                                              .@                                                      2@      >@      �?                      .@       @                                              *@                                                      1@      &@                              $@       @                                              (@                                                      "@      @                              @       @                                              �?                                                       @      @                              @                                                       @                                                      �?      3@      �?                      @                                                                                                              �?      @                              @                                                       @                                                              (@      �?                       @                                                      7@      �?      1@                                     @`@     �P@      �?              @      C@      0@                                               @      �?      1@                                     �Z@     �I@      �?              @      B@      $@                                              @      �?      .@                                     �W@      D@                      �?      ;@      @                                              �?                                                      .@      0@                              �?      �?                                              @      �?      .@                                     �S@      8@                      �?      :@      @                                              �?               @                                      *@      &@      �?               @      "@      @                                                               @                                      &@      @                       @       @      �?                                              �?                                                       @      @      �?                      �?      @                                              .@                                                      7@      0@                       @       @      @                                              @                                                      5@      &@                       @       @      @                                               @                                                      *@      $@                      �?      �?      @                                              @                                                       @      �?                      �?      �?                                                       @                                                       @      @                                                                                     �P@      @     �I@      �?      @              @     �W@     �V@       @      @      ,@      X@     �F@              @      @      &@       @      C@      �?      0@              @              @     �N@      N@      �?      @      "@     �G@      :@              @              @      @      ,@      �?      @              @              @      ,@      *@      �?       @      @      4@       @               @              @      @      @              �?                                      @      @      �?              @      "@                                       @              �?                                                      �?       @                               @                                                      @              �?                                       @       @      �?              @      @                                       @               @      �?      @              @              @      &@      "@               @      �?      &@       @               @              �?      @      @      �?                      @              @                               @              @       @                                       @      @              @               @                      &@      "@                      �?      @      @               @              �?       @      8@              (@              �?                     �G@     �G@               @      @      ;@      2@              �?              �?       @      .@               @                                      7@     �A@              �?      �?      1@      @                              �?       @      &@               @                                      4@     �@@              �?      �?      0@      @                                       @      @                                                      @       @                              �?                                      �?              "@              $@              �?                      8@      (@              �?      @      $@      .@              �?                              @              $@                                      5@      "@              �?      �?      "@       @              �?                              @                              �?                      @      @                      @      �?      @                                              <@      @     �A@      �?                       @      A@      >@      �?       @      @     �H@      3@               @      @      @       @      5@      �?     �@@      �?                              4@      3@      �?       @      @     �F@      1@                      �?      @       @      0@      �?      6@      �?                              "@      1@               @      @      5@      .@                      �?      @       @      &@      �?      6@      �?                              @      0@                      @      3@      $@                              @       @      @                                                       @      �?               @               @      @                      �?                      @              &@                                      &@       @      �?                      8@       @                                              @              $@                                      @       @      �?                      1@       @                                                              �?                                      @                                      @                                                      @       @       @                               @      ,@      &@                      �?      @       @               @       @       @              @       @                                      �?      @       @                      �?      @       @               @       @      �?               @       @                                              @      @                      �?              �?                       @      �?              @                                              �?      �?      @                              @      �?               @                               @               @                              �?      @      @                              �?                                      �?               @              �?                              �?      @                                                                                                              �?                                      �?      @                              �?                                      �?             pu@     �Q@      r@      ?@     �R@      2@      Q@     @q@     �x@      P@      R@     �`@      |@     `u@      @      M@      =@     �Z@     �H@     �m@      5@      c@      "@      B@      @     �@@     @j@     �q@      ;@      D@      Q@      r@     �f@              6@      .@     �M@      1@     �d@      "@     @U@      @      7@       @      7@      e@     �h@      $@      9@      H@      f@     �`@              $@      @      H@       @      O@      @      7@       @      ,@       @      "@      N@     @Y@      �?       @      5@      O@     �Q@              @       @      6@      @      8@       @      "@              @      �?      @      =@     �O@               @      @     �C@      =@               @              $@       @      ,@              @                              �?      0@      <@               @      @      ?@      $@                              @      �?      $@       @       @              @      �?       @      *@     �A@                      @       @      3@               @              @      �?      C@       @      ,@       @       @      �?      @      ?@      C@      �?      @      ,@      7@     �D@              @       @      (@      �?      <@      �?      (@       @      @      �?      @      =@     �@@      �?      @      ,@      3@      C@              @       @      (@      �?      $@      �?       @              �?              @       @      @              �?              @      @                                             �Y@      @      O@      @      "@              ,@      [@     �W@      "@      1@      ;@     �\@     �O@              @      @      :@      @     �S@      �?      E@      @      "@               @      V@     �R@      @      (@      ,@      R@      ?@              @      �?      .@      @      A@              &@              @              @      C@     �C@      @      @      �?     �B@      "@              @               @      �?     �F@      �?      ?@      @      @              @      I@      B@               @      *@     �A@      6@              �?      �?      *@       @      8@      @      4@                              @      4@      4@      @      @      *@     �E@      @@              �?      @      &@       @      *@       @      .@                              �?      ,@      .@      @      @      @      =@      ;@                              @       @      &@       @      @                              @      @      @      �?               @      ,@      @              �?      @      @              R@      (@     �P@      @      *@       @      $@      E@     @V@      1@      .@      4@     @\@     �G@              (@      "@      &@      "@      G@      @     �M@              "@       @      @      3@     �A@      .@      (@      (@      O@      >@              "@      @      @      "@     �@@      @     �C@              @              @      "@      .@      @      @       @     �F@      6@               @       @      @      @      ;@      @      >@              @              @      "@      .@      @      @      @     �B@      3@               @       @       @      @      @              "@                                                                      @       @      @                              �?              *@      @      4@              @       @              $@      4@      $@      @      @      1@       @              �?      @       @      @      $@      @      @               @      �?              @      .@      "@                      @      �?              �?      @              �?      @              ,@               @      �?              @      @      �?      @      @      $@      @                               @      @      :@      @       @      @      @              @      7@      K@       @      @       @     �I@      1@              @       @      @              &@       @                       @                      1@     �A@              @       @      @@      $@                               @              "@                                                      "@      <@              @              1@      @                              �?               @       @                       @                       @      @                       @      .@      @                              �?              .@      @       @      @       @              @      @      3@       @              @      3@      @              @       @      @              ,@      @      @       @                      @      @      3@       @              @      3@      @              @       @      @              �?              @      �?       @                       @                               @              �?                                             �Z@     �H@     @a@      6@     �C@      ,@     �A@     �P@     @\@     �B@      @@      P@      d@     @d@      @      B@      ,@     �G@      @@     �H@      ;@     �Q@      "@      <@      "@      1@      @     �I@      3@      7@      F@     @Q@     �R@      @      8@      (@      ;@      <@      @@      4@      J@      @      1@      @      &@      @     �C@      *@      (@      >@     �N@     @P@              (@      @      ,@      (@      7@      "@      ?@       @      ,@      @      @      @      >@      (@      $@      9@      F@     �M@              @      @      (@      @       @      @      *@              @      �?      @       @       @      @      @      @      3@      (@              �?      �?      @              .@      @      2@       @       @      @       @      �?      <@      "@      @      3@      9@     �G@              @      @       @      @      "@      &@      5@      @      @              @      @      "@      �?       @      @      1@      @              @      �?       @      @       @      @      4@      @      @              @      @      "@      �?       @      @      ,@      @              @      �?       @      @      �?      @      �?                                                                              @                                                      1@      @      2@      @      &@      @      @      �?      (@      @      &@      ,@       @      $@      @      (@      @      *@      0@      �?      @      @              @              @      �?      @       @               @      @      @              �?       @              @              @                                      �?                                               @      @                                              �?      @      @              @               @      �?      @       @               @      �?      �?              �?       @              @      0@      �?      &@      @      @      @      @              @      @      &@      @      @      @      @      &@      @      *@      (@      0@      �?      $@      @      @      @      @              @      @       @       @      @      @              &@      @      *@       @                      �?               @                               @      �?      @      @                      @              �?              @     �L@      6@      Q@      *@      &@      @      2@     �M@      O@      2@      "@      4@     �V@     �U@      �?      (@       @      4@      @     �K@      3@      P@      *@      &@      @      1@     �M@     �N@      $@      "@      4@     �V@     �T@      �?      (@       @      4@      @      7@      (@      ?@      (@      @      @      @      8@      D@      "@      @      "@      =@      @@              @       @      @      �?      *@      @      *@      @      �?               @      (@      9@                      @      0@      "@              @               @              $@      "@      2@      "@      @      @      @      (@      .@      "@      @      @      *@      7@              @       @      @      �?      @@      @     �@@      �?      @      �?      &@     �A@      5@      �?      @      &@      O@     �I@      �?      @              *@      @      8@      @      ,@      �?      @      �?      "@      =@      2@               @      @     �H@      A@              �?              @       @       @      @      3@                               @      @      @      �?       @      @      *@      1@      �?      @               @      �?       @      @      @                      �?      �?              �?       @                              @                                              �?      @       @                      �?                      �?      @                               @                                              �?               @                              �?                      @                               @                                        �t�bub��      hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�<hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKuhnh4h7K ��h9��R�(KKu��hu�B�         6                   �4@�wr����?�	           ��@                          �0@����jX�?u           ؛@                           @n-xX�?y            �g@                           @�D�+��?A            �Z@                           @���Um�?4            @V@                           �?����I��?(            �Q@������������������������       �p�u=q��?             7@������������������������       ��鿈���?            �G@	       
                    �?ԍx�V�?             3@������������������������       �x�5?,�?             "@������������������������       �                     $@                            @F��ӭ��?             2@������������������������       �և���X�?             @������������������������       �t�E]t�?             &@                           @������?8            @T@                           @"�uq�?&             I@������������������������       ��&5D�?             1@                           @t�Qe6�?            �@@������������������������       �ףp=
�?             4@������������������������       ��q-�?             *@                           �?r֛w���?             ?@������������������������       ��g���e�?             &@������������������������       �)\���(�?             4@       '                     @D*ɔĒ�?�           �@                           �3@���D��?�           T�@                            �?~XM-Q��?           @�@                           �?ƌ@�9�?�            Pu@������������������������       ��~��p�?J            �^@������������������������       �bc�N��?�            `k@                           �?_[U�r�?:           0@������������������������       �JG��S��?!             K@������������������������       ���o���?           �{@!       $                    @��T~K��?�            �p@"       #                    @Z� X��?k            @c@������������������������       �	Y���|�?6            �S@������������������������       �:W��S��?5             S@%       &                     �?&(v���?J            �\@������������������������       �x�	8��?4            �T@������������������������       �     ��?             @@(       /                    �?�,1:�?;           P~@)       ,                    �?���(�?b            �c@*       +                    @�}</*��?1            @S@������������������������       �AW/���?"            �H@������������������������       �Y�Cc�?             <@-       .                    �?4]�I��?1            �T@������������������������       ��1G����?             *@������������������������       �5 �=s�?+            @Q@0       3                    �?$%�7�?�            `t@1       2                    �?(���F��?            �g@������������������������       ��5�膫�?-            @Q@������������������������       �1u��A��?R             ^@4       5                   �3@�ѷ���?Z             a@������������������������       �N贁N�?N             ^@������������������������       ��ѳ�w�?             1@7       V                    �?H�1�7�?R           ��@8       G                    �?Z:~8|�?�           |�@9       @                    �?��C��?           0y@:       =                   �6@     b�?T             `@;       <                     �?�q�q�?             B@������������������������       �<ݚ�?             2@������������������������       ������H�?             2@>       ?                   �:@���^|�?<             W@������������������������       �ʵ�:"�?            �E@������������������������       �R|�6_c�?            �H@A       D                    @�`��K��?�            0q@B       C                    �?v��:ө�?f            �c@������������������������       ��m��?6            �U@������������������������       ��z�G��?0            �Q@E       F                   �>@~qZ�!�?K            �]@������������������������       ��HPS!��?A             Z@������������������������       �؂-؂-�?
             .@H       O                   �=@e��"���?�           `�@I       L                    @j`��RB�?g           ��@J       K                    �?�E��F��?�            �m@������������������������       ��n����?U            �^@������������������������       ������?M            @]@M       N                     @`[>��@�?�            �r@������������������������       �9R�U>�?w            �e@������������������������       ��N	����?N             `@P       S                   �>@��Kz�?C            �[@Q       R                    @�Cc}h��?             <@������������������������       �     @�?             0@������������������������       ��q�q�?             (@T       U                   @@@�h�T�?1            �T@������������������������       �     ��?             @@������������������������       ��>W[���?             I@W       f                    �?�%����?�           А@X       _                    �?�_�;��?�             t@Y       \                   �5@��'[3�?g            �d@Z       [                     �?���%�?             J@������������������������       �4և����?             @������������������������       ��d�+H�?            �F@]       ^                     �?ZĄ�~��?I            �\@������������������������       �N<+	��?             >@������������������������       ��x�P���?3             U@`       c                    @��v���?_            �c@a       b                   �9@&���^B�?*             R@������������������������       ��w��#��?             I@������������������������       ��T�x?r�?             6@d       e                     �?�8��8��?5             U@������������������������       �R����?            �@@������������������������       �y�j�
�?             �I@g       n                    �?T�����?�           ��@h       k                     �?�$�>*�?�            �u@i       j                    @G4��"�?�            �j@������������������������       �\�CZY��?_            @b@������������������������       �٫~Q$�?%             Q@l       m                   �:@�Tkט��?U            �`@������������������������       ��Q�}e��?D             Z@������������������������       ���QN�?             ?@o       r                    @��6� �?           Py@p       q                   �6@�J��}��?�            �t@������������������������       �\,��#	�?B            �\@������������������������       �8¢���?�            �j@s       t                    @�6��K�?2            @S@������������������������       ����s�4�?)            @P@������������������������       ��������?	             (@�t�bh�h4h7K ��h9��R�(KKuKK��h��BxE       �{@     �U@     �s@     �B@      P@      7@      V@     �@     ��@     �Q@     �W@     �c@     X�@     p{@      &@     �P@      N@     �`@      M@     `n@      4@     �Z@      @      @      �?      ,@     x@     �u@      0@      8@     �L@      r@     `f@              5@      "@      G@      &@      <@              @               @                     �Q@     �H@              �?              4@      (@                                              1@              @               @                      <@     �A@              �?              &@      "@                                              0@              @                                      8@      8@              �?              &@      "@                                              0@              @                                      5@      "@              �?              $@      "@                                              @              @                                      @      @                                                                                      "@                                                      .@      @              �?              $@      "@                                                                                                      @      .@                              �?                                                                                                              @      @                              �?                                                                                                                      $@                                                                                      �?                               @                      @      &@                                                                                                                                              @      @                                                                                      �?                               @                      �?      @                                                                                      &@              �?                                     �E@      ,@                              "@      @                                               @                                                      A@      @                              @      �?                                                                                                      "@      @                              @                                                       @                                                      9@       @                              @      �?                                                                                                      2@       @                                                                                       @                                                      @                                      @      �?                                              "@              �?                                      "@      @                              @       @                                              @                                                      @                                      �?                                                      @              �?                                       @      @                               @       @                                             �j@      4@     @Y@      @      @      �?      ,@     �s@     �r@      0@      7@     �L@     �p@     �d@              5@      "@      G@      &@     �b@      0@      O@       @      �?               @     p@      k@      @      $@     �A@     `g@     �Y@              (@       @      9@      "@     @[@      .@     �I@      �?                      @     `j@     �e@      @      @      7@     �`@     @R@              @      @      3@      @     �E@      $@      2@      �?                      �?      Q@     �R@       @      @      *@      N@     �@@                       @      "@      @      8@      @      "@                              �?      .@      2@                      @      9@      .@                              @       @      3@      @      "@      �?                             �J@      L@       @      @      "@     �A@      2@                       @      @      �?     �P@      @     �@@                              @     �a@     @Y@      @              $@      R@      D@              @       @      $@      �?      0@              @                               @      @       @       @              @      @      @               @                              I@      @      =@                              @      a@     @W@      @              @     @Q@      B@              @       @      $@      �?     �D@      �?      &@      �?      �?              �?      G@      E@              @      (@     �K@      >@              @      @      @      @      :@              "@      �?                      �?      4@      ;@               @       @      9@      8@              @              @      @      (@              @                                      $@      ,@              �?      �?      5@      (@                               @      �?      ,@              @      �?                      �?      $@      *@              �?      @      @      (@              @               @       @      .@      �?       @              �?                      :@      .@              @      @      >@      @              @      @       @       @      @              �?              �?                      6@      *@              @      @      7@      �?              @      @      �?       @      $@      �?      �?                                      @       @                      �?      @      @                              �?             @P@      @     �C@      @      @      �?      @     �L@      T@      "@      *@      6@     �T@      P@              "@      �?      5@       @      A@      @      "@       @      @      �?      @      4@      7@      �?      @      @      4@      4@              @              @              ,@      �?      @              �?      �?              "@      (@      �?              �?      (@      ,@              �?              @              ,@      �?                      �?      �?              @      @      �?              �?       @       @              �?              @                              @                                      @      @                              @      @                                              4@       @      @       @      @              @      &@      &@              @      @       @      @              @                                                               @                      @                                      @                      �?                              4@       @      @       @      �?              @      @      &@              @      @      @      @              @                              ?@      �?      >@      @                      @     �B@     �L@       @      $@      1@     �O@      F@              @      �?      0@       @      ,@              8@      �?                       @      .@      <@      @      @      (@     �B@      @@               @      �?      $@       @      @              @                               @      $@      5@              �?      @      &@      @                              �?      �?      $@              2@      �?                              @      @      @       @      @      :@      :@               @      �?      "@      �?      1@      �?      @       @                      �?      6@      =@       @      @      @      :@      (@              �?              @              *@      �?      @       @                      �?      2@      =@       @      @      @      7@      (@              �?               @              @              �?                                      @                              �?      @                                      @             `i@     �P@     `j@      >@     �L@      6@     �R@      d@     �q@     �K@     �Q@     �X@     �r@     @p@      &@     �F@     �I@      V@     �G@      X@      @@      Z@      2@     �C@      1@      E@      C@     �U@     �A@     �H@     �P@     �a@     �a@      @      ;@      B@     �D@     �C@      F@      $@     �D@      @       @       @      3@      8@     �I@      @      2@      1@     �L@      M@       @      @      ,@      *@      "@      &@      �?       @              �?              @      *@      :@      @      *@      @      6@      @               @      �?      @       @      �?              @                              @      @      @              @      �?      $@      @              �?                              �?               @                              @              @                              @       @                                                               @                                      @                      @      �?      @      �?              �?                              $@      �?      @              �?              �?      @      7@      @      $@      @      (@      @              �?      �?      @       @      @      �?                                              @      .@              @       @      @      �?              �?              @      �?      @              @              �?              �?      @       @      @      @      @      "@       @                      �?              �?     �@@      "@     �@@      @      @       @      ,@      &@      9@              @      &@     �A@      J@       @      @      *@      @      @      9@      �?      6@       @      �?      �?      @      $@      &@              @      @      0@      D@      �?      @      @      @       @      3@      �?      $@       @      �?              @      @      @              �?       @      $@      2@      �?      �?              @       @      @              (@                      �?              @      @               @      @      @      6@              @      @       @               @       @      &@      @      @      �?      &@      �?      ,@               @      @      3@      (@      �?              "@       @      @      @       @      $@      @      @      �?      @      �?      ,@               @      @      3@      (@                      @       @      @       @              �?              @              @                                                              �?               @                      J@      6@     �O@      *@      ?@      .@      7@      ,@     �A@      >@      ?@      I@     �U@     �T@      @      5@      6@      <@      >@      J@      4@     �K@      @      7@       @      5@      ,@     �@@      6@      2@      B@      U@     �S@      �?      *@      .@      9@      5@      4@      "@      1@       @      $@      @      @      "@      5@      &@      @      &@     �G@      A@      �?      @       @      ,@      @      &@       @       @      �?      @      @       @       @      (@      @      @      @      8@      2@      �?      @      @      @      @      "@      @      "@      �?      @              @      @      "@       @       @      @      7@      0@              @       @      "@       @      @@      &@      C@      �?      *@      @      0@      @      (@      &@      (@      9@     �B@      F@              @      @      &@      0@      6@      @      4@              "@      �?      @      @      "@      @      @      *@      :@      2@              @      @      "@      $@      $@       @      2@      �?      @      @      $@      �?      @      @      @      (@      &@      :@                               @      @               @       @      $@       @      @       @               @       @      *@      ,@       @      @       @       @      @      @      "@               @      �?      @      �?               @                      �?       @               @       @              @      �?       @                       @      �?      @      �?               @                      �?                       @      �?              �?               @                                                                                               @                      �?               @      �?                                      @      @      @      @                       @      @      @      ,@              @       @      @      @      �?      "@                       @              @      @                      �?      @       @      @               @              @                       @                      @      @      @      �?                      �?      @      @      @              �?       @       @      @      �?      @     �Z@      A@     �Z@      (@      2@      @      @@     �^@     �h@      4@      6@      @@     @c@     �]@      @      2@      .@     �G@       @      @@      2@      :@      @      @      @      "@     �B@      U@      @      @      @     �A@      B@              @      @      @      @      5@      @      0@              �?              @      ,@     �L@       @      �?      @      5@      3@              �?              @              @              �?                              @      @      7@              �?      �?      @      �?                              @               @                                                      �?                      �?               @      �?                                              @              �?                              @      @      7@                      �?      @                                      @              ,@      @      .@              �?              �?      "@      A@       @               @      ,@      2@              �?                              @              �?                              �?              ,@      �?               @      �?      @                                              "@      @      ,@              �?                      "@      4@      �?                      *@      *@              �?                              &@      .@      $@      @       @      @      @      7@      ;@      @      @      @      ,@      1@              @      @       @      @      "@      @       @      @       @      @      @      @      @      �?              @      @      "@              @              �?               @      @      @                      @      @      @      @                      @      @       @              @                              �?              @      @       @                      �?              �?              �?      �?      @                              �?               @      $@       @                      �?      �?      0@      5@      @      @               @       @              �?      @      �?      @      �?               @                                      *@      @               @              @      @              �?                              �?      $@                              �?      �?      @      .@      @       @              @      @                      @      �?      @     �R@      0@     @T@      "@      .@      �?      7@     @U@     �\@      ,@      1@      9@     �]@     �T@      @      (@      (@      E@      @      ?@      @     �B@      @      @              @      K@     �N@      @      &@      (@      N@      C@              @      �?      (@      �?      ;@      @      3@              @              @      :@     �D@      @      @      @      A@      ;@              @      �?      @      �?      &@      @      1@              @              @      7@      :@      �?       @      �?      7@      5@              @      �?      @              0@               @                                      @      .@       @      @      @      &@      @               @              �?      �?      @      �?      2@      @      @                      <@      4@      @      @      @      :@      &@                              @              @      �?      (@      @      �?                      :@      *@      �?      �?      @      8@      @                              @                              @               @                       @      @      @      @               @      @                              �?              F@      (@      F@      @       @      �?      3@      ?@     �J@      @      @      *@     �M@     �F@      @      @      &@      >@      @      C@      (@      B@      @      �?      �?      (@      9@      G@      @      @       @      J@      B@      @      @      &@      7@       @      9@      @      @      @                       @      *@      2@              @              *@      &@               @               @              *@      @      @@      �?      �?      �?      @      (@      <@      @       @       @     �C@      9@      @      @      &@      .@       @      @               @       @      @              @      @      @      �?      �?      @      @      "@       @                      @       @      @              @              @              @      @      @      �?      �?      @      @      @       @                      @       @      �?              @       @      �?              �?       @                                               @                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ=�flhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmK{hnh4h7K ��h9��R�(KK{��hu�B�         >                    �?5ko[��?�	           ��@       !                    �?��q9�?           ��@                           �?K��S��?>           �@                            �?ʭ�bJ�?~            @i@                          �4@��ݓ���?             I@                          �2@;U��j�?             =@������������������������       �     @�?             0@������������������������       �/y0��k�?             *@	       
                   �6@�5;j��?             5@������������������������       ��(\����?             $@������������������������       ���!pc�?             &@                           �?J�w�"w�?a             c@                          �6@W��LF�?+            �R@������������������������       ������?            �I@������������������������       �r�q��?             8@                          �1@��̆��?6            @S@������������������������       �      �?              @������������������������       ���xJ���?0            @Q@                            �?*x9/��?�            @s@                           �?*f��N�?3            �S@                          �7@T�r
^N�?             <@������������������������       �F]t�E�?             &@������������������������       ��l� {�?	             1@                          �2@t$���~�?"             I@������������������������       ��q-�?             *@������������������������       �к����?            �B@                           �?����?�            �l@                          �1@r��ճC�?<             V@������������������������       �Y�����?             &@������������������������       �Ө*��?5            @S@                             �?zv�|F��?Q            �a@������������������������       ��Q��X�?             C@������������������������       ��B�����?<             Z@"       1                    �?#|�3�?�           �@#       *                    �?]����c�?           �y@$       '                     �?B>��VY�?o            �d@%       &                   �5@J�w�"w�?"            �L@������������������������       ���Ĝ�?             =@������������������������       �$I�$I��?             <@(       )                     �?fw���?M             [@������������������������       ��"��Q�?             E@������������������������       �� ����?2            �P@+       .                     �?X����?�            �n@,       -                   �<@Xǰy��?/            �P@������������������������       � Q���E�?)            �L@������������������������       ���"e���?             "@/       0                    @�C{���?o            @f@������������������������       �;�g��J�?.            �S@������������������������       �`�[9��?A            �X@2       7                   �5@z7u?�I�?�           �@3       6                    @��y�4��?�            ps@4       5                   �0@#�/t��?�            �r@������������������������       �ݾ�z�<�?             *@������������������������       �������?�            �q@������������������������       ��T�6|��?             *@8       ;                     �?R���?           �z@9       :                     �?�	3�<f�?}            @j@������������������������       ��i
��2�?P            ``@������������������������       �#����?-            �S@<       =                   �>@�J�GT��?�             k@������������������������       ����>�?p            `f@������������������������       �",4D��?            �B@?       \                    �?Lol�A��?�           ��@@       M                   �1@�}����?�           <�@A       F                   �0@.(����?�             m@B       E                    @+7���?;             W@C       D                     �?���=A�?0             S@������������������������       �      �?             0@������������������������       �f�����?(             N@������������������������       �     ��?             0@G       J                    @��NV��?_            �a@H       I                     �?�r
^N��?             <@������������������������       ���Kh/�?             2@������������������������       �      �?	             $@K       L                    @������?J             \@������������������������       ��>��R�?$            �M@������������������������       �������?&            �J@N       U                   �9@�$���?7           8�@O       R                    @�,�k88�?�           ��@P       Q                     �?�.��Q�?�           ؄@������������������������       �xM����?�            �w@������������������������       �[�|���?�            �q@S       T                    @և���X�?)             L@������������������������       ����c���?              E@������������������������       ��>4և��?	             ,@V       Y                   �=@�Rͦ$�?[            �b@W       X                    �?$v̐���?C            �[@������������������������       �/�����?             <@������������������������       �,o����?3            �T@Z       [                    �?�lO��?             C@������������������������       ��������?             (@������������������������       ���N��N�?             :@]       l                     @�MPr��?�           �@^       e                   �3@j[�p���?=           Ќ@_       b                    �?�2A6+��?�             u@`       a                    @V�k{���?J            �_@������������������������       �Am��?$            �M@������������������������       �>z��.�?&             Q@c       d                   �1@ȇrb��?�            `j@������������������������       ��qǡ�?6             X@������������������������       ��Cp]�?Q            �\@f       i                    @��U��?l           @�@g       h                   �9@��΃��?           `{@������������������������       �1�\F���?�             u@������������������������       ��J�4�?@             Y@j       k                    @�fn��?a            @b@������������������������       �<�:�k+�?U             _@������������������������       ��袋.��?             6@m       t                   �5@�w�3��?�             m@n       q                    @��;��+�?W             `@o       p                    �?����{�??            �V@������������������������       �ޒ�� w�?             E@������������������������       �r�qG�?"             H@r       s                   �1@�B�����?            �C@������������������������       �ZZZZZZ�?	             1@������������������������       �h���eP�?             6@u       x                   �9@�zB�B��?>            �Y@v       w                   �6@d�_p�<�?              K@������������������������       ��E��ӭ�?             2@������������������������       �R�n��?             B@y       z                    @`ל�<��?            �H@������������������������       ��ח���?            �B@������������������������       �r�q��?             (@�t�bh�h4h7K ��h9��R�(KK{KK��h��BI       �z@     �R@     Pu@      @@      S@     �@@      U@     Ѐ@     H�@     �N@     �T@     @c@     ��@      |@       @     @R@      M@     �a@      M@     �g@      A@      f@      .@      I@      =@     �B@     �^@     �e@      ?@     �K@     �S@     �p@      j@      @      B@     �@@     @Q@     �F@     �U@      $@     �F@      @      *@       @       @      G@     �Q@      @      *@      3@      S@     �I@      @      "@      "@      9@       @      ?@       @      &@               @              @      ;@     �A@      �?      "@      "@      <@      9@              @      @       @      @      @              @                               @      @      ,@                              $@      @                      @                       @               @                               @      @      @                              $@      @                                               @               @                                      @      @                               @      @                                                                                               @              @                               @                                                      @              @                                       @       @                                                              @                      @              �?                                       @       @                                                               @                       @               @                                              @                                                              �?                      8@       @      @               @              �?      5@      5@      �?      "@      "@      2@      6@              @      @       @      @      *@       @      @                                      ,@      &@      �?      @      @      @      @              @               @       @      @              @                                      *@      &@      �?              @       @      @              @               @              @       @                                              �?                      @              @       @                                       @      &@              �?               @              �?      @      $@              @      @      &@      1@              @      @               @      �?                                                      �?      �?                              @                                                      $@              �?               @              �?      @      "@              @      @      @      1@              @      @               @      L@       @      A@      @      &@       @      @      3@      B@       @      @      $@      H@      :@      @       @      @      7@      @      0@              @      �?                      �?      @      &@                      @      1@      @      �?                      &@              "@              �?      �?                      �?       @      �?                              @      �?                              @              �?              �?                              �?       @      �?                              @                                                       @                      �?                                                                       @      �?                              @              @              @                                      @      $@                      @      $@      @      �?                      @              �?                                                              @                       @      @                                                      @              @                                      @      @                       @      @      @      �?                      @              D@       @      =@      @      &@       @      @      ,@      9@       @      @      @      ?@      4@      @       @      @      (@      @      (@      @      (@              �?               @      $@      "@              @              1@      @      @                       @      �?      �?                                                      @      �?                              �?      �?                                              &@      @      (@              �?               @      @       @              @              0@      @      @                       @      �?      <@      @      1@      @      $@       @       @      @      0@       @      �?      @      ,@      *@               @      @      @      @       @      @      "@                               @       @      @      �?                      �?      @                               @      �?      4@       @       @      @      $@       @               @      (@      �?      �?      @      *@       @               @      @       @       @     �Y@      8@     ``@      $@     �B@      5@      =@     @S@      Z@      <@      E@      N@     �g@     �c@      @      ;@      8@      F@     �B@     �G@      @      B@              (@      �?      @     �A@     �A@      1@      $@      4@     �W@      H@              @      @      4@      (@      1@              @              @              @      6@      7@      @      @      @      G@      3@              �?      �?      @      @      @               @                                      @      @      �?      �?      @      8@      $@                               @               @                                                      @      @                      @      .@      �?                                              �?               @                                              @      �?      �?              "@      "@                               @              ,@              @              @              @      1@      1@      @      @      @      6@      "@              �?      �?       @      @      (@              �?              @              �?       @      @      @      @       @      @      @                                               @              @                              @      .@      (@      �?              �?      0@      @              �?      �?       @      @      >@      @      =@              "@      �?      �?      *@      (@      (@      @      ,@     �H@      =@              @      @      0@      "@      @      @      @              @      �?              @       @                      @      7@      @               @              @      @      @      @      @                      �?              @       @                              7@      @                              @      @                      �?              @                                                      @                               @                              :@      @      7@              @              �?      $@      $@      (@      @      &@      :@      8@               @      @      "@      @      (@       @      (@              @                       @      @      �?       @      @      .@       @              �?      �?      @      �?      ,@       @      &@               @              �?       @      @      &@      @       @      &@      0@              �?       @      @      @      L@      1@     �W@      $@      9@      4@      8@      E@     @Q@      &@      @@      D@     @W@     @[@      @      6@      4@      8@      9@     �E@       @     �D@       @      @              @      B@      C@              @      "@      M@      J@              @              "@      �?      E@       @     �D@       @      @               @      A@      C@              @      @     �L@     �G@              @              "@              @               @                                       @      @                                      �?                                              C@       @     �C@       @      @               @      @@      A@              @      @     �L@      G@              @              "@              �?                                              �?       @                               @      �?      @                                      �?      *@      .@      K@       @      5@      4@      5@      @      ?@      &@      9@      ?@     �A@     �L@      @      0@      4@      .@      8@      @      $@      B@       @       @      @      $@      @      .@      @      (@      *@      5@      6@              "@      @      (@      ,@      @      "@      5@      �?      @      @      @      �?      &@      @      @      @      *@      3@              �?      @      @      "@              �?      .@      �?      @              @      @      @      @      @      @       @      @               @      �?      @      @       @      @      2@      @      *@      .@      &@      �?      0@      @      *@      2@      ,@     �A@      @      @      .@      @      $@       @      @      1@      @      (@      *@      "@      �?      0@       @      @      1@      ,@      @@              @      $@      @      @                      �?      �?      �?       @       @                      @      @      �?              @      @      @      @              @     �m@     �D@     �d@      1@      :@      @     �G@     �y@     �y@      >@      ;@     �R@     @w@     @n@      �?     �B@      9@     �Q@      *@     @[@      .@      O@      @      @              (@      p@     �m@      $@      *@      8@     �g@     �]@              &@       @      6@      @      9@      �?      @                               @     �Y@     �L@              �?      @      B@      �?                              �?              *@              �?                                     �E@      6@              �?              (@                                                      *@              �?                                      E@      &@              �?               @                                                                                                              ,@      �?              �?                                                                      *@              �?                                      <@      $@                               @                                                                                                              �?      &@                              @                                                      (@      �?       @                               @     �M@     �A@                      @      8@      �?                              �?                                                                      @      .@                              @                                      �?                                                                      @      $@                                                                      �?                                                                              @                              @                                                      (@      �?       @                               @      J@      4@                      @      3@      �?                                               @      �?                                       @     �A@      @                              @                                                      @               @                                      1@      *@                      @      *@      �?                                              U@      ,@     �M@      @      @              $@     �c@     �f@      $@      (@      5@      c@     @]@              &@       @      5@      @     �M@      @     �H@      @      �?              $@     �a@     �c@      @      $@      3@     �^@     �Z@              @       @      2@      �?     �J@      @     �E@      @      �?              @     @`@     �b@      @      $@      1@     �[@     �Z@              @      @      1@      �?      :@       @      7@      @                      @      G@     @Z@      @      @      "@     @R@     @P@              @      @      @      �?      ;@      @      4@      �?      �?                      U@      G@       @      @       @     �B@     �D@                      �?      $@              @              @                              @      (@      @      �?               @      (@      �?                       @      �?              @              @                              @      &@      @                       @      "@      �?                              �?                               @                              @      �?       @      �?                      @                               @                      9@      @      $@       @      @                      ,@      7@      @       @       @      >@      $@               @              @       @      7@      @      @       @      @                      *@      3@       @      �?      �?      1@      @              @              @       @      @      �?      �?                                      @      &@                      �?      �?       @               @                              1@      @      @       @      @                      $@       @       @      �?              0@      @              @              @       @       @              @              @                      �?      @       @      �?      �?      *@      @              @                                                              �?                                                              $@                      �?                               @              @               @                      �?      @       @      �?      �?      @      @               @                             @`@      :@     �Y@      &@      3@      @     �A@     �c@     �e@      4@      ,@     �I@      g@      _@      �?      :@      1@     �H@      $@     @Z@      5@     �S@      @      ,@      @      ;@     �`@     �a@      1@      *@      <@     @c@      V@      �?      8@      .@     �D@       @     �D@       @      .@              �?              @      U@     �Q@      @       @      @     �K@      <@              @      @      @      @      $@              @                               @     �G@      9@               @      �?      "@      *@              @       @      �?      @      "@               @                                      1@       @               @      �?      @      @              @                      @      �?              @                               @      >@      1@                              @      @              �?       @      �?              ?@       @      $@              �?              @     �B@     �F@      @              @      G@      .@               @      �?      @              (@      @      �?                                      0@      6@                      @      7@       @                              @              3@       @      "@              �?              @      5@      7@      @              �?      7@      @               @      �?                      P@      *@     �O@      @      *@      @      6@     �I@      R@      ,@      &@      6@     �X@      N@      �?      1@      (@      B@      @     �F@      &@     �D@      @      @      @      2@     �D@     �P@      &@      $@      (@      U@     �F@      �?      (@      @      2@              C@      @      ?@      @               @      .@     �C@     @P@      �?      @      @     @Q@      @@              &@      �?      &@              @      @      $@              @       @      @       @       @      $@      @      @      .@      *@      �?      �?      @      @              3@       @      6@      �?      @              @      $@      @      @      �?      $@      .@      .@              @      @      2@      @      1@       @      *@      �?      @              @      $@      @      @      �?      @      *@      ,@              @      @      .@       @       @              "@                              �?                                      @       @      �?                              @      �?      9@      @      9@      @      @               @      6@      ?@      @      �?      7@      >@      B@               @       @       @       @      1@       @      4@      @                      @      1@      .@              �?      &@      7@      "@              �?              @      �?      ,@       @      4@       @                      @      *@      @                      @      0@      @              �?                      �?      "@       @      @       @                      @       @      �?                      @       @      @                                              @              *@                              �?      &@      @                      �?       @       @              �?                      �?      @                       @                      �?      @      "@              �?      @      @      @                              @                                                                      @       @                      @      @      @                               @              @                       @                      �?              @              �?       @      @      �?                              �?               @      @      @              @              @      @      0@      @              (@      @      ;@              �?       @      @      �?      @              @               @                      @      *@                      @       @      (@                       @      @      �?      �?                               @                      @      @                              �?      @                              �?              @              @                                      �?       @                      @      �?       @                       @       @      �?      �?      @      �?              @              @              @      @              "@      @      .@              �?               @              �?      @                      �?              �?              @      @              "@      @      "@              �?              �?                              �?               @               @                                                      @                              �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�Q�=hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKmhnh4h7K ��h9��R�(KKm��hu�B�         8                    �?�u�����?�	           ��@                           �?�$*�F6�?           �@                          �;@Y�?$���?=           �~@                          �5@w������?           �z@                           �?���h� �?�            �n@                           �?�"p�� �?K            �[@������������������������       �y�j�
�?#            �I@������������������������       �xwwwww�?(             N@	       
                     @2ǋ���?X            �`@������������������������       �}�-����?1            �S@������������������������       �I�$I�$�?'             L@                          �:@��v���?o            @f@                            �?��t�4&�?b            �c@������������������������       �.��g���?            �D@������������������������       ��V��I�?I            �\@                            �?��J��?             6@������������������������       ��������?             $@������������������������       ��8��8��?             (@                           �?�O��K��?+            @P@                          �=@�>���T�?            �A@������������������������       �r�q��?             8@������������������������       ��9����?	             &@                          �=@�q�q�?             >@������������������������       �     @�?             0@������������������������       ��r
^N��?
             ,@       )                   �4@�h���G�?�           @�@       "                   �2@�m�� �?           Py@                            �?�vHr��?�            �l@                           �?���&��?)            @P@������������������������       ���S�
�?             ?@������������������������       ������?             A@        !                    �?��]�3��?j            �d@������������������������       �-�R���?0            �R@������������������������       �����?:             W@#       &                    �?���rm�?s            �e@$       %                    �?;K��?3            �T@������������������������       ���92���?             =@������������������������       ��b-����?            �J@'       (                    @
;&����?@             W@������������������������       �q`����?6            �S@������������������������       �������?
             ,@*       1                     �?��q�݇�?�           ؇@+       .                    �?�P�B��?�             l@,       -                   �9@�ڛ�xt�?,            �S@������������������������       �颋.���?             F@������������������������       �bq�����?             A@/       0                   �?@�0�>��?Z            `b@������������������������       �e�7�
t�?T             a@������������������������       ���ˠ�?             &@2       5                   �>@IW����?J           Ѐ@3       4                    �?��āq�?$           �}@������������������������       �Ǩ�M��?r             h@������������������������       ���#��Z�?�            �q@6       7                    �?�UB���?&            �M@������������������������       ��q�q�?             (@������������������������       ����D���?            �G@9       T                    �?��r)��?�           ��@:       G                     @��WJ �?�           ��@;       B                    @��'�ǯ�?2           ��@<       ?                    @��.|�?           ��@=       >                   �2@%z��?           �z@������������������������       �����B��?b            @c@������������������������       ��	o.���?�            0q@@       A                    @�;�%��?�            �x@������������������������       �������?            �F@������������������������       �nn��M��?�            �u@C       F                    @�	�~�n�?*            @P@D       E                     �?�Cc}h�?#             L@������������������������       �     @�?
             0@������������������������       ���Q���?             D@������������������������       ��2�tk~�?             "@H       O                    @���m���?�            `m@I       L                   �5@�A�����?F            �^@J       K                   �4@�0���?.            �T@������������������������       �m}����?&            @P@������������������������       � )O��?             2@M       N                    @�G�z�?             D@������������������������       �L$e?���?             7@������������������������       �	6c����?	             1@P       Q                   �1@T�r
^��?>             \@������������������������       �VUUUUU�?             8@R       S                    @�zv��?2             V@������������������������       ��.sxQ��?             ;@������������������������       �$�ߥ��?%            �N@U       d                   �6@�N��T��?�           ��@V       ]                   �0@��L��?�           �@W       Z                     �?&bV��?0            �Q@X       Y                     �?0���p��?            �D@������������������������       � �Cc}�?             <@������������������������       �؉�؉��?             *@[       \                    @�:m���?             >@������������������������       �      �?             0@������������������������       �d}h���?
             ,@^       a                     @�mQ��?�           ��@_       `                    @������?S           (�@������������������������       �N�F��r�?�            �u@������������������������       ���Q0�x�?v            �e@b       c                    @F��d���?d            �b@������������������������       ��I��s�?O            �_@������������������������       �c�ZB>��?             9@e       l                   �@@9�C�?�            �x@f       i                    @;�;(�?�            @w@g       h                   �>@�F����?�            �p@������������������������       �6���Z��?�            �n@������������������������       �V�Lt�<�?             3@j       k                   �8@ġ���?@            �Z@������������������������       ��8��8N�?             H@������������������������       �$:9$A��?"             M@������������������������       ��a����?             7@�t�bh�h4h7K ��h9��R�(KKmKK��h��B�@       �|@     �P@     �u@     �D@     �T@      D@     @W@     ��@     ��@     �L@     @T@     �f@     x�@     �y@      &@      T@     �H@     ``@      L@     �h@      >@      e@      3@      O@      >@     �E@     �`@     `d@      ;@     �H@     �X@     @l@     �j@       @      I@      @@     �P@     �C@      U@      $@      H@      @      2@      @      (@     �B@     �L@       @      $@      ;@      P@     �K@      @       @      @      8@      $@     �Q@      @      G@      @      (@      @      @     �B@      H@      @      @      ;@      O@      H@      @      @      @      6@      @      I@       @      ;@              @       @       @      :@     �A@              @      "@      A@      8@              @       @      1@      @      2@      �?      &@               @                      *@      ,@              �?      @      ,@      1@              �?              *@       @      (@              @                                      @      &@                      @      @      @              �?               @              @      �?      @               @                      @      @              �?              $@      *@                              &@       @      @@      �?      0@              @       @       @      *@      5@               @      @      4@      @               @       @      @      �?      5@              "@                               @      @      0@                      @      $@      @                              @      �?      &@      �?      @              @       @              @      @               @       @      $@      �?               @       @                      5@      @      3@      @      @      �?      @      &@      *@      @      �?      2@      <@      8@      @      @      @      @      @      2@      @      3@      @      @      �?      @      &@      $@      @      �?      *@      5@      6@      @      @      @      @      @      @               @                               @      @       @       @                      $@      &@      �?              �?       @              ,@      @      1@      @      @      �?       @      @       @      @      �?      *@      &@      &@       @      @      @      @      @      @                              �?                              @      �?              @      @       @                                               @                              �?                               @      �?              @              �?                                              �?                                                              �?                       @      @      �?                                              *@      @       @              @      �?      @              "@       @      @               @      @               @      �?       @      @      (@      @      �?              @              �?              @               @               @      @               @                              "@      @      �?              @                               @              �?                      @                                              @                                              �?               @              �?               @                       @                              �?              �?              @      �?      @              @       @      @                       @                      �?       @      @                                      �?              @              @              �?                      �?                                      @      �?              �?               @      �?                               @      @                      �?                      �?       @             �\@      4@     @^@      0@      F@      :@      ?@     �W@     �Z@      3@     �C@     �Q@     @d@     �c@      @      E@      9@     �E@      =@     �I@             �C@      @       @               @      O@      J@      @      @      4@     @S@     �G@              $@      �?      4@      @      <@              6@      @                       @      G@      @@       @      @      "@     �G@      5@              @              "@       @      @              @                                      2@      @      �?       @      @      6@      �?                                      �?      @                                                       @      @                       @      *@                                                      �?              @                                      $@      �?      �?       @       @      "@      �?                                      �?      7@              0@      @                       @      <@      ;@      �?       @      @      9@      4@              @              "@      �?      @              @                              �?      4@      (@               @      �?      0@      @              �?              @              1@              $@      @                      �?       @      .@      �?              @      "@      ,@               @              @      �?      7@              1@               @                      0@      4@      @      @      &@      >@      :@              @      �?      &@      @      ,@               @               @                      &@      ,@      �?       @      @      *@      @              @                      @      @                               @                      @      @      �?              �?      @      @                                              "@               @                                      @      $@               @       @      @       @              @                      @      "@              "@                                      @      @       @      �?       @      1@      3@              @      �?      &@      �?       @              @                                      @      @      �?      �?       @      1@      *@              @      �?       @      �?      �?               @                                              �?      �?                              @                              @              P@      4@     �T@      (@      E@      :@      =@     �@@      K@      ,@      @@     �I@     @U@      \@      @      @@      8@      7@      7@      4@      "@      @@       @      &@       @      &@      @      $@       @       @      "@      :@      E@              ,@      @      "@      @      @      @      @               @              @              @      �?      @       @      (@      1@              @      @      @      �?      @              @               @               @              @               @       @      @      ,@              @               @              @      @       @                               @              @      �?      �?              @      @                      @      @      �?      *@      @      ;@       @      "@       @      @      @      @      �?      @      @      ,@      9@              $@       @       @       @      *@      @      ;@      �?      "@       @      @      @      @      �?      @      @      ,@      9@               @       @       @      �?                              �?              @                                              �?                               @                      �?      F@      &@      I@      $@      ?@      2@      2@      =@      F@      (@      8@      E@     �M@     �Q@      @      2@      3@      ,@      4@      E@      &@     �H@       @      2@      *@      2@      =@      E@      &@      6@     �A@     �M@     �P@              *@      ,@      *@      .@      8@      @      4@              @      �?       @      2@      4@      @      @      "@     �C@      .@              @      @      @      "@      2@       @      =@       @      ,@      (@      $@      &@      6@      @      3@      :@      4@      J@               @       @      "@      @       @              �?       @      *@      @                       @      �?       @      @              @      @      @      @      �?      @       @                              @                                                       @                                              �?                              �?       @      @      @                       @      �?       @      @              @      @      @      @              @     0p@      B@     �e@      6@      5@      $@      I@     @y@     �{@      >@      @@     �T@     �v@     �h@      @      >@      1@      P@      1@     �`@      .@     �S@      @      "@      �?      0@     �n@     �p@      $@      *@      =@      f@     �U@              "@      @      5@      @     �X@      *@     �J@      @       @              &@     �j@     �k@      @      $@      <@     �`@      O@              @      �?      *@      @     @V@      *@     �E@      @      @               @      i@      k@      @      $@      ;@     �^@      M@              @              *@       @      I@      (@      4@       @       @               @     @V@     �Z@      @       @      5@     @Q@     �@@              @              @              "@              @                              @      L@      H@              �?      @      7@      @                                             �D@      (@      0@       @       @              @     �@@      M@      @      �?      1@      G@      ;@              @              @             �C@      �?      7@      �?      @                     �[@     �[@       @       @      @     �J@      9@              �?              @       @      �?              @                                      >@      @                              @      @                                              C@      �?      2@      �?      @                     @T@      [@       @       @      @      I@      6@              �?              @       @      "@              $@              @              @      ,@      @      �?              �?      *@      @                      �?               @      "@              @              @              @      (@      @                      �?      &@      @                                       @      @              @                                                                              @      @                                              @              �?              @              @      (@      @                      �?       @      �?                                       @                      @                                       @              �?                       @                              �?                     �A@       @      :@      �?      �?      �?      @     �@@     �F@      @      @      �?      E@      8@              @       @       @              1@       @      .@      �?      �?      �?              ,@      <@       @                      =@      @              �?       @      @              *@              @                      �?              @      7@       @                      8@      @                       @      @              $@              @                      �?              @      6@       @                      0@      @                                              @                                                              �?                               @                               @      @              @       @      $@      �?      �?                       @      @                              @      @              �?                              @              @      �?      �?                       @      @                              @      �?              �?                                       @      @                                      @                                       @       @                                              2@              &@                              @      3@      1@      �?      @      �?      *@      2@               @              @               @                                                      "@       @                              @                                                      0@              &@                              @      $@      "@      �?      @      �?       @      2@               @              @              @               @                                      @      �?                              �?      @                                              $@              @                              @      @       @      �?      @      �?      @      *@               @              @             �_@      5@      X@      2@      (@      "@      A@     �c@     �e@      4@      3@      K@     �g@     �[@      @      5@      ,@     �E@      *@      V@      @      K@      "@      @      �?      .@     �`@      a@      @      &@      =@     �]@     �S@              "@      @      8@      "@      @              �?               @                      6@      4@                      �?      "@       @                              �?              @                                                       @      3@                      �?      @      @                              �?              @                                                      @      .@                      �?       @                                                      �?                                                       @      @                              �?      @                              �?               @              �?               @                      ,@      �?                              @      @                                              �?              �?                                      @                                      @      �?                                              �?                               @                      @      �?                                      @                                             @T@      @     �J@      "@      @      �?      .@     �[@     @]@      @      &@      <@     �[@     �Q@              "@      @      7@      "@      O@      @      ?@      @      @      �?      $@      Y@     @W@      @      $@      6@     �R@     �M@              @      @      1@      @      H@      @      4@              @      �?      @     @T@     �M@       @      @      &@      G@      E@              @      �?      @      @      ,@       @      &@      @                      @      3@      A@      �?      @      &@      <@      1@               @      @      &@      @      3@      �?      6@      @      �?              @      &@      8@              �?      @      B@      (@               @              @       @      1@      �?      6@      @      �?              @      @      2@              �?      @      ?@      @                              @       @       @                                                      @      @                              @      @               @                              C@      .@      E@      "@      @       @      3@      8@      C@      1@       @      9@     @Q@      @@      @      (@       @      3@      @     �@@      .@      D@      "@      @      @      1@      8@      C@      *@       @      2@     @Q@      @@       @      (@       @      3@      @      7@       @      5@       @      @      @      ,@      0@     �A@      &@       @      ,@     �J@      7@      �?       @       @       @      @      7@       @      5@       @      �?      @      ,@      .@      =@      "@       @      *@     �I@      4@      �?       @      �?       @      @                                      @                      �?      @       @              �?       @      @                      �?                      $@      @      3@      �?      �?              @       @      @       @              @      0@      "@      �?      @      @      &@      �?      @      @       @                                       @      @                      �?      *@      @      �?      �?       @       @              @      @      1@      �?      �?              @      @               @              @      @      @              @      @      @      �?      @               @                       @       @                      @              @                      �?                                �t�bub�     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�yQhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKmhnh4h7K ��h9��R�(KKm��hu�B�         2                   �2@�"-���?�	           ��@                          �0@yK&0��?�           �@                           @!
A^�?{            �h@                           �?���FJ�?r            �f@                           �?
P����?-            �Q@                           @a���?            �H@������������������������       ���>4և�?             ,@������������������������       �np�_��?            �A@	       
                    �?�Ń����?             5@������������������������       ��x?r���?             &@������������������������       �
ףp=
�?             $@                           @փW�_�?E            �[@                           �?�/ᚶ��?#            �M@������������������������       �<�O��n�?             9@������������������������       ���.Lj�?             A@                           @\�5��?"             J@������������������������       ��T�6|��?             *@������������������������       �!�;\�O�?            �C@������������������������       ��h$���?	             .@       #                    @~���?           ��@                            @B '����?�             y@                           �?��Y];�?�            `m@                           �?����p9�?]             c@������������������������       ��f�W�?(             Q@������������������������       ��J����?5             U@                           �?֋�ܓ��?5            �T@������������������������       �o�ŏ1�?!             I@������������������������       �T]���b�?            �@@                            @c4Y���?l            �d@                           �?{��?���?U            �`@������������������������       ��o���?            �E@������������������������       ��M��?8            @V@!       "                    �?�M�v��?            �A@������������������������       �      �?              @������������������������       ���e/
�?             ;@$       +                    @˵`X�?           �z@%       (                     �?�W���?�            �s@&       '                    �?
N�AB!�?4            �T@������������������������       �!��-f�?            �E@������������������������       �
ףp=
�?             D@)       *                    @��!w �?�            �l@������������������������       �V^�q�0�?y            �g@������������������������       ���[�@��?            �E@,       /                    �?�~"���?F            �\@-       .                    @*Z�����?&            �M@������������������������       ���(\���?             D@������������������������       �0\�Uo��?             3@0       1                   �1@:/����?              L@������������������������       ���J��?             6@������������������������       �(s�	U��?             A@3       N                    �?<�~���?#           ��@4       C                   �>@ �P(6�?E           ��@5       <                   �7@�[ڑ� �?            �@6       9                     �?&f7��?�           H�@7       8                    �?�갇0�?�            pt@������������������������       �d�z���?`            `a@������������������������       ��s;�b��?x            �g@:       ;                   �6@�3{���?�             v@������������������������       �̤sk���?�            �r@������������������������       �~*_�#�?#             K@=       @                   �9@��j�G�?H           ��@>       ?                    �?�rя��?�             m@������������������������       �w�qG�?4            �U@������������������������       ��WXt�?W            `b@A       B                    @N�]Ԗ�?�            `s@������������������������       �I�}s���?�            q@������������������������       ���ͽ1��?            �B@D       I                   �@@����)��?D            �W@E       H                     @��"AM�?%             J@F       G                    �?��Kh/�?             B@������������������������       ��T�x?r�?	             &@������������������������       ���e�c]�?             9@������������������������       �      �?
             0@J       M                     @���tT��?            �E@K       L                    @���+��?             5@������������������������       �ܶm۶m�?             @������������������������       ����S�r�?
             ,@������������������������       ��!pc��?             6@O       ^                   �8@\�=/9l�?�           |�@P       W                   �5@��Pa��?�           ԑ@Q       T                    @�ަ���?�           P�@R       S                    @�=���?�           �@������������������������       ���On���?b            �b@������������������������       ����3���?3           `~@U       V                   �4@Oz�?%            @S@������������������������       ��%7)��?             E@������������������������       ��/<�׿�?            �A@X       [                    �?`�`{��?           �z@Y       Z                    �?״����?�            �h@������������������������       �ʵ�:"�?6            �U@������������������������       �������?K            �[@\       ]                   �6@�2�߱#�?�            �l@������������������������       �j��"z�?9            �X@������������������������       ��?�B�?X            ``@_       f                    �?��b �?           �z@`       c                    @!���O�?U            �`@a       b                    �?]0�kz�?<            @W@������������������������       ���8��8�?             H@������������������������       ��c��R��?            �F@d       e                     �?��n=���?            �C@������������������������       �X�3�R�?             3@������������������������       �ףp=
��?             4@g       j                    @��̈́���?�            `r@h       i                     @?(?����?�            �n@������������������������       �ܰh���?y            �f@������������������������       ��噮��?$            �O@k       l                     �?��q���?              I@������������������������       ��������?             >@������������������������       �ffffff�?             4@�t�bh�h4h7K ��h9��R�(KKmKK��h��B�@       @|@     �U@      u@      ?@     �S@      ;@     @V@      �@     H�@     @R@     @W@     �c@     ��@     `{@      (@      Q@     �F@      a@     �L@     �^@      (@     �O@              @              $@     �r@     �g@      *@      &@      >@     `c@      T@              @      @      5@      @      >@              @                                      S@      H@               @       @      4@      &@                              �?              >@              @                                     �R@     �G@               @       @      1@      @                              �?              *@              @                                     �A@      $@               @              @      �?                                              @               @                                      <@      @               @              @                                                      @                                                      @       @               @                                                                       @               @                                      7@      @                              @                                                      @              �?                                      @      @                              �?      �?                                              @                                                      @       @                                      �?                                              �?              �?                                      @      @                              �?                                                      1@                                                     �C@     �B@                       @      &@      @                              �?              $@                                                      *@      :@                              @      @                                               @                                                       @      ,@                              �?                                                       @                                                      @      (@                              @      @                                              @                                                      :@      &@                       @      @                                      �?              �?                                                      $@      �?                              �?                                                      @                                                      0@      $@                       @      @                                      �?                              @                                       @      �?                              @      @                                              W@      (@     �L@              @              $@      l@     �a@      *@      "@      <@     �`@     @Q@              @      @      4@      @     �I@      @      ;@              @              @     �T@     �P@       @       @      .@      R@      @@              @      @      (@      @     �A@      @      .@              @              @      N@      C@      @      @      (@     �B@      &@                      @      �?      @      6@      @      &@              @              �?      @@      4@       @       @      &@     �A@      @                              �?       @      *@      @       @                                      7@      @              �?      @      ,@      @                                              "@              "@              @              �?      "@      ,@       @      �?       @      5@       @                              �?       @      *@              @                               @      <@      2@      @       @      �?       @      @                      @              �?      @               @                                      3@      0@                      �?      �?      @                                              @               @                               @      "@       @      @       @              �?       @                      @              �?      0@      @      (@              �?               @      6@      <@      @      @      @     �A@      5@              @              &@      �?      .@      @      @              �?               @      5@      3@      �?       @      @      @@      0@               @              @              @      �?                      �?                      @      @      �?       @       @      "@      @                              @              "@      @      @                               @      2@      *@                      �?      7@      "@               @               @              �?              @                                      �?      "@       @       @              @      @               @              @      �?                                                                       @                                      �?                              @      �?      �?              @                                      �?      @       @       @              @      @               @                             �D@      @      >@                              @     �a@      S@      @      �?      *@     �O@     �B@              �?      �?       @              @@      @      5@                              @     �Z@     �N@      @      �?      @      J@      7@              �?                              (@      @       @                               @      2@      =@                              &@      @                                              (@               @                              �?      @      0@                              @      @                                                      @                                      �?      (@      *@                               @       @                                              4@      �?      3@                               @      V@      @@      @      �?      @     �D@      2@              �?                              (@      �?      3@                              �?     �S@      9@       @      �?      @      B@      $@                                               @                                              �?      $@      @      @                      @       @              �?                              "@              "@                              �?     �B@      .@                      $@      &@      ,@                      �?       @              @              @                                      =@       @                      �?      @      @                                              @              @                                      3@      @                               @      @                                              @                                                      $@       @                      �?       @                                                       @              @                              �?       @      @                      "@      @       @                      �?       @                                                                      @       @                      @      @      @                               @               @              @                              �?      @      @                      @      �?       @                      �?      @             �t@     �R@     0q@      ?@     @R@      ;@     �S@     `n@     �x@      N@     �T@     �_@     |@     `v@      (@     �O@     �D@     �\@     �J@     �a@      A@     �a@      2@     �F@      2@     �B@      D@     �`@      ;@     �H@     @S@      g@     �g@      $@     �C@      @@     �N@      E@     �a@     �@@     �`@      .@     �C@      0@     �@@      D@      `@      4@      E@     �P@      g@      g@      @      @@      6@      K@     �A@     @W@      &@     �T@      @      4@      @      $@      @@     �S@      &@      :@      <@      ^@     @W@       @      ,@      "@      ;@      &@     �J@      @     �F@      �?       @               @      $@      =@      @      5@      &@      P@      F@              @       @      &@      @      =@      �?      0@              @               @      @      "@      �?      @      @      D@      ,@               @              �?      �?      8@       @      =@      �?       @              @      @      4@       @      0@      @      8@      >@              @       @      $@      @      D@       @      C@      @      (@      @       @      6@      I@       @      @      1@      L@     �H@       @      @      @      0@      @      A@      @      @@      @      $@      @       @      2@      B@      @      @      *@     �J@      G@              @      @      0@      @      @       @      @               @       @              @      ,@      @              @      @      @       @              @                      H@      6@      J@      "@      3@      $@      7@       @     �H@      "@      0@     �C@      P@     �V@       @      2@      *@      ;@      8@      8@      "@      8@              @      �?      ,@      @      4@      @      @      .@      ;@     �J@              @      @      (@      @      "@       @      @              �?      �?              @      $@      �?      @       @      2@      .@               @      @      @      @      .@      @      1@              @              ,@       @      $@      @       @      *@      "@      C@              @       @       @              8@      *@      <@      "@      .@      "@      "@       @      =@      @      &@      8@     �B@      C@       @      (@      @      .@      5@      4@      *@      3@      "@      .@      "@      @       @      <@      @      &@      7@      ?@      <@       @      &@      @      .@      5@      @              "@                              @              �?                      �?      @      $@              �?                               @      �?      @      @      @       @      @              @      @      @      $@              @      @      @      $@      @      @      �?      �?       @       @       @       @      @              @      @      @       @              @              @       @      @       @      �?      �?       @       @       @      �?      @              @      @      �?       @              @              �?      @      @                              �?              �?                               @      @               @              �?                              �?              �?      �?      �?       @      �?      �?      @              �?              �?                      @              �?      @      @                                                      �?                               @       @                      �?              @      @               @      �?              @      �?      @              �?              �?       @      @       @                      @      �?       @       @      @      �?              @      �?      �?                              �?       @      �?      @                              �?      �?       @      �?                      �?              �?                                      �?      �?      �?                              �?      �?                      �?              @      �?                                      �?      �?              @                                               @      �?                      �?              @              �?                              @      @                      @              �?              @     `g@      D@     �`@      *@      <@      "@      E@     `i@     pp@     �@@     �@@     �H@     �p@      e@       @      8@      "@      K@      &@      c@      1@      U@      &@      *@      @      8@     �e@      l@      &@      8@     �A@     �h@      [@       @      .@       @      A@      @     @[@      @     �F@      @      @      @      2@      _@     �a@      @      5@      7@      ^@      K@              @      �?      2@      @     �V@      @     �C@      @      @      @      &@     �]@     �`@      @      3@      7@      X@     �J@              @      �?      1@      @      *@       @      "@      �?              @      "@      6@      D@                      @      2@      1@                              $@             �S@      @      >@      @      @               @      X@     @W@      @      3@      1@     �S@      B@              @      �?      @      @      2@              @                              @      @       @      @       @              8@      �?                              �?              $@                                              �?      @       @                              2@      �?                              �?               @              @                              @      @              @       @              @                                                      F@      $@     �C@      @      @              @     �I@      U@      @      @      (@     �S@      K@       @      "@      �?      0@              3@      @      3@              @              �?     �A@      I@       @      @      @      :@      <@               @      �?       @              (@      @      @              @                      @      =@      �?              @      *@      &@                      �?                      @              *@                              �?      ?@      5@      �?      @              *@      1@               @               @              9@      @      4@      @      @              @      0@      A@       @              "@     �J@      :@       @      @              ,@               @      �?      ,@      @       @              �?      $@      "@       @              @      1@      ,@              @              $@              1@      @      @      @       @              @      @      9@                      @      B@      (@       @      @              @              A@      7@     �H@       @      .@      @      2@      <@      C@      6@      "@      ,@     �P@     �N@              "@      @      4@      @      $@      @      (@       @      @       @      @      0@      0@      &@      @      @      0@      *@              @       @      @       @      $@      @      (@              �?       @      @      @      *@      @      @      @      &@      $@              @      �?      @              @       @      "@              �?               @      @       @              �?      @      @      @              @                              @       @      @                       @      @              @      @       @      �?       @      @                      �?      @                      �?               @       @              �?      (@      @      @              �?      @      @                      �?               @                                                              &@       @      @                              @                                                      �?               @       @              �?      �?      �?      @              �?      @                              �?               @      8@      2@     �B@              (@      @      (@      (@      6@      &@      @      @      I@      H@              @      @      1@      @      3@      2@      :@               @      @      @      $@      4@      $@      @      @      F@      C@              @      @      .@      @      1@      "@      5@               @      �?      @       @      ,@       @      @      @      B@      6@              @      @      *@       @       @      "@      @                       @      @       @      @       @      @               @      0@               @               @      �?      @              &@              @              @       @       @      �?                      @      $@                               @      �?      @              @               @              @                      �?                      @      @                                      �?                      @               @              @       @       @                                      @                               @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJF�@3hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         @                    �?X������?�	           ��@       !                    �?�5� ��?           T�@                           �?y`��ƕ�?q           ��@                            �?F�?X��?�            �l@                           �?�qH|�?,            �N@                           3@fP*L��?             6@������������������������       ����!pc�?             &@������������������������       �������?             &@	       
                    @:ֈ�?            �C@������������������������       �d�ϙ�?             ;@������������������������       ��q�q�?             (@                          �1@�
�%��?r            �d@                           @<5rԹ��?             7@������������������������       �r�q��?	             (@������������������������       �2(&ޏ�?             &@                           �?O��E
�?b             b@������������������������       �o_Y�K�?%             J@������������������������       ��x�W��?=             W@                            �?���h��?�            �u@                           @�W�g��?=            �Y@                          �2@�H
����?0            �R@������������������������       �$߼�x�?	             .@������������������������       �k'(���?'            �M@                          �6@�Cc}�?             <@������������������������       �����>4�?             ,@������������������������       �������?             ,@                            �?�����?�            @n@                          �<@˲,˲,�?6             U@������������������������       �_O�N�v�?0            �R@������������������������       �|	�%���?             "@                           �8@MQ��.��?`            �c@������������������������       ���3h�?G            @]@������������������������       �+���i�?            �D@"       1                    �?F�f|E�?�           d�@#       *                    �?[��5���?           p{@$       '                     @���H8�?\             b@%       &                     �?��ym�K�?,            @Q@������������������������       ��)x9/�?             <@������������������������       �G0b���?            �D@(       )                   �:@�o�2z�?0            �R@������������������������       �P���T�?%            �N@������������������������       �����>4�?             ,@+       .                   �3@c+���?�            pr@,       -                    @�n#،�?*             Q@������������������������       �����W�?             *@������������������������       �"'�q"�?#            �K@/       0                    @�����?�            `l@������������������������       �0����??             [@������������������������       �� �*n��?N            �]@2       9                   �4@ޘ��Re�?�           �@3       6                   �0@bi0&���?�            �k@4       5                    @J���#�?             6@������������������������       �9��8���?             (@������������������������       ���Q��?             $@7       8                     @NbX9��?�             i@������������������������       �`*���Q�?9            @U@������������������������       �4�nτ{�?L            �\@:       =                    @��E���?�            @x@;       <                    �?����?�?�            �m@������������������������       �"��EA��?A            �Y@������������������������       �C4%��?\             a@>       ?                     �?=������?^            �b@������������������������       �[$��m�?             J@������������������������       �͐�Jƈ�?@            @X@A       ^                   �2@���O��?�           �@B       O                     �?榙�R��?�           ��@C       J                    @NbX9��?~             i@D       G                    �?���.�?[            �a@E       F                   �1@Vp���<�?+            @P@������������������������       �Z������?            �F@������������������������       ��(\����?             4@H       I                    @      �?0             S@������������������������       �o��UbQ�?#            �J@������������������������       ��a����?             7@K       L                   �0@F~��;��?#            �M@������������������������       ��(\����?             4@M       N                    �?�(�Tw��?            �C@������������������������       ����!pc�?             6@������������������������       �{�/��>�?
             1@P       W                   �0@c�"���?1           �~@Q       T                    �?�РX4��?M            �`@R       S                    @� �9��?            �I@������������������������       ��n���?             2@������������������������       �z;Cb���?            �@@U       V                     �?��¦��?2            �T@������������������������       �ښØ}��?            �A@������������������������       �`㖪@��?            �G@X       [                    @]�=���?�            �v@Y       Z                     @��exi��?�             o@������������������������       �"���X��?s            �f@������������������������       ��paRC4�?+             Q@\       ]                    @w��7 �?F            @\@������������������������       �3�c	O�?            �G@������������������������       ���]1�[�?*            �P@_       n                   �:@ģn��v�?�           ��@`       g                     @S��5�?X           ,�@a       d                    @"T���?�           �@b       c                    @�����?{           �@������������������������       �醫���?c           @�@������������������������       �������?           P{@e       f                    @pS�sG�?5            @W@������������������������       ������Y�?'            �Q@������������������������       �H��	,�?             7@h       k                    @���^��?�            q@i       j                    �?�B�����?a            �c@������������������������       ��y��T�?-            @R@������������������������       �gݪzcS�?4            �T@l       m                    �?SX�W��?G            @]@������������������������       ���=��?%            �O@������������������������       �uk~X��?"             K@o       t                    @�VW�?�            @n@p       s                   @A@�� ��?}             i@q       r                    @��ƭ�?v            �g@������������������������       ��U,�F�?<            �W@������������������������       �	����?:            �W@������������������������       �b���i��?             &@u       v                    @�ܤ��?             E@������������������������       � )O��?
             2@������������������������       ��q�q�?             8@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       �|@     �U@      u@     �C@     �N@      9@     �Z@     ��@     ��@     �K@     �T@      e@      �@     @|@      *@      O@     �F@      _@      K@      j@      C@      c@      .@     �D@      3@     �J@     �`@     @e@      >@      P@      U@     �l@     `j@      @      C@      ;@     �P@     �B@     �V@      @      I@              &@              ,@      M@     @P@      0@      .@     �B@     @Y@      M@               @      "@      6@      *@      @@       @      3@              �?              @     �B@     �C@      @       @      .@     �B@      1@              @      �?      @      @      @      �?      @                                      @      $@      �?      @      @      *@      @                      �?      �?       @       @              @                                      @      @                               @      �?                      �?                       @              @                                      @      �?                              �?      �?                                                              @                                              @                              �?                              �?                      @      �?                                              �?      @      �?      @      @      &@      @                              �?       @       @                                                               @      �?      @      @      @      @                                       @       @      �?                                              �?      �?                              @      �?                              �?              :@      �?      *@              �?              @     �@@      =@      @      @       @      8@      &@              @              @      @      �?              �?                                      @      $@      �?               @      �?                                                                                                              @       @      �?               @      �?                                                      �?              �?                                      �?       @                                                                                      9@      �?      (@              �?              @      :@      3@       @      @      @      7@      &@              @              @      @      @      �?      @                                       @      "@              @              @      @              @              �?       @      2@              @              �?              @      2@      $@       @       @      @      1@      @              �?               @      �?     �M@       @      ?@              $@              &@      5@      :@      (@      @      6@      P@     �D@              @       @      2@       @      *@       @      ,@              @               @      "@       @              �?      @      ;@      @              �?      �?      @       @      @       @      (@              @              �?      "@      @              �?      @      2@       @              �?      �?      @       @      @              �?                                      @                                       @                                       @               @       @      &@              @              �?       @      @              �?      @      0@       @              �?      �?      @       @       @               @                              �?              @                              "@      @                                                               @                                              @                              @       @                                               @                                              �?              �?                              @      �?                                              G@              1@              @              "@      (@      2@      (@      @      0@     �B@      B@              @      @      &@      @      3@              @                              @      �?      $@       @       @      @      2@      *@               @                              3@              @                                      �?      "@       @       @      @      2@      (@               @                                                                              @              �?                      �?              �?                                              ;@              (@              @              @      &@       @      $@      @      $@      3@      7@              �?      @      &@      @      ;@              "@               @              @      &@       @      @      @      "@      "@      0@                      @      @      @                      @              @                                      @              �?      $@      @              �?       @      @      @     @]@      A@     �Y@      .@      >@      3@     �C@     �R@     @Z@      ,@     �H@     �G@     @`@      c@      @      >@      2@      F@      8@      J@      (@      G@       @      &@      @      (@      C@     �K@              1@      2@     @P@     �K@       @      *@      @      6@      "@      ;@      @      &@      �?      @              �?      $@      5@              @       @      7@      0@      �?      @              ,@      �?      &@               @      �?      @              �?       @      &@               @       @      &@      @              @              @              @              @      �?      @              �?              @              �?      �?      @                                      �?              @              @              �?                       @      @              �?      �?      @      @              @               @              0@      @      @               @                       @      $@              �?              (@      (@      �?      �?              &@      �?      "@      �?      @               @                       @      $@                              $@      &@      �?                      &@      �?      @       @                                                                      �?               @      �?              �?                              9@      "@     �A@      �?      @      @      &@      <@      A@              ,@      0@      E@     �C@      �?      "@      @       @       @      @      @       @                               @      2@      1@                              0@       @                              �?                              �?                               @      @      @                                      �?                                              @      @      �?                                      (@      ,@                              0@      �?                              �?              4@      @     �@@      �?      @      @      "@      $@      1@              ,@      0@      :@     �B@      �?      "@      @      @       @      @              .@              �?      @      @      @      @              "@      @      @      6@              "@      @      @      @      ,@      @      2@      �?      @              @      @      *@              @      "@      4@      .@      �?              @              @     @P@      6@     �L@      *@      3@      0@      ;@      B@      I@      ,@      @@      =@     @P@     �X@       @      1@      &@      6@      .@     �@@      @      :@       @       @              �?      :@      6@              @      @     �D@      E@              @      �?      @       @       @              @                                      @       @                              �?                                                      @              @                                       @                                      �?                                                       @              �?                                      @       @                                                                                      9@      @      6@       @       @              �?      3@      4@              @      @      D@      E@              @      �?      @       @      $@              @              �?              �?      0@      $@               @      �?      1@      0@                              @       @      .@      @      0@       @      �?                      @      $@              @      @      7@      :@              @      �?      @              @@      2@      ?@      &@      1@      0@      :@      $@      <@      ,@      :@      8@      8@      L@       @      ,@      $@      0@      *@      >@      &@      3@      @      &@      @      @       @      9@      $@      @      (@      3@      E@              @      @      "@      @      1@      @      ,@      �?      �?      @       @      @      (@      @              @      &@      (@              �?      @      @       @      *@      @      @      @      $@      �?      @      @      *@      @      @      @       @      >@              @              @      @       @      @      (@      @      @      &@      3@       @      @      @      3@      (@      @      ,@       @      @      @      @      @                      @              @      @      @      �?                      &@      @              @              @       @      @      @       @      @       @      @      @      @      .@      �?      @      @       @      "@      @      $@       @      @      @      �?      @     @o@     �H@     �f@      8@      4@      @     �J@     �z@     Py@      9@      2@     @U@     �w@      n@      "@      8@      2@      M@      1@      P@      "@      @@                               @     @l@      c@      @       @      1@     @\@     �I@              @      @      @      @      9@      @                                      @      G@     �I@              �?      (@      <@      0@              �?      @      @      @      4@      @                                      @      B@      6@              �?      $@      8@      &@              �?              @      @      "@                                               @      6@      *@                      @      &@      @                                              @                                               @      2@      @                       @      $@                                                      @                                                      @      @                      �?      �?      @                                              &@      @                                      �?      ,@      "@              �?      @      *@      @              �?              @      @      $@                                                      "@       @              �?      @      "@      @              �?                      @      �?      @                                      �?      @      �?                              @      �?                              @              @                                                      $@      =@                       @      @      @                      @      �?               @                                                      �?      1@                                                                                      @                                                      "@      (@                       @      @      @                      @      �?              @                                                      @      @                       @      @       @                                                                                                      @      @                              �?      @                      @      �?             �C@       @      @@                              @     �f@     �Y@      @      �?      @     @U@     �A@              @               @              &@              @                                      P@     �@@                              3@      �?                              �?              @              @                                      ?@       @                              @                                                                      �?                                      "@      @                              @                                                      @               @                                      6@      @                               @                                                      @              �?                                     �@@      9@                              ,@      �?                              �?              @                                                      @      ,@                              $@                                      �?               @              �?                                      <@      &@                              @      �?                                              <@       @      <@                              @      ]@     @Q@      @      �?      @     �P@      A@              @              �?              2@       @      4@                              @     @R@     �M@      �?      �?       @      H@      1@               @              �?              &@       @      @                              @      Q@      E@      �?      �?      �?      ;@      .@               @              �?              @              *@                               @      @      1@                      �?      5@       @                                              $@               @                                     �E@      $@       @              @      2@      1@               @                              @              �?                                      7@       @      �?                      @      "@              �?                              @              @                                      4@       @      �?              @      (@       @              �?                             @g@      D@     �b@      8@      4@      @     �F@     �i@     �o@      6@      0@      Q@     �p@     �g@      "@      3@      .@      J@      ,@     �e@      8@     @^@      4@      (@      @     �B@      h@     �l@      ,@      .@     �J@     �l@     �b@      @      ,@      "@      D@      "@     �a@      2@     @Y@      (@      "@      �?      8@     `e@     �h@      $@      ,@     �D@      g@     �Z@      @      $@      @      :@      @     �^@      2@     �V@      "@      @      �?      3@     �c@      h@      @      *@      D@     @d@     �Y@      @      $@      @      :@      @     �P@      @     �K@      @      @      �?      .@     �P@     �]@      @      @      <@     @X@     �N@              @      �?      ,@      �?      L@      &@      B@      @      @              @     �V@     �R@      @      @      (@     @P@      E@      @      @      @      (@      @      4@              $@      @       @              @      .@      @      @      �?      �?      7@      @                      �?                      "@               @      @       @              @      .@      @      @      �?              0@      �?                      �?                      &@               @                                                                      �?      @       @                                              ?@      @      4@       @      @      @      *@      5@     �@@      @      �?      (@      F@      F@      @      @       @      ,@      @      .@      @      (@       @      �?      @      @      (@      5@              �?      &@      >@      0@              �?       @       @      @       @      @              @      �?      @              &@      &@              �?      @      ,@      @                       @      @      �?      @              (@      @                      @      �?      $@                      @      0@      $@              �?              @      @      0@       @       @               @               @      "@      (@      @              �?      ,@      <@      @      @              @              @              @                               @      @      @      @              �?      "@      3@               @              @              (@       @      @               @              @       @      @                              @      "@      @      �?               @              *@      0@      >@      @       @      �?       @      (@      5@       @      �?      .@     �A@      D@       @      @      @      (@      @      "@      ,@      9@      @      @      �?      @      (@      0@       @      �?      .@     �@@      =@       @      @      @      $@      @      "@      ,@      7@      @      @      �?      @      (@      .@      @      �?      .@     �@@      8@       @       @      @      $@      @      @              *@      @      @      �?      @      @      @      @              @      8@      "@       @      �?      �?      @       @      @      ,@      $@      �?                      �?      @       @      �?      �?      $@      "@      .@              �?      @      @       @                       @                                              �?       @                              @              �?                              @       @      @              @              @              @                               @      &@               @               @      �?      �?                              @              @                                                       @               @                              @       @      @                              �?              @                               @      @                               @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���'hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         8                   �4@۪�~���?�	           ��@                           �?=h\��_�?v           �@                          �1@��a��?�           �@                           @F\���?k            �e@                          �0@�G�z��?b             d@                           �?<�F-�?            �K@������������������������       �΃�\�?             =@������������������������       �h��9J�?             :@	       
                    @�
��-�?F            @Z@������������������������       ��ĕ�(�?:             U@������������������������       �^�:|z�?             5@������������������������       �      �?	             (@                           �?~��`�N�?!           `{@                            �?&�wإ��?v             f@                          �3@��-,�?$            �K@������������������������       �=���D�?            �@@������������������������       �@r��ճ�?             6@                           �?�L�� ��?R            �^@������������������������       ��&�L��?%            �M@������������������������       �87�1��?-            �O@                           @�@A5m�?�            Pp@                           @X�Qǃc�?�            �n@������������������������       �^Z�b�?u            �f@������������������������       ��#1U��?,            @P@������������������������       �����>4�?
             ,@       )                    �?�����?�           ��@       "                   �1@"YCGK��?}           ��@                            @������?�            �o@                           @R5��\�?{            `h@������������������������       ��y�.���?t             g@������������������������       ���Q��?             $@        !                    @��V�D.�?"             M@������������������������       �h�d0ܩ�?             7@������������������������       �"��\��?            �A@#       &                    @���Т��?�            v@$       %                    @�(W3	A�?�            �p@������������������������       ����Ɩ�?t            @g@������������������������       ��3_�?5             U@'       (                     �?H�)����?7            �T@������������������������       �~K$e?��?             G@������������������������       �h�m��?            �B@*       1                    �?�f�x}�?m           �@+       .                    @��nO��?�             k@,       -                   �1@
�GN��?             F@������������������������       �������?             ,@������������������������       �p^M<+�?             >@/       0                    @\_<>t�?u            �e@������������������������       �W��>���?P            �^@������������������������       � A�c�]�?%             I@2       5                     �?M=󨣰�?�            �v@3       4                   �3@>�����?|            @i@������������������������       �q`�+e�?_            �c@������������������������       �ڤ�:�^�?            �F@6       7                    @��Q���?f             d@������������������������       �      �?             @@������������������������       �     ~�?Q             `@9       X                   �:@����.�?,           ��@:       I                     �?�\����?�           ��@;       B                    �?���Y��?           |@<       ?                    @�1=�J�?v            `i@=       >                   �5@�e��v��?H            �]@������������������������       �\x ~�c�?            �@@������������������������       �σ�V#�?6            �U@@       A                   �6@�������?.             U@������������������������       �������?            �B@������������������������       �m�w6�;�?            �G@C       F                   �9@ec>����?�            �n@D       E                   �6@�P���?�             k@������������������������       ��k�Uo�??            @X@������������������������       �z>�*���?I            �]@G       H                    �?�o^M<+�?             >@������������������������       ��������?             1@������������������������       ���1G���?             *@J       Q                    �?����q��?�           ��@K       N                    @d;��K�?.           0~@L       M                     @~�Q� :�?�            w@������������������������       ��z�gU��?\            @c@������������������������       ��������?�            �j@O       P                   �9@& �����?G            �\@������������������������       �q? �h��?<            @Y@������������������������       �؉�؉��?             *@R       U                    �?���w��?�            �@S       T                   �9@
�D�#&�?�             o@������������������������       ��&�'��?�            @m@������������������������       ���2Tv�?	             .@V       W                     �?���b{@�?�            �x@������������������������       ��@N�h��?o            �f@������������������������       ���w���?�            �j@Y       h                   �>@�������?a           ��@Z       a                   �;@(cc��p�?�            �w@[       ^                    �?T�r���?X            �a@\       ]                     �?/�6�G��?             7@������������������������       �����X�?             ,@������������������������       ��2�tk~�?             "@_       `                     �?-�Մ	[�?J            @]@������������������������       �r�8�+��?+            �P@������������������������       �l	��g��?             I@b       e                     �?�]���?�            �m@c       d                   �<@�V�:Vm�?/            @R@������������������������       ���d�7��?             A@������������������������       ����%�?            �C@f       g                   �=@��$��?r            �d@������������������������       �6���q�?O            �\@������������������������       �C�����?#             J@i       p                    �?��A-�A�?h            `d@j       m                    �?*S��/��?7            �T@k       l                    @>��^�?             ?@������������������������       ���8��8�?
             (@������������������������       ����,�?
             3@n       o                    @�9J���?#             J@������������������������       �     p�?             @@������������������������       ����(\��?             4@q       t                    @�z�G��?1             T@r       s                    @��(��(�?             E@������������������������       ��@�Y��?             =@������������������������       ��q-�?             *@u       v                    �?�].��?             C@������������������������       �؉�؉��?	             *@������������������������       ��������?             9@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       P{@     @S@     `u@      =@      P@     �B@     �V@     ��@     ��@      N@      X@     �d@     p�@     �z@      0@     �P@      D@      `@     �J@      j@      ,@     �`@      @       @       @      3@     �v@     �v@      *@      :@      H@     �s@     �f@              :@      @      J@      &@      W@      @     �M@              @              @     �S@     �W@      @      .@      5@      Z@     �R@              "@      �?      >@      "@      =@              &@              �?               @     �B@      ?@      �?      �?      @      >@      2@              �?              @      �?      ;@              $@              �?               @     �A@      ?@      �?      �?      @      9@      2@              �?              @              0@              @                                      *@      &@                              @      "@                                              "@              @                                      @      $@                              �?                                                      @                                                      @      �?                               @      "@                                              &@              @              �?               @      6@      4@      �?      �?      @      6@      "@              �?              @              $@              @              �?               @      2@      "@      �?      �?      @      5@      @              �?               @              �?              �?                                      @      &@                              �?       @                              �?               @              �?                                       @                              �?      @                                              �?     �O@      @      H@              @              @     �D@      P@      @      ,@      .@     �R@     �L@               @      �?      ;@       @      <@              $@               @               @      2@      >@      @       @       @     �B@      8@              @      �?      @      @      @               @                              �?       @      @                      @      3@      @                              @      �?      @              @                                      �?      @                      @      @      @                              @              �?              @                              �?      �?       @                              *@                                              �?      5@               @               @              �?      0@      9@      @       @      @      2@      2@              @      �?      �?      @       @               @              �?                      *@      ,@                              (@       @              �?                              *@                              �?              �?      @      &@      @       @      @      @      $@               @      �?      �?      @     �A@      @      C@              @              �?      7@      A@       @      (@      @     �B@     �@@              @              7@      @      <@      @      C@              @              �?      7@      A@              &@      @     �A@      @@              @              6@      @      :@      @      6@              @              �?      0@      >@              @      @      8@      8@              @              (@      @       @              0@                                      @      @              @      �?      &@       @                              $@              @                                                                       @      �?               @      �?                              �?              ]@      "@     �R@      @       @       @      ,@     �q@     �p@      @      &@      ;@     �j@     �Z@              1@      @      6@       @      N@       @      4@      �?               @      @     �e@      d@      @      @       @     �X@      I@              @              *@              5@              @                              �?     @U@      U@               @      @      G@      @                               @              &@              @                              �?      R@     �P@               @      @      ?@      @                               @              &@              @                              �?     �P@     @P@               @      �?      =@      @                               @                                                                      @      �?                       @       @                                                      $@               @                                      *@      2@                              .@                                                       @                                                               @                              *@                                                       @               @                                      *@      $@                               @                                                     �C@       @      ,@      �?               @      @     �V@      S@      @      �?      @      J@     �G@              @              &@              <@              $@      �?               @      @      T@     �L@      @              @      A@     �A@                              &@              5@              "@      �?               @      @      G@      G@                      @      9@      3@                               @              @              �?                                      A@      &@      @                      "@      0@                              @              &@       @      @                               @      $@      3@      �?      �?              2@      (@              @                              $@       @      �?                                      @      &@      �?                      @      @               @                              �?              @                               @      @       @              �?              &@      @              �?                              L@      @      K@      @       @              @     �[@     �Z@      @       @      3@      ]@      L@              ,@      @      "@       @      9@      �?      ,@                               @      J@      I@              @       @     �B@      ,@               @      �?              �?      @              @                                      @      *@                       @      &@      @               @                                               @                                       @       @                       @                                                              @              @                                      �?      @                              &@      @               @                              6@      �?      "@                               @     �H@     �B@              @      @      :@      "@              @      �?              �?      *@              @                                     �D@      <@              @      @      1@      @                                      �?      "@      �?       @                               @       @      "@                              "@      @              @      �?                      ?@      @      D@      @       @              @     �M@     �L@      @      @      &@     �S@      E@              @      @      "@      �?      8@      @      (@      @      �?              @      B@      ?@      �?       @      @      B@      :@              @      @      @              1@      @      "@      �?                      @      A@      >@      �?      �?       @      =@      ,@              @       @      @              @              @       @      �?                       @      �?              �?      @      @      (@              �?       @      �?              @       @      <@              �?              �?      7@      :@       @       @      @     �E@      0@              �?              @      �?              �?      @                              �?      @       @               @              @       @                                              @      �?      5@              �?                      3@      8@       @              @      B@       @              �?              @      �?     �l@     �O@      j@      9@      L@     �A@      R@     �d@     �p@     �G@     �Q@     �]@      s@     @o@      0@      D@      A@      S@      E@     �e@     �D@     @b@      0@      >@      0@      J@     `c@     �l@      >@     �I@     �T@     �o@     �e@      "@      =@      ,@      I@      4@     �G@      @      K@       @      @      @      3@      :@      H@      "@      *@      8@      U@     �M@              (@       @      :@       @      8@      @      5@      �?      �?               @      (@      A@      @      @      &@     �A@      >@              @              @              @              @      �?      �?              @      $@      <@      @      �?      @      6@      3@              @              @              @                                                      @      @              �?      �?      .@       @                              �?              @              @      �?      �?              @      @      9@      @              @      @      1@              @              @              1@      @      .@                              @       @      @              @      @      *@      &@                              �?              @      �?       @                               @              @                      @       @      �?                                              $@      @      @                               @       @      �?              @              @      $@                              �?              7@      @     �@@      @      @      @      &@      ,@      ,@      @      @      *@     �H@      =@               @       @      3@       @      5@      @      @@      @       @      @      &@      ,@      *@      @      @      $@     �G@      2@              @      �?      0@      �?      $@      �?      &@      @              @      @      @      $@      �?      �?      @      "@      &@                      �?      *@              &@       @      5@               @      �?      @      "@      @      @      @      @      C@      @              @              @      �?       @              �?               @                              �?                      @       @      &@              @      �?      @      �?       @              �?               @                              �?                                      @              �?      �?      @      �?                                                                                              @       @      @               @                             �_@      A@      W@       @      9@      (@     �@@      `@     �f@      5@      C@     �M@     `e@      ]@      "@      1@      (@      8@      2@     �J@      .@      H@      @      0@      (@      5@      6@      K@      (@      <@      <@     �P@     �M@      @      &@      @      "@      *@     �B@      .@      C@       @      .@       @      ,@      &@     �H@      &@      3@      3@      J@      F@      @      $@      @      "@      @      6@      @      3@              @              "@      @      &@       @      0@      @      8@      0@                      �?      @      @      .@      "@      3@       @      (@       @      @      @      C@      @      @      .@      <@      <@      @      $@      @      @      @      0@              $@       @      �?      @      @      &@      @      �?      "@      "@      .@      .@      �?      �?                      @      0@              $@      �?      �?      @      @      &@      @      �?      @      "@      &@      .@              �?                      @                              �?                      �?                               @              @              �?                              @     �R@      3@      F@      @      "@              (@     �Z@      `@      "@      $@      ?@      Z@     �L@      @      @      @      .@      @      ?@      @      1@       @      @              @     �@@      R@               @      *@     �A@      3@               @      @      @      �?      >@      @      (@       @       @              @      >@      R@               @      "@      A@      3@               @      @      @      �?      �?              @              �?                      @                              @      �?                                                     �E@      (@      ;@       @      @              @     �R@      L@      "@       @      2@     @Q@      C@      @      @      @      &@      @      :@      @      "@              @               @      =@     �D@      @       @      $@      7@      .@              @       @      �?              1@      "@      2@       @      @              @     �F@      .@      @               @      G@      7@      @      �?      �?      $@      @     �K@      6@     �O@      "@      :@      3@      4@      (@     �A@      1@      3@     �A@     �H@     �R@      @      &@      4@      :@      6@      I@      5@      B@      @      3@      "@      0@      &@      :@      $@      ,@      .@     �@@      L@               @      *@      6@      1@      .@      $@      (@              @      �?      @      @      $@      @      @      "@      $@     �@@              @      @      @       @      @       @                      �?                       @       @                      �?      @      @                      @       @      �?      @       @                      �?                               @                              @                              @                                                                               @                              �?              @                               @      �?      (@       @      (@               @      �?      @      @       @      @      @       @      @      >@              @      �?      @      �?      @      �?      $@              �?               @      @      @      @      @      @      @      ,@              @              @              @      @       @              �?      �?      @              @                      @      @      0@                      �?              �?     �A@      &@      8@      @      0@       @      &@      @      0@      @      $@      @      7@      7@              @      "@      0@      .@      *@      �?      @              @       @      �?      �?      @              @      �?      (@      "@                       @      �?      @      @               @              �?              �?              �?                              "@      @                      @              @      $@      �?      @              @       @              �?       @              @      �?      @      @                       @      �?      �?      6@      $@      3@      @      "@      @      $@      @      *@      @      @      @      &@      ,@              @      �?      .@      "@      1@      @      (@      @      @      @      $@       @      &@      @      @       @      @       @               @      �?      "@      "@      @      @      @              @       @              �?       @       @      @      @      @      @              �?              @              @      �?      ;@      @      @      $@      @      �?      "@      @      @      4@      0@      3@      @      @      @      @      @      @      �?      &@      @      @      @      @              @              @      &@      @      @      @      �?      @      @      @       @      �?      @              @               @              @              @              @      �?      �?              �?      �?       @      �?      �?                                                      �?              @              @                                      �?       @      �?              @              @               @               @                                      �?      �?              �?                      �?              @      @       @      @       @              �?               @      &@               @      @      �?      @       @      @                      @      �?       @       @                      �?               @      @               @      @      �?      @              @      �?                      @              @       @                                      @                      @                       @               @              0@      �?      �?      @              �?      @      @              "@      *@      0@               @      �?      �?                              @      �?                              �?      �?      @              @      $@      (@               @      �?                                       @      �?                              �?      �?      @              @      "@      @               @      �?                                      @                                                       @                      �?      @                                               @              &@              �?      @                      @      �?              @      @      @                              �?              �?              @                                                                       @      @      @                                              �?               @              �?      @                      @      �?              @                                              �?        �t�bub��     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�UJhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKmhnh4h7K ��h9��R�(KKm��hu�B�         0                    �?�p)��?�	           ��@                          �2@֗ƎQ��?a           ��@                            @��� MC�?F           �~@                           @7:���F�?�            �v@                           @l�����?�            0s@                           �?�
Gp�?�            @i@������������������������       �v��`��?             =@������������������������       �F{�	�Z�?r            �e@	       
                     �?L�w�Z��?F            @Z@������������������������       �X|�W|��?            �A@������������������������       �[e�Ӟ�?,            �Q@                          �1@ �/��?$            �K@                           @(C� ��?            �C@������������������������       ��������?             8@������������������������       �
ףp=
�?             .@������������������������       �      �?             0@                           @Q�(���?W            �`@                           @(iv���?C            �X@                           �?�������?5             T@������������������������       ���Q��?             4@������������������������       ��6�i��?(             N@������������������������       ��8	���?             3@������������������������       �6�d�M6�?            �@@       '                   �6@�v��K�?           <�@                            �?3��x�?�           �@                            �?��F`���?�            �l@                           @g�˹�?K            �\@������������������������       �^N��)x�?'             L@������������������������       �?��2��?$             M@                           �?�㰞j�?I            �\@������������������������       �r�q��?             B@������������������������       ���%&��?2            �S@!       $                     @�6���?	           �y@"       #                    @�dY�>��?�            �t@������������������������       �ndG�+�?M             _@������������������������       �$B`~��?�            �i@%       &                   �3@�����?8             U@������������������������       ��r��_�?             7@������������������������       �1M.��1�?(            �N@(       /                   �@@������?~           p�@)       ,                    @7#c1w��?s           ��@*       +                   �8@�����?'           �|@������������������������       ��QT�<q�?n            �e@������������������������       �Z�&Ӣ��?�            �q@-       .                    �?�M �w�?L             ]@������������������������       ����I��?             A@������������������������       ��"\��?8            �T@������������������������       �����K�?             2@1       P                    �?{2H���?C           �@2       A                     �?M�(�>�?z           Џ@3       :                    �?D9fL�?H           ��@4       7                   �9@�H
����?X            �b@5       6                    �?{sL�n�?F            �]@������������������������       �<�bj*R�?            �G@������������������������       �Lh/����?*             R@8       9                     �?��𡌢�?             =@������������������������       ����S�r�?	             ,@������������������������       �VUUUUU�?	             .@;       >                   �2@zZ u��?�             x@<       =                   �1@0�����?(            �O@������������������������       ���Kh/�?             B@������������������������       ��k���?             ;@?       @                    �?&;_���?�            0t@������������������������       �>��R	�?L             _@������������������������       �I-�a*��?|            �h@B       I                    �?~C���?2           @~@C       F                    @l����?c            @d@D       E                   �7@���4�g�?H            �\@������������������������       ��U&k{�?1            �R@������������������������       ��������?             D@G       H                    @     ��?             H@������������������������       �8�q_��?            �@@������������������������       ��X�%��?
             .@J       M                     @�w�P�?�             t@K       L                    7@     p�?             @@������������������������       ��������?             $@������������������������       �F]t�E�?
             6@N       O                   �9@��K<<�?�             r@������������������������       �o���{��?�            �k@������������������������       �9�\@��?-            @Q@Q       ^                    �?�<���j�?�           H�@R       Y                    @����\.�?�            �t@S       V                     @�w�.��?�            �n@T       U                    @@c7�K�?z            �h@������������������������       ���6��?D            �\@������������������������       �����X�?6             U@W       X                   �4@U��`�?            �G@������������������������       ��ӭ�a��?             B@������������������������       �t�E]t�?             &@Z       ]                   �7@d��c��?6            @V@[       \                     �?��Jr�?+            �P@������������������������       �2�^��"�?             A@������������������������       �     �?             @@������������������������       ����Q��?             7@_       f                     @51�5th�?�           �@`       c                    @�h��a6�?�           `�@a       b                   �5@=d��z�?d            �d@������������������������       �<�D�^��?3            �U@������������������������       �\��,<e�?1            �S@d       e                   �5@��5QK��?-           p~@������������������������       �V��,c��?�            pq@������������������������       ����3���?�             j@g       j                    @�?����?l            �f@h       i                    @r�0��D�?^            �c@������������������������       ������?<            @Y@������������������������       ��D�M��?"            �K@k       l                   �7@��k���?             ;@������������������������       ����#���?             &@������������������������       �     ��?             0@�t�bh�h4h7K ��h9��R�(KKmKK��h��B�@       0|@     �U@     0r@      E@      Q@      @@     �P@      �@     ��@     �Q@     @W@     @h@      �@     �|@      1@      M@     �B@     @`@     �L@      l@     �@@     �]@      @      7@       @      ,@     �r@     �t@      2@     �C@     �L@     �r@     �d@      @      5@      ,@     �D@      4@     �R@      @      5@                               @     �c@     �]@      @              *@     @S@      0@                              @              J@       @      "@                              �?     @`@      X@                      $@      I@      &@                              �?              C@              "@                              �?     @]@     �T@                      @     �E@      "@                              �?              (@              @                              �?     �V@     �L@                      @      8@       @                                              @              @                                       @      @                              @      @                                              @               @                              �?     �T@      J@                      @      5@      @                                              :@               @                                      ;@      :@                      @      3@      �?                              �?              @                                                      $@      *@                       @      @                                      �?              5@               @                                      1@      *@                      �?      .@      �?                                              ,@       @                                              *@      *@                      @      @       @                                              @                                                      (@      "@                      @      @      �?                                              @                                                      @      @                      �?      @      �?                                                                                                      @      @                      @       @                                                      @       @                                              �?      @                              �?      �?                                              7@      @      (@                              �?      <@      6@      @              @      ;@      @                              @              .@      @      $@                              �?      9@      (@      @              @      4@      @                               @              .@      @      @                              �?      4@      "@      @              @      2@      @                               @              @                                                      @              @              �?      @      �?                                              $@      @      @                              �?      .@      "@                       @      *@       @                               @                              @                                      @      @                               @       @                                               @               @                                      @      $@       @                      @                                      �?             �b@      <@     �X@      @      7@       @      (@     `a@     �j@      *@     �C@      F@     �k@     �b@      @      5@      ,@     �B@      4@     @T@      @     �B@      �?      *@       @      @     �Y@      `@      @      @      5@     �`@      Q@              @       @      4@      @     �A@              2@              &@       @      �?      @@      >@      �?       @      "@      H@      9@               @              @      @      6@              $@              @              �?      *@      0@      �?              @      @@       @              �?                      �?      @              $@                              �?      @      ,@                              0@      �?                                      �?      .@                              @                      @       @      �?              @      0@      @              �?                              *@               @              @       @              3@      ,@               @      @      0@      1@              �?              @      @      @               @                                      (@      @                              @      @              �?              �?              @              @              @       @              @      $@               @      @      &@      (@                              @      @      G@      @      3@      �?       @              @     �Q@     �X@      @      @      (@      U@     �E@               @       @      ,@             �C@      @      ,@      �?       @              �?     �J@     �V@      @       @      &@      O@     �@@              �?      �?      "@              (@      @      @      �?       @              �?      &@     �E@                      @      3@      0@                              @              ;@              "@                                      E@     �G@      @       @      @     �E@      1@              �?      �?      @              @              @                               @      2@       @      �?      @      �?      6@      $@              �?      �?      @              �?                                              �?      @      @               @      �?      @       @              �?                              @              @                              �?      ,@      �?      �?      �?              2@       @                      �?      @             @Q@      6@     �N@      @      $@               @      B@      U@       @      @@      7@     �V@     @T@      @      1@      (@      1@      *@      Q@      6@      N@      @       @               @      B@      U@      @      @@      6@     @V@     @T@      @      "@      (@      1@      (@      O@      4@      J@       @       @               @      9@      L@      @      5@      4@     �P@     @P@      @      @      (@      (@      &@      >@      @      2@      �?       @               @      $@     �@@      @      "@      (@      3@      1@      @       @      @      @       @      @@      1@      A@      �?      @              @      .@      7@       @      (@       @      H@      H@              @      @      "@      "@      @       @       @      �?                              &@      <@      �?      &@       @      6@      0@               @              @      �?      �?      �?      @                                      @      3@              �?               @       @                                              @      �?      @      �?                              @      "@      �?      $@       @      4@      ,@               @              @      �?      �?              �?               @                                       @              �?      �?              �?       @                      �?     @l@      K@     �e@      C@     �F@      >@     �J@     `k@      q@      J@      K@      a@     Pu@     `r@      *@     �B@      7@     @V@     �B@     �X@      =@     @Z@      5@      ;@      4@      7@     �I@     @U@      4@      C@     �S@     �a@     @c@      @      9@      .@     �I@      >@     �N@      ,@     �F@      (@      0@      @      .@      @@      F@      &@      4@      F@      S@     �Q@              5@      @      :@      .@      ?@      �?      @              @              �?       @      .@      @      @      (@      4@      <@                      @      &@              >@      �?      @                              �?       @      ,@      �?       @      "@      2@      3@                      @      @              &@              �?                                      @       @               @       @      @       @                       @      @              3@      �?      @                              �?      @      @      �?              �?      (@      1@                       @      @              �?              �?              @                              �?      @      �?      @       @      "@                              @                              �?              @                                       @      �?      @              �?                              @              �?                                                              �?      �?                       @       @                               @              >@      *@      C@      (@      *@      @      ,@      8@      =@      @      1@      @@      L@      E@              5@       @      .@      .@      �?              @              �?              @      $@      &@              �?      @      5@      @                              �?      �?                       @              �?              @      @       @              �?      �?      ,@      @                              �?      �?      �?              @                                      @      "@                       @      @       @                                              =@      *@     �@@      (@      (@      @      &@      ,@      2@      @      0@      =@     �A@     �B@              5@       @      ,@      ,@      1@      $@      &@      �?      @              @       @      @      @      @      "@      4@      *@              @               @      $@      (@      @      6@      &@      @      @      @      (@      &@      @      *@      4@      .@      8@              .@       @      (@      @      C@      .@      N@      "@      &@      ,@       @      3@     �D@      "@      2@      A@      P@      U@      @      @      "@      9@      .@      4@      @      2@               @              �?      &@      @      @      @      ,@      6@      >@              �?      �?      ,@      @      ,@      @      @               @              �?      "@      @      @       @      "@      2@      8@              �?      �?      @      @       @       @      @              �?              �?       @      @      @       @       @      ,@      $@              �?                      @      @       @                      �?                      �?              �?              �?      @      ,@                      �?      @       @      @              &@                                       @      �?      �?      @      @      @      @                              @      �?      @              @                                      �?              �?      @      @       @      @                              @      �?      �?              @                                      �?      �?                               @       @                               @              2@      &@      E@      "@      "@      ,@      @       @      A@      @      (@      4@      E@      K@      @      @       @      &@      "@                      @                                       @      @                       @      @      $@                      @       @                              �?                                       @      �?                      �?      @                                       @                              @                                              @                      �?       @      $@                      @                      2@      &@      C@      "@      "@      ,@      @      @      >@      @      (@      2@     �B@      F@      @      @      @      "@      "@      1@      &@      :@      @      @      @      @      @      9@      @      @      1@     �A@     �C@               @      @      "@      �?      �?              (@      @       @      $@       @              @      �?      @      �?       @      @      @      �?       @               @     �_@      9@     �P@      1@      2@      $@      >@      e@     �g@      @@      0@     �M@      i@     �a@      @      (@       @      C@      @      :@       @      1@      @      @      @      $@      M@     @P@      &@       @      .@      F@     �G@               @      �?      @      @      0@      @      *@      @       @      @      @      H@      J@      @       @      *@     �C@      ?@              @               @      �?      *@      @       @      �?       @      @      @      G@      F@      @       @      @      =@      7@              @              �?      �?      @              @      �?       @      @      @      ;@      2@      @              @      4@      *@              @                      �?      @      @      �?                      @      �?      3@      :@               @       @      "@      $@                              �?              @              @      @                               @       @                      @      $@       @                              �?              @              @      @                               @      @                      @      $@      �?                                                                                                              �?                       @              @                              �?              $@      @      @              �?              @      $@      *@      @               @      @      0@              @      �?      @       @      $@              @                              �?      @      *@                       @      @      .@              @      �?       @      �?      @                                                      @      (@                       @      �?      @                      �?       @              @              @                              �?              �?                              @      "@              @                      �?              @                      �?              @      @              @                              �?                               @      �?     @Y@      1@      I@      (@      .@      @      4@     �[@      _@      5@      ,@      F@     �c@     @W@      @      @      @      @@      @      U@      *@     �C@      &@      "@       @      $@      W@     @X@      4@      (@     �@@     �`@      N@       @      �?      @      :@       @      1@       @      $@      �?       @       @      @      (@      >@      "@      @       @      7@      ;@                       @      "@              &@              @              �?              @      $@      9@      @                      @      ,@                       @      @              @       @      @      �?      �?       @       @       @      @      @      @       @      1@      *@                              @             �P@      &@      =@      $@      @              @      T@     �P@      &@      @      9@     @[@     �@@       @      �?      @      1@       @      D@      @      (@      @      �?              �?      P@     �C@              @      .@      P@      6@                      �?      @              ;@      @      1@      @      @              @      0@      <@      &@      �?      $@     �F@      &@       @      �?      @      &@       @      1@      @      &@      �?      @       @      $@      2@      ;@      �?       @      &@      9@     �@@      @      @              @       @      1@      @      &@      �?      @       @      @      1@      9@      �?              "@      8@      <@       @      @              @       @      &@      @      $@              �?       @      @      "@      *@      �?              @      .@      8@       @      @                      �?      @      �?      �?      �?       @              �?       @      (@                      @      "@      @                              @      �?                                      @              @      �?       @               @       @      �?      @       @                      @                                              �?                      �?       @               @       @      �?               @                                                                       @              @                                                      @                              @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJzm�HhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         :                    �?m^�O��?�	           ��@                           �?��	�?'           �@                           @�����?�           Є@                          �6@{��>��?J           �@                          �3@�E�����?�            �r@                           �?�1���?e             d@������������������������       ����#2�?0            @T@������������������������       �������?5             T@	       
                   �5@���Y��?_            `a@������������������������       ��>�آ��?A            �W@������������������������       ��
�GN�?             F@                           �?'vb'v��?�             j@                           �?�>v·��?9            �T@������������������������       �V�Lt�<�?             3@������������������������       �     @�?)             P@                           @�wb֋��?M            @_@������������������������       � ��]��?5            �T@������������������������       ��q�q�?             E@                           �?�)�{U�?l            �c@                          �6@\;U���?(             M@                            �?���3c�?            �@@������������������������       ��"w����?             3@������������������������       �������?
             ,@                           @��0�*�?             9@������������������������       �\��"e��?             2@������������������������       �����X�?             @                          �?@�~j�t��?D             Y@                          �4@c�� �?>            �V@������������������������       ��fG-B��?             5@������������������������       �5 �=s�?+            @Q@������������������������       ��G�z��?             $@        /                   �9@b���9�?q           P�@!       (                    �?2�ݡ�?�           ��@"       %                   �7@��`Α?�?�             o@#       $                    @d��h'��?�            @k@������������������������       ����d��?E            �\@������������������������       ���.
���?B            �Y@&       '                   �8@"?ӧ
��?             ?@������������������������       ��������?             4@������������������������       ���ˠ�?             &@)       ,                    �?�.����?*           �}@*       +                     �?     4�?P             `@������������������������       �5yy8,�?             ?@������������������������       ��e��=�?:            @X@-       .                     @�</s���?�            �u@������������������������       �R����?k            `f@������������������������       �z�=Ig��?o            �e@0       7                    @b�dD��?�             q@1       4                   �:@R�ڵ���?�            �n@2       3                    @m��1G��?             J@������������������������       �'a����?             3@������������������������       �mo�<~'�?            �@@5       6                   �?@G/����?�             h@������������������������       �'a����?a             c@������������������������       �%�Ѿ��?            �D@8       9                     �?���Kϟ�?             =@������������������������       ��t����?             1@������������������������       ���8��8�?             (@;       X                    �?�f�����?�           ��@<       K                     @�m���?�           |�@=       D                     �?E�ߩ�?=           (�@>       A                    @ś�G���?�           X�@?       @                    @�`�/�?`             d@������������������������       �b��@��?A            �[@������������������������       �x$(~��?             I@B       C                   �1@8"W��?-           �|@������������������������       �i���1d�?E            �Y@������������������������       �{�譫@�?�            @v@E       H                    @����sv�?�            �q@F       G                    @�/E7�5�?�            `i@������������������������       ��Jє���?s            �e@������������������������       �P*�n���?             =@I       J                    @��yǡ�?+            �S@������������������������       ���S���?#            �P@������������������������       �؉�؉��?             *@L       S                   �6@�6z��?�            @k@M       P                   �3@��$c��?e            �d@N       O                    �?�w�����?<            �W@������������������������       �Iє�?             A@������������������������       �>
ףp=�?%             N@Q       R                    @1t4]2�?)            �Q@������������������������       �-�.v!��?#            �M@������������������������       �t�E]t�?             &@T       W                   �<@�������?#             K@U       V                    @�Z=;n�?             F@������������������������       ���]�2��?             ?@������������������������       ��s�n_�?             *@������������������������       �
ףp=
�?             $@Y       h                   �:@�����?�           ��@Z       a                     @S����?m           h�@[       ^                   �5@P��� �?�           0�@\       ]                    �?�5Z-X�?R           ��@������������������������       �'{���.�?k            �d@������������������������       ����[z��?�            �v@_       `                     �?��OU���?�            �n@������������������������       �[T�D$��?5            �T@������������������������       �~*_�#�?h            @d@b       e                   �0@�V)�?~            �h@c       d                    @Lh/����?             2@������������������������       �ffffff�?             $@������������������������       �      �?              @f       g                    @ �m���?r            �f@������������������������       �     ��?O             `@������������������������       ��v*���?#            �J@i       n                    @TM�?9�?b             c@j       m                    @����?H            �Z@k       l                     �?�e|���?=            �V@������������������������       �5^�I�?             I@������������������������       ����Q��?              D@������������������������       �{�/��>�?             1@o       r                     �?�˫���?             G@p       q                    @L�9���?             6@������������������������       �؉�؉��?	             *@������������������������       ���"e���?             "@������������������������       �9��8���?             8@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       P|@     @U@     0v@      9@     �P@      ?@      S@     ��@     8�@     @R@     �V@      c@     ��@     0|@      0@     �Q@     �E@     @\@     �P@     �h@      I@     �f@      .@      D@      6@      D@     �Z@     �f@      @@     �K@      U@     `p@      j@      &@      E@      8@     �N@      J@     �T@      7@     �R@       @      *@       @      *@     �P@     �W@      @      6@      7@      \@      S@      @      &@      "@      2@      (@     �R@      3@     �N@      �?      @      �?      &@     �L@     �P@      @      1@      .@     �S@      L@              $@      @      1@      @     �F@       @      >@              @      �?      @     �K@      B@      @      @      @      N@      <@               @      �?      $@      �?      6@       @      *@                               @      E@      1@      @      �?      @      >@      2@              �?              @              0@              "@                                      0@       @      @               @      *@      (@              �?              �?              @       @      @                               @      :@      "@              �?      �?      1@      @                              @              7@              1@              @      �?       @      *@      3@              @      @      >@      $@              @      �?      @      �?      3@              "@              @              �?       @      &@              �?      @      4@       @              @              @      �?      @               @               @      �?      �?      @       @               @              $@       @                      �?                      =@      1@      ?@      �?      �?              @       @      >@       @      *@      "@      3@      <@               @      @      @      @      2@      "@      "@      �?      �?                      �?      *@               @       @      $@       @              �?               @                      @       @                                      �?      @              @              @                                      �?              2@      @      @      �?      �?                               @              @       @      @       @              �?              �?              &@       @      6@                              @      �?      1@       @      @      @      "@      4@              �?      @      @      @      "@      �?      0@                              @      �?      &@       @       @      @      @      2@              �?       @      @      @       @      @      @                              @              @              @       @      @       @                       @              @      "@      @      ,@      �?      @      �?       @      $@      <@       @      @       @     �@@      4@      @      �?      @      �?      @      @      @      �?               @                      @      ,@       @       @              .@      @              �?              �?              @              �?               @                      @      $@       @       @              @      �?                                              @              �?               @                      @      @       @      �?              �?                                                                                                              @      @              �?              @      �?                                              �?      @                                                      @                              $@      @              �?              �?              �?      @                                                      @                              @      @              �?              �?                                                                                                              @       @                                              @      �?      *@      �?      @      �?       @      @      ,@              @       @      2@      ,@      @              @              @      @      �?      &@      �?       @      �?       @      @      ,@              @       @      2@      ,@                      @              @      @              @                                      @      �?              @      �?      @      �?                                                      �?      @      �?       @      �?       @              *@                      @      ,@      *@                      @              @      �?               @               @                                                                              @              �?                     �\@      ;@      [@      *@      ;@      4@      ;@     �C@     @V@      9@     �@@     �N@     �b@     �`@      @      ?@      .@     �E@      D@     �X@      7@     �S@      @      &@       @      .@     �A@     @T@      0@      ,@     �F@     �`@     @X@              1@      @     �A@      (@      C@       @      1@      �?      @      �?      @       @      ?@      @      @      0@     �L@      8@               @      @      *@      @      >@       @      .@      �?      @              @      @      ?@      @      @      .@      E@      5@               @      @      *@      @      1@      @       @              �?              �?      @      1@      @      @      "@      >@      @              @      �?       @      �?      *@      @      @      �?       @              @      �?      ,@      �?      @      @      (@      .@              �?       @      &@      @       @               @                      �?              �?                              �?      .@      @                                              @               @                                                                      �?      $@      @                                              @                                      �?              �?                                      @                                                     �N@      .@      O@      @       @      @      "@      ;@      I@      (@       @      =@     �R@     @R@              "@       @      6@      @      9@      @      ,@      �?      @      @              "@      4@      �?              @      1@      .@                              @      @      @              @                                      �?      "@      �?              �?      @      @                              �?              6@      @      &@      �?      @      @               @      &@                      @      &@      "@                               @      @      B@       @      H@       @      @       @      "@      2@      >@      &@       @      8@      M@      M@              "@       @      3@      @      7@      �?      6@      �?      @              @      *@      0@       @      @      *@      ;@      2@              @       @      &@      @      *@      @      :@      �?      �?       @      @      @      ,@      @       @      &@      ?@      D@              @               @      �?      0@      @      =@      "@      0@      (@      (@      @       @      "@      3@      0@      2@     �A@      @      ,@      $@       @      <@      ,@      @      8@      "@      0@       @      &@      @       @       @      .@      &@      2@      >@      @      ,@      $@       @      ;@      @               @      �?      �?      @                      �?              �?      @      @       @       @      @               @      1@      �?               @      �?              @                                              �?       @      �?      �?       @               @      @       @                              �?                              �?              �?       @      @      @      �?      �?                      ,@      &@      @      6@       @      .@      @      &@      @      @       @      ,@       @      *@      6@      @      &@      $@      @      $@      $@      @      4@      @      &@      @      &@      @      @      @      @      @      *@      5@              "@      "@      @       @      �?               @      @      @       @                               @       @      @              �?      @       @      �?       @       @       @      �?      @                      @      �?                      �?      @      @              @                                      �?       @              @                       @                                      @       @               @                                      �?              �?      �?                       @      �?                      �?              @              @                                             �o@     �A@     �e@      $@      ;@      "@      B@     �z@      y@     �D@      B@     @Q@     w@     `n@      @      <@      3@      J@      ,@     �_@      $@     @S@      �?      $@       @      (@     �p@      l@      0@      1@      9@      h@      ^@              @      �?      $@      @      Y@      @      K@      �?       @              "@     @l@      i@      (@      *@      4@     �a@      Y@              �?      �?       @       @     �R@      @     �A@      �?       @              @     ``@     �`@      $@      &@      1@     �[@     @R@              �?      �?      @       @      ;@              .@              �?              �?      9@     �A@       @      @      @      8@      6@                               @              $@              &@                                      8@      ;@       @       @      @      1@      *@                              �?              1@              @              �?              �?      �?       @              �?              @      "@                              �?              H@      @      4@      �?      �?              @     �Z@     �X@       @       @      *@     �U@     �I@              �?      �?      @       @      @              @                              �?     �G@      7@                      @      2@                                                      E@      @      1@      �?      �?              @     �M@      S@       @       @      "@      Q@     �I@              �?      �?      @       @      9@              3@              @               @     �W@     �P@       @       @      @     �@@      ;@                               @              3@              (@               @               @     �O@     �M@      �?       @      @      2@      5@                              �?              .@              &@              �?               @     �M@     �H@      �?      �?      @      2@      ,@                                              @              �?              �?                      @      $@              �?                      @                              �?              @              @              @                      @@      @      �?                      .@      @                              �?              @              @              @                      >@      @      �?                      &@      @                              �?                              @              �?                       @      @                              @                                                      :@      @      7@               @       @      @      C@      9@      @      @      @     �H@      4@              @               @      @      5@              .@                       @      @     �B@      1@      @      @       @      F@      ,@              �?              �?              0@               @                              �?      7@      0@      @       @       @      2@      @              �?                              @              @                                      $@      �?                              $@      @                                              *@              �?                              �?      *@      .@      @       @       @       @      �?              �?                              @              @                       @       @      ,@      �?      �?      �?              :@      $@                              �?              @              @                       @              *@      �?      �?      �?              3@      "@                              �?                                                               @      �?                                      @      �?                                              @      @       @               @                      �?       @              �?      @      @      @              @              �?      @      @      @      @               @                      �?      @                      @      @      @              �?              �?      @      @      @                       @                      �?      @                      �?       @      @                              �?      @              @      @                                                                       @       @      �?              �?                                              @                                              �?              �?              �?                      @                              `@      9@     �W@      "@      1@      @      8@      d@     �e@      9@      3@      F@      f@     �^@      @      6@      2@      E@      "@     �\@      .@     �S@      @      ,@      �?      2@      d@     �d@       @      1@      @@     �d@     @Y@      @      5@      &@      ;@       @     �W@      (@      P@      @      $@      �?      &@     �a@     �a@       @      ,@      8@     @^@      R@       @      1@      "@      6@      @     �Q@      @      D@              @      �?      @     �^@     @Z@      @      "@      ,@      R@      I@              @      @      *@      @      ,@               @                      �?      @      E@     �G@      �?      @       @      4@      0@               @                      @      L@      @      @@              @               @      T@      M@       @      @      (@      J@      A@              @      @      *@       @      9@      @      8@      @      @              @      3@      B@      @      @      $@     �H@      6@       @      &@      @      "@              @              *@      @                      �?      @      &@      @       @      @      &@      "@              "@              @              3@      @      &@      �?      @              @      0@      9@       @      @      @      C@      *@       @       @      @       @              4@      @      ,@       @      @              @      4@      :@              @       @      G@      =@      @      @       @      @      @      �?                              �?                      @      @                                      @                                              �?                                                      @       @                                      @                                                                              �?                      @      �?                                      @                                              3@      @      ,@       @      @              @      *@      7@              @       @      G@      7@      @      @       @      @      @       @      @      *@      �?      @              @      "@      2@              @       @     �@@      2@              �?              @      �?      &@              �?      �?                       @      @      @                              *@      @      @      @       @      �?       @      ,@      $@      1@       @      @      @      @               @      1@       @      (@      $@      6@              �?      @      .@      �?      @      $@      @       @      @      @                       @      1@       @      &@      @      ,@                      @      $@      �?      @       @      @       @      �?      @                       @      .@       @       @      @      ,@                      @      $@      �?      �?              @                       @                      �?      (@              @       @      &@                      @      @              @       @       @       @      �?       @                      �?      @       @      @      �?      @                      �?      @      �?               @                       @       @                      @       @              @                                                              @              $@                              @                                      �?      @       @              �?      �?      @              @              �?                               @                                      �?      @      @              �?      �?       @              @              �?                                                                              @      �?              �?               @                                                               @                                      �?      �?      @                      �?                      @              "@                              @                                               @      @                              @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ^�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         >                   �4@M�]���?�	           ��@       !                     @��"��;�?W            �@                           @�f���?
            �@                           �?x2�g+*�?�           h�@                           �??a0�Di�?�            �u@                          �3@�妹�?`            `c@������������������������       ��|�j��?E             ^@������������������������       �(N:!���?            �A@	       
                    @P�!D!��?w            �h@������������������������       �=�M8���?Z            @c@������������������������       �˲,˲,�?             E@                          �1@(�\Ha�?�            �t@                            �?�Z�Jl^�?G            �X@������������������������       �7�K���?:            �T@������������������������       ��
t�F��?             1@                            �?ɀJ��{�?�            `m@������������������������       ����Q�w�?p            �e@������������������������       �G����?&            �N@                           @�����k�?V           ��@                            �?��Ɂs��?�            pv@                           �?8���`��?�             k@������������������������       ����a1)�?;            @X@������������������������       ��a�|6�?K            �]@                           @I��Np�?\            �a@������������������������       �]�l� �?,             Q@������������������������       ���n~�?0            �R@                           �?W���7�?t            �e@                           �?W3%_�q�?=            �W@������������������������       ��������?             H@������������������������       �K����?"             G@                           �3@���_&�?7            �S@������������������������       �����q�?*            �O@������������������������       �N贁N�?             .@"       /                    �?7�R'��?M           @�@#       (                   �1@\��R٪�?l             e@$       %                   �0@Vr����?'            �Q@������������������������       �d�
��?
             6@&       '                    @��')>Y�?            �H@������������������������       �^�k���?            �A@������������������������       �^N��)x�?	             ,@)       ,                    @ک'N��?E            �X@*       +                   �3@�7�����?5            �S@������������������������       �Ũ�oS��?            �F@������������������������       �t�Qe6�?            �@@-       .                    �?q=
ףp�?             4@������������������������       �9��8���?	             (@������������������������       �      �?              @0       7                    �?���:`��?�            �u@1       4                   �2@*�1%m�?e            �c@2       3                    @rZCVi��?6            �S@������������������������       ��3};��?%            �L@������������������������       ��9����?             6@5       6                   �3@�V)�?/            �S@������������������������       ��F<�A�?             C@������������������������       �q=
ףp�?             D@8       ;                    @��(��?|            @h@9       :                   �3@�z�G!�?h             d@������������������������       �E~�O��?Q             _@������������������������       �n�����?             B@<       =                   �2@%����?             A@������������������������       ��	j*D�?             :@������������������������       �      �?              @?       ^                   �=@h��)u*�?a           �@@       O                    @�Q�����?�           t�@A       H                   �7@��i�#�?            �@B       E                    �?I�$I���?`           ��@C       D                   �6@�6����?�            �m@������������������������       �L(���?g            �c@������������������������       ��⺴
�?1            �S@F       G                     @����Z�?�            @t@������������������������       �LšO��?{            �i@������������������������       �������?M            @]@I       L                    �?AB��?�           `�@J       K                     �?�*�M���?h            �c@������������������������       ����@m�?             �I@������������������������       �tT�A-��?H            �Z@M       N                    �?�3�s�?8           �~@������������������������       �HcT!)��?Z             c@������������������������       ��'�����?�            `u@P       W                    @��� ��?�           �@Q       T                   �;@BĎ�>+�?           P{@R       S                    @2�jp�&�?�            y@������������������������       �/ ��E�?�             p@������������������������       ������ �?U            �a@U       V                    @����[��?             B@������������������������       ����Q��?             .@������������������������       �~VC�1��?             5@X       [                   �5@>î ���?�            �r@Y       Z                     @� G���?0            �U@������������������������       �>����\�?'            �Q@������������������������       �{�/��>�?	             1@\       ]                     @��r]��?�            �j@������������������������       �ףp=
��?d             d@������������������������       ��?��?#            �J@_       f                    �?����?�            �l@`       c                     �?b���Ly�?/            �P@a       b                    @y����0�?            �B@������������������������       ���c����?             :@������������������������       ��ˠT�?	             &@d       e                    @��-�?             =@������������������������       �\���(\�?             4@������������������������       �h/�����?             "@g       l                   �>@��*<�{�?i            @d@h       k                    @����[�?             B@i       j                     �?      �?             8@������������������������       ��r
^N��?             ,@������������������������       ��G�z��?             $@������������������������       �      �?             (@m       p                     @ģ��nH�?O            �_@n       o                    �?(W�7�?3             U@������������������������       ��V����?            �C@������������������������       ���M1j��?            �F@q       r                    @=��<���?             E@������������������������       ��Pk�w�?             9@������������������������       �4%���?
             1@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD        |@     �S@      t@      9@     @R@     �A@     @R@     ��@     `�@     �P@      T@     �f@     �@     �|@      &@     �O@     �I@     `d@      M@     @j@      3@     @Z@      @      (@      @      *@      x@     �s@      (@      5@     �L@     �t@     @c@              1@      @     �I@      *@      a@      &@     �P@       @      @              &@     t@     �n@      @      &@      C@     �k@     @V@               @      @      >@      @     �U@      @     �F@       @                      @     �`@      b@      @      "@      :@     �`@     �M@              @      �?      .@      @     �M@      @      :@                               @      Q@     �H@       @      @      3@      R@      ;@              @              (@      @     �B@      @      @                                     �F@      7@              @       @      :@      @               @                      �?      @@      @      @                                      D@      2@               @       @      ,@      @                                              @               @                                      @      @              �?              (@       @               @                      �?      6@              4@                               @      7@      :@       @              1@      G@      4@              @              (@      @      3@              *@                               @      *@      3@      �?              *@     �D@      0@              @              &@      @      @              @                                      $@      @      �?              @      @      @                              �?              <@      @      3@       @                      @     @P@      X@      @      @      @      O@      @@              �?      �?      @       @      @      @      @                               @      =@      <@              @              1@      @                                              @       @      @                              �?      8@      :@              @              *@      �?                                                      �?      �?                              �?      @       @                              @      @                                              6@              .@       @                       @      B@      Q@      @              @     �F@      <@              �?      �?      @       @      2@              *@       @                       @      4@      J@      �?              @      A@      5@              �?      �?      @       @      @               @                                      0@      0@       @              @      &@      @                                              I@      @      5@              @              @     �g@     �Y@       @       @      (@     @V@      >@               @      @      .@      �?      ;@              $@                              �?      c@      N@       @       @      @     �P@      5@                       @      @      �?      4@              @                              �?     @S@      @@      �?       @      @     �J@      1@                       @       @      �?      @               @                                      E@      ,@                       @      >@      @                                              1@              �?                              �?     �A@      2@      �?       @      @      7@      *@                       @       @      �?      @              @                                     �R@      <@      �?               @      ,@      @                              @              @              @                                     �D@      @      �?                      $@       @                                              @              @                                      A@      5@                       @      @       @                              @              7@      @      &@              @              @      B@      E@                      @      6@      "@               @       @       @              0@              @                                      <@      8@                      @      $@      @                                               @              �?                                      3@      &@                      �?      @      @                                               @              @                                      "@      *@                       @      @      �?                                              @      @      @              @              @       @      2@                       @      (@      @               @       @       @              @      @       @                              @       @      0@                              &@      @              �?       @      @              @               @              @                               @                       @      �?                      �?              �?             @R@       @     �C@      �?      "@      @       @     @P@     �Q@      @      $@      3@      \@     @P@              "@       @      5@      @     �B@      @      *@              @      @      �?      ,@      6@       @              @      B@      *@               @               @      �?      ,@              @              @                      $@      (@       @              @      1@       @                                              @                                                      @      @                              @                                                       @              @              @                      @      @       @              @      (@       @                                              @                              @                      �?      @       @              @      "@       @                                              �?              @                                      @      �?                       @      @                                                      7@      @      "@               @      @      �?      @      $@                      �?      3@      &@               @               @      �?      6@      @       @               @      @               @      "@                      �?      0@      @              �?               @      �?      &@       @       @                                      �?      @                              $@      @              �?               @              &@       @                       @      @              �?      @                      �?      @       @                                      �?      �?              @                              �?       @      �?                              @      @              �?                              �?              @                                      �?      �?                               @      @                                                              @                              �?      �?                                      �?                      �?                              B@      @      :@      �?      @              �?     �I@     �H@      @      $@      (@      S@      J@              @       @      *@      @      2@              &@                              �?     �B@      6@       @      @      @      >@      .@              @              @      @      *@              @                                      =@       @       @                      0@      @               @              �?              $@              @                                      :@      �?                              (@      @                                              @                                                      @      @       @                      @                       @              �?              @              @                              �?       @      ,@              @      @      ,@      &@              �?              @      @       @               @                              �?       @      "@              @       @      @      "@              �?                      @      @              @                                      @      @              @       @      $@       @                              @              2@      @      .@      �?      @                      ,@      ;@      �?      @       @      G@     �B@              @       @       @       @      .@      @      ,@      �?      @                       @      1@      �?      @      @     �E@      A@               @       @      @      �?      &@      @      &@      �?      @                       @      (@              @      @      ;@      <@               @       @      @      �?      @      �?      @                                              @      �?                      0@      @                                              @              �?                                      @      $@                      @      @      @               @              �?      �?       @                                                      @      @                      @       @      @               @              �?      �?      �?              �?                                              @                              �?                                                     �m@     �M@      k@      6@     �N@      @@      N@      b@     �m@     �K@     �M@     @_@     0s@     �r@      &@      G@      F@      \@     �F@     `l@      K@     �h@      .@     �G@      4@      L@     �a@     �k@     �C@     �G@     �X@     0r@     0q@       @     �C@     �B@     �X@     �A@      a@      ?@     @`@      (@     �B@      4@      E@      F@      _@      9@      @@      R@     �e@     `g@      @      =@      ;@     �M@      =@     �S@      &@     �P@      @      "@      &@      1@      8@     �K@      0@      1@      A@      W@     �P@       @      "@      *@      :@       @      E@      �?      C@       @      @      @      @      .@      6@      �?       @      *@      H@      <@       @       @      �?      @      �?      4@              8@       @      @      @       @      *@      .@              �?      @     �B@      6@               @      �?      @      �?      6@      �?      ,@              �?               @       @      @      �?      �?       @      &@      @       @                      �?              B@      $@      =@       @      @      @      *@      "@     �@@      .@      .@      5@      F@     �C@              @      (@      5@      @      >@      @      4@                               @      @      9@      @      @      "@      @@      ?@              @      @      .@      @      @      @      "@       @      @      @      @      @       @       @      "@      (@      (@       @              @      @      @       @      M@      4@     �O@       @      <@      "@      9@      4@     @Q@      "@      .@      C@      T@      ^@       @      4@      ,@     �@@      5@      6@      @      &@      @      @               @      @      =@      @      @      @      3@      7@              @      @      $@      �?      @              �?       @      @                      �?      1@      �?              �?      @       @                      �?      @              1@      @      $@      @       @               @      @      (@       @      @      @      .@      .@              @       @      @      �?      B@      0@      J@      @      5@      "@      7@      ,@      D@      @      (@      ?@     �N@     @X@       @      1@      &@      7@      4@      1@      @      $@               @      �?      @      @      &@      @      @      @      ;@      9@              @      �?      $@      $@      3@      "@      E@      @      *@       @      3@      "@      =@       @       @      ;@      A@      R@       @      *@      $@      *@      $@     �V@      7@     @Q@      @      $@              ,@     �X@     @X@      ,@      .@      :@     �]@      V@      @      $@      $@      D@      @     �I@      ,@      <@              @              @      R@      N@      @      $@      .@     �T@     �K@       @       @      @      .@      @     �F@      &@      <@              @              @     �Q@     �M@      @      @      .@     �P@     �K@      �?      @      @      .@      @     �A@      "@      7@              @               @      B@     �A@      @      @      .@      A@     �E@              �?      �?      $@      �?      $@       @      @               @              @      A@      8@               @              @@      (@      �?      @      @      @      @      @      @                                               @      �?      �?      @              0@              �?      @                              @                                                                                              "@                                                              @                                               @      �?      �?      @              @              �?      @                              D@      "@     �D@      @      @              "@      :@     �B@      $@      @      &@     �B@     �@@       @       @      @      9@      �?      2@              "@               @              @      *@      .@       @       @      @      @       @                              @      �?      0@              @               @               @      &@      .@               @      @      @      @                              @      �?       @              @                              @       @               @                               @                                              6@      "@      @@      @      �?              @      *@      6@       @      @      @      @@      9@       @       @      @      6@              5@      @      >@      @                      �?      &@      2@      @      @      @      2@      *@               @      @      1@              �?      @       @              �?              @       @      @      �?              �?      ,@      (@       @                      @              &@      @      2@      @      ,@      (@      @       @      1@      0@      (@      ;@      0@      ;@      @      @      @      *@      $@      $@       @      �?               @               @              @       @      @      @      $@      (@      �?      @      �?               @       @       @      �?                               @              @       @      @      @      �?      @              @                      �?      @       @                                      �?              @       @      @      @              �?              @                      �?      @              �?                              �?              �?                              �?      @                                               @                               @                              �?              @              "@      @      �?       @      �?              �?       @                               @                                              @              @      @      �?       @      �?              �?                                                                      �?                              @      @                                              �?      @      1@      @      (@      (@       @       @      &@      ,@      @      7@      @      .@       @       @      @      *@       @              �?      @      �?      @       @                      �?               @      �?       @      "@                      �?      @                      �?      @      �?      @       @                      �?               @              �?      @                      �?      @                      �?       @              �?       @                      �?                              �?      @                      �?       @                               @      �?      @                                               @                                                      �?                                                                                                      �?      �?      @                              @              �?       @      *@      @      @      $@       @       @      $@      ,@      @      6@      @      @       @       @      @      @       @      �?              (@      @      @      @       @              @      $@      �?      4@      @      @              �?       @      @      �?                      @      @      @      @                      �?      �?      �?      .@              �?              �?      �?      @      �?      �?               @              @               @              @      "@              @      @      @                      �?      @                       @      �?       @      �?      @               @      @      @      @       @               @       @      �?      @              @               @              �?      �?      @                      @      @      �?       @               @      �?      �?      �?              �?                      �?      �?               @               @                       @                              �?               @              @�t�bub��      hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ>*xhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKyhnh4h7K ��h9��R�(KKy��hu�Bx         >                    �?V��j��?�	           ��@                           �??s�z�?!           �@                           �?��g���?�           H�@                           @羅�?�            q@                            �?K׆���?            �i@                           �?��X#��?O            �_@������������������������       �]4��!�?&            �M@������������������������       ��ҼI�?)            �P@	       
                   �6@
ףp=��?0             T@������������������������       �	6c����?            �I@������������������������       � �^�@��?             =@                           @۝����?(            �P@������������������������       �*L�9��?             F@                          �4@��JÝ�?             7@������������������������       ���!pc�?             &@������������������������       �r�q��?             (@                            @ɖd2 ��?           �y@                           �?���6F��?�            `j@                            �?�G�z��?4             T@������������������������       ��2����?+            �P@������������������������       ��T�6|��?	             *@                          �3@8{�$��?Q            ``@������������������������       ����U��?             A@������������������������       � ��qg��?>            @X@                          �3@+�%sP��?�            �h@                           �?��O�+�?&             K@������������������������       �躍`3�?             1@������������������������       �J�?�b�?            �B@                          �=@��Œ���?d            �a@������������������������       �h}(�=T�?[             `@������������������������       �����X�?	             ,@        /                    �?��S̪=�?k           Ȏ@!       (                   �5@b�|=���?�            �v@"       %                    �?��)Jk�?b            @e@#       $                   �4@�2q�{�?             E@������������������������       ��Էr�?            �@@������������������������       ��<ݚ�?             "@&       '                    @     s�?J             `@������������������������       �|���?$            �P@������������������������       �6�`��V�?&             O@)       ,                   �<@�� ����?            @h@*       +                   �6@�G�z��?g             d@������������������������       ���	h"�?             I@������������������������       ���W�J�?L            �[@-       .                   �?@�V�e�t�?             A@������������������������       �S�!�uq�?             9@������������������������       ��2�tk~�?             "@0       7                    �?�#y��D�?�           h�@1       4                     @ z��/?�?l            �c@2       3                     �?֌��^�?=            �U@������������������������       �����?            �F@������������������������       ��ܤ��?             E@5       6                   �4@>�֕�?/            �Q@������������������������       ��������?             B@������������������������       ��g+�v�?             A@8       ;                    @	�|/D�?            }@9       :                   �4@R�
�%��?G            @\@������������������������       �     ��?             @@������������������������       ����k���?5            @T@<       =                   �6@��n;�X�?�            �u@������������������������       �r��ճC�?k             f@������������������������       �����?l            �e@?       Z                    @S�����?�           ��@@       O                    @���Ol��?5           0�@A       H                   �1@�@?��?>           �@B       E                     @�65��?�            �m@C       D                    �?ZAl��?{             f@������������������������       ��u����?D            �Y@������������������������       �b��^��?7            �R@F       G                    @� =�	��?(             O@������������������������       �(}�'}��?             >@������������������������       �     ��?             @@I       L                   �9@�D�mVA�?�           \�@J       K                     �?\�����?            ��@������������������������       �Ϋ�gE��?7            ~@������������������������       �_|�!��?�             w@M       N                     @,9��HA�?{            �h@������������������������       �03�i�3�?d            �c@������������������������       ���Q��?             D@P       W                    @�cް�?�            `x@Q       T                   �0@6Ws5Ws�?�            �v@R       S                    �?���{��?             I@������������������������       ���8��8�?             B@������������������������       ��X�C�?             ,@U       V                   �8@,yi��?�            �s@������������������������       ��xGQ[�?�             q@������������������������       ��������?             D@X       Y                   �4@�k���B�?             :@������������������������       ��q�q�?             (@������������������������       ���S�r
�?             ,@[       j                   �5@��p�U�?w           ؁@\       c                     @�hP�vC�?�            �t@]       `                     �?؎mz��?�             o@^       _                    �?hs��h�?            �h@������������������������       �M��>z�?2             Q@������������������������       �LΞ��i�?M             `@a       b                   �1@�wɃg�?!             J@������������������������       ��q�q�?
             (@������������������������       ���Q��?             D@d       g                    �?%���Qz�?.            �S@e       f                   �3@4�����?             ?@������������������������       �B{	�%��?             "@������������������������       ��J����?	             6@h       i                    @UUUUU��?             H@������������������������       ��i�6��?             >@������������������������       ��n���?             2@k       r                    �?����?�            `n@l       o                   �:@�/鳗�?H            @Y@m       n                     @�������?1             R@������������������������       �����>4�?'             L@������������������������       �      �?
             0@p       q                   �;@^s]ev�?             =@������������������������       ��zv��?             &@������������������������       �Ix�5?�?             2@s       v                   �>@mv$Ҷ��?a            �a@t       u                     �?6�����?T            �^@������������������������       �ie��#�?)            �N@������������������������       �� �kRB�?+            �N@w       x                    @��(\���?             4@������������������������       ����!pc�?             &@������������������������       ��n���?             "@�t�bh�h4h7K ��h9��R�(KKyKK��h��B�G       ~@     @T@     t@      @@     @Q@      ?@      Q@     ��@     ��@      Q@     �S@     �e@     ��@     �{@      ,@     �J@     �J@      `@      P@     �i@      E@     �c@      4@     �C@      1@      C@     @a@     @f@      ?@     �J@     �W@      l@     `m@      &@      :@      ?@     �Q@      L@     �U@      &@      M@      @      ,@      �?      &@     @U@      V@      @      0@      >@     �\@      T@      @      *@      *@      ;@      5@      B@      @      .@              @               @      D@      J@      @      @      ,@     �H@      6@              @      @      @       @      ?@      @      .@              @              �?      @@     �C@      @      �?       @      A@      3@              @      @      @      @      8@      @      @              @              �?      &@      <@       @      �?       @      .@      ,@               @       @       @      @      @      @      @                                      @      3@              �?       @      @      @                       @       @      @      2@               @              @              �?      @      "@       @              @      $@      "@               @                      �?      @              "@                                      5@      &@       @                      3@      @              �?       @      �?       @      @               @                                      3@       @                              .@      @              �?              �?              �?              @                                       @      "@       @                      @                               @               @      @       @                                      �?       @      *@       @      @      @      .@      @              @              @       @      @       @                                              @      @       @      �?      @      $@      @              @              �?              �?                                              �?      @      @               @              @                                      @       @                                                                      @               @               @                                      �?              �?                                              �?      @                                      @                                       @       @      I@      @     �E@      @      &@      �?      "@     �F@      B@              (@      0@     @P@      M@      @      @      "@      4@      *@      =@      @      5@      �?      @              @      9@      2@              $@      @      >@      ?@              @      @      $@      @      .@      �?      @      �?       @              �?      0@      @              @       @      "@      &@              �?              @              $@      �?      @      �?       @              �?      ,@      @              @      �?      "@      &@                              @              @               @                                       @      �?                      �?                              �?              �?              ,@      @      .@              @              @      "@      *@              @      @      5@      4@               @      @      @      @       @                                                      @       @                              $@                                              @      @      @      .@              @              @      @      @              @      @      &@      4@               @      @      @      @      5@              6@      @      @      �?      @      4@      2@               @      $@     �A@      ;@      @      @      @      $@      @      @              @                              �?      ,@      @                      @      &@      @              �?              @      �?       @                                                              @                              @      @                              @              �?              @                              �?      ,@       @                      @      @       @              �?              �?      �?      2@              3@      @      @      �?       @      @      *@               @      @      8@      6@      @      @      @      @      @      ,@              3@      @      @      �?       @      @      *@               @      @      8@      5@              �?      @      @      @      @                              �?                                                                      �?      @       @      �?               @     �]@      ?@     �X@      0@      9@      0@      ;@     �J@     �V@      9@     �B@      P@     �[@     `c@       @      *@      2@      F@     �A@     �M@      $@      @@      @      $@       @      @      9@      B@      @      *@      :@      K@     �E@              @       @      ,@      *@      =@      @      ,@              �?                      1@      =@      @      @      3@      5@      &@              �?      @      @      @      "@              �?              �?                      (@       @              @      @       @                                      �?              "@                              �?                      (@      @              �?      �?       @                                      �?                              �?                                               @               @      @                                                              4@      @      *@                                      @      5@      @      @      ,@      3@      &@              �?      @      @      @      @      @       @                                      @      @              @      "@      ,@      @              �?                      @      .@              @                                       @      ,@      @              @      @      @                      @      @      �?      >@      @      2@      @      "@       @      @       @      @      @      @      @     �@@      @@               @      @       @      "@      =@      @      ,@      @      @       @              @      @      @      @      @     �@@      =@               @      �?      @       @      @              @      @                              �?      @       @                      @      "@               @              @      �?      6@      @      "@              @       @              @      �?      �?      @      @      :@      4@                      �?      �?      @      �?      �?      @              @              @       @                      @      @              @                      @      �?      �?              �?       @              @              @       @                              �?              @                      @      �?      �?      �?               @              �?                                              @       @                                                              N@      5@     �P@      (@      .@      ,@      5@      <@      K@      3@      8@      C@     �L@      \@       @      $@      $@      >@      6@     �A@      @      .@       @      @      @      @       @      .@      �?              @      6@      6@      �?              @      @      @      6@      �?      @              �?              @      @      "@      �?              @       @      3@      �?              @      @      �?      *@                              �?                              @                       @      @      &@      �?              @      @              "@      �?      @                              @      @      @      �?               @      @       @                                      �?      *@      @      $@       @      @      @              @      @                      @      ,@      @                              �?       @      (@      @      @              @                      @      @                      �?      @      @                              �?              �?              @       @       @      @                      @                       @      $@                                               @      9@      1@     �I@      $@      "@      "@      2@      4@     �C@      2@      8@      ?@     �A@     �V@      @      $@      @      9@      3@       @      "@      ,@       @       @              @      @      &@       @      @      �?      &@      :@       @      @      @      @      @      �?              (@                                      �?      @               @              @       @                              @              �?      "@       @       @       @              @      @      @       @       @      �?      @      8@       @      @      @      @      @      7@       @     �B@       @      @      "@      &@      0@      <@      0@      4@      >@      8@      P@      @      @      @      2@      0@      0@      @      .@      @              �?      @      0@      2@      @      @      $@      2@     �E@                      �?      *@      @      @      @      6@      @      @       @      @              $@      $@      0@      4@      @      5@      @      @      @      @      *@     @q@     �C@     �d@      (@      >@      ,@      >@     �z@      |@     �B@      :@     �S@     �t@      j@      @      ;@      6@      M@       @     �g@      9@     @^@      @      :@      (@      9@     `u@     v@      :@      2@      N@     0p@      b@      �?      .@      $@      A@      @     �c@      5@     @Y@      @      8@      (@      4@     @k@     @p@      :@      (@     �H@      i@     @]@              ,@      $@      @@      @      8@      @      *@                               @     @U@     �O@      @      �?      @      >@       @                               @      �?      .@      @      "@                               @     @R@     �G@              �?       @      3@      @                              �?      �?      &@       @                                       @      J@      <@                      �?      @                                      �?              @      �?      "@                                      5@      3@              �?      �?      *@      @                                      �?      "@              @                                      (@      0@      @               @      &@      @                              �?              �?                                                      @      (@      @              �?       @      �?                              �?               @              @                                      "@      @                      �?      @      @                                             �`@      2@      V@      @      8@      (@      2@     �`@     �h@      7@      &@     �F@     @e@     @[@              ,@      $@      >@      @     �\@      (@     �Q@      @      @      @      *@     �^@      f@      $@      "@     �B@     �b@     �S@              @       @      0@       @      P@      @     �B@      @      �?      �?      @     �I@     @[@      @      @      7@     @U@     �J@              @       @      *@             �I@       @      A@       @      @      @      @      R@     �P@      @      @      ,@      P@      :@                              @       @      3@      @      1@              1@      @      @      $@      5@      *@       @       @      5@      >@              @       @      ,@       @      .@      @      &@              1@      @       @       @      0@      *@       @      @      3@      6@              @       @      &@      �?      @      �?      @                              @       @      @                      @       @       @                              @      �?     �@@      @      4@               @              @      _@     @W@              @      &@     �M@      <@      �?      �?               @      �?      ?@      @      3@               @              @     �^@     �V@              @      &@      F@      :@      �?      �?               @      �?      @                                                     �@@      "@                      @      �?                                                      @                                                      9@      @                              �?                                                      �?                                                       @       @                      @                                                              ;@      @      3@               @              @     @V@     @T@              @       @     �E@      :@      �?      �?               @      �?      6@      �?      ,@                              @     �U@      S@              @      @     �@@      8@      �?      �?               @      �?      @      @      @               @              �?      @      @               @       @      $@       @                                               @              �?                              �?       @      @                              .@       @                                               @                                                      �?      @                              @      �?                                                              �?                              �?      �?                                      $@      �?                                             @U@      ,@      F@      @      @       @      @     @U@     @X@      &@       @      3@      S@      P@       @      (@      (@      8@       @     �J@      @      0@               @                     �Q@     @P@      @      @      &@      G@      A@              $@       @       @      �?      F@      @      (@               @                      J@     �L@       @      �?      &@      =@      2@               @       @      @      �?      A@      @      "@              �?                     �F@      B@       @      �?      &@      8@      ,@               @       @      @      �?      @              @                                      1@      0@                       @       @      &@              �?       @      �?              ;@      @      @              �?                      <@      4@       @      �?      "@      0@      @              @              @      �?      $@              @              �?                      @      5@                              @      @                              �?              @                                                      @       @                              �?       @                                              @              @              �?                      @      3@                              @       @                              �?              "@              @                                      3@       @      �?       @              1@      0@               @              �?              @                                                      @                                      @      *@               @                                                                                       @                                      @       @               @                              @                                                      @                                              &@                                              @              @                                      (@       @      �?       @              ,@      @                              �?              @              @                                      $@      @               @              @       @                                                                                                       @      @      �?                      $@      �?                              �?              @@      &@      <@      @       @       @      @      ,@      @@       @      @       @      >@      >@       @       @      $@      0@      �?      3@      @      @      �?                               @      8@      @      @      �?      .@       @              �?              @      �?      .@      @       @                                      @      5@       @      @              "@      @              �?              @              ,@      @       @                                      @      0@              @              @      @                              �?              �?                                                       @      @       @                      @                      �?               @              @      @       @      �?                              �?      @      �?      �?      �?      @      @                               @      �?       @      �?                                                              �?      �?              @                                       @               @       @       @      �?                              �?      @                      �?       @      @                                      �?      *@      @      8@      @       @       @      @      @       @      @              @      .@      6@       @      �?      $@      &@              $@      @      1@      @       @              @      @      @      @              @      .@      6@       @      �?      $@      $@              @              &@      @                      �?      @       @                      @      &@      @              �?       @      @              @      @      @      �?       @               @              @      @              �?      @      .@       @               @      @              @              @                       @       @              �?      �?              @                                              �?              @              @                       @                      �?      �?                                                              �?                              @                               @                                      @                                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��khG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKohnh4h7K ��h9��R�(KKo��hu�BH         8                    �?�x-ω��?�	           ��@                          �2@t�:-?�?'           �@                           �?ᗭ��?�            Pu@                           @R�;&	��?T            @`@                           @�̚��?M            �^@                            �?4ܪ'z�?&            �O@������������������������       ���R[s�?            �A@������������������������       ���X��?             <@	       
                   �1@�������?'            �M@������������������������       ��a�2�t�?             B@������������������������       ��\@˜��?             7@������������������������       �      �?              @                          �1@�`+H��?�            `j@                            @�h
uI�?C            �[@                            �?�
Yg��?!            �J@������������������������       ��ˠT��?             6@������������������������       �p��N�?             ?@                           �?|�%~oI�?"            �L@������������������������       ��"w����?             3@������������������������       ��].��?             C@                           @�/鳗�?@            @Y@                           @�*3��F�?1            �S@������������������������       �ܚ�R��?             G@������������������������       �     0�?             @@                           �?�r��_�?             7@������������������������       �R���Q�?             $@������������������������       ��T�6|��?             *@       +                    @��b�?P           ��@       $                     �?��~�)�?           ؈@       !                    �?����"��?�            �n@                            �?����i2�?Q            �`@������������������������       �G ��h�?            �E@������������������������       �C��/\��?6            �V@"       #                    �?��Nݍ�?G            @\@������������������������       ��2q�{�?             E@������������������������       ���>�S�?-            �Q@%       (                    �?�s���:�?o            �@&       '                     �?挛:|�?�            @r@������������������������       ���K7�A�?D             Y@������������������������       �������?�             h@)       *                     �?    @D�?�             p@������������������������       �,R�n��?-             R@������������������������       �SvLB�?z             g@,       3                   �>@�qi���?I           X�@-       0                    �?J��J�i�?*           �}@.       /                   �8@X�	�S)�?g            �d@������������������������       �
^N��)�?G             \@������������������������       �~4��?             �J@1       2                   �4@�)q$D�?�            `s@������������������������       ��$ğӯ�?*            �O@������������������������       ���<;k�?�            �n@4       5                    @9��8�#�?             H@������������������������       ���8��8�?	             (@6       7                   �@@����H�?             B@������������������������       �ƵHPS!�?             *@������������������������       ���/��@�?             7@9       V                   �2@��+���?�           ��@:       G                    @C��|�?�           x�@;       B                     @�#R����?_             c@<       ?                   �1@4�~#��?C            �Z@=       >                   �0@�����?+            �P@������������������������       ��h9����?            �B@������������������������       ��;N��?             =@@       A                     �?��Z���?            �D@������������������������       �v��`��?             =@������������������������       ��������?             (@C       D                    �?��4c�?             G@������������������������       �����W�?	             *@E       F                    �?h�����?            �@@������������������������       �)O���?	             2@������������������������       �������?
             .@H       O                   �0@��\���?W           ��@I       L                    �?6<�R��?>             Y@J       K                    �?�q���?             H@������������������������       ����ؓ�?             ?@������������������������       �8߄*�u�?
             1@M       N                    @���3�E�?!             J@������������������������       ����B�(�?            �A@������������������������       �*�8�G��?	             1@P       S                   �1@�8.j��?            {@Q       R                    @Gi�e��?�            �k@������������������������       �f�z`��?g            �c@������������������������       ���M��?)             O@T       U                    @�xWx��?�            �j@������������������������       �:e��^��?k            �d@������������������������       �UUUUU��?             H@W       f                   �8@N$�ɲ}�?�           |�@X       _                     @L��G�?�           ��@Y       \                    �?�ٕ-n��?T           H�@Z       [                     �?k���f�?�            �v@������������������������       ��A;����?�            �n@������������������������       ���?N��?G            @\@]       ^                     �?�3�z�A�?n           �@������������������������       �1*�a��?           z@������������������������       ����(\�?h             d@`       c                    �?P�4��>�?�            �j@a       b                    @Y�5�?A            �Y@������������������������       �ްS��k�?(            �M@������������������������       ����#���?             F@d       e                   �5@���}�?I            �[@������������������������       �/�6�G��?-            @Q@������������������������       ���뺮��?             E@g       n                   @A@��9J'�?
            z@h       k                    @������?            �x@i       j                    @�:��]��?�            �p@������������������������       �vo��?w            �f@������������������������       ��R���?;            @U@l       m                    �?     �?N             `@������������������������       ���;�?             =@������������������������       �y�R��{�?9            �X@������������������������       ���(\���?
             4@�t�bh�h4h7K ��h9��R�(KKoKK��h��B�A       `y@     �T@     Pv@      G@     �P@      <@     �X@     �@     ��@     @R@     @U@      f@     @�@     �z@      *@     @R@     �I@     �[@     @P@      f@      C@     `f@      9@      H@      4@      I@      ^@      i@     �@@      I@     @Y@      l@     @h@      "@     �D@      B@     @Q@      F@     �F@      @      B@      �?      @              @      L@     �P@      �?       @      ,@      J@      9@              @      �?      &@      @      2@      �?      $@                               @     �A@      7@              �?      @      4@      @              @              @              .@      �?       @                               @     �A@      6@                      @      4@      @              @              @              @      �?      @                               @      1@      "@                       @      @      @              @              @              @              @                                      *@      "@                       @      �?      @                                              @      �?      @                               @      @                                      @       @              @              @               @               @                                      2@      *@                      @      ,@                                                      @               @                                      *@      &@                              @                                                       @                                                      @       @                      @      $@                                                      @               @                                              �?              �?                                      �?                              ;@      @      :@      �?      @              @      5@      F@      �?      @       @      @@      3@               @      �?      @      @      .@              &@              @                      .@      3@              @      @      0@      &@               @      �?      @       @       @               @              �?                      @      ,@              �?      @      (@       @                              �?       @      �?                                                      @       @              �?      �?       @       @                                      �?      @               @              �?                              @                      @      $@                                      �?      �?      @              "@              @                      "@      @              @      �?      @      "@               @      �?       @              @                              @                      �?       @              @              @       @                                              @              "@                                       @      @                      �?      �?      @               @      �?       @              (@      @      .@      �?                      @      @      9@      �?      @      @      0@       @                              @      �?      @      @      $@      �?                      @      @      7@      �?      @      @      &@      @                              @              @      @      @                                      @      $@              @      �?      "@      @                              @               @              @      �?                      @              *@      �?               @       @      @                              �?              @              @                                      @       @                              @       @                                      �?      �?              @                                               @                              @                                              �?      @               @                                      @                                       @       @                                             �`@      A@     �a@      8@      E@      4@     �F@      P@     �`@      @@      E@     �U@     �e@      e@      "@     �A@     �A@      M@     �D@     �W@      ,@     @T@      .@      ?@      $@      1@      D@     @V@      *@      5@      H@     �Z@     �[@      @      6@      2@     �A@      5@      ?@      "@      5@      @       @              "@      @     �@@      @       @      0@     �D@      A@       @      @      @      2@      @      8@       @      &@               @              @      @      5@      @              @      6@      (@       @      �?      @      0@              @              @               @              �?      �?      &@                       @      (@      �?                      @       @              5@       @      @                              @       @      $@      @              @      $@      &@       @      �?              ,@              @      @      $@      @                      @       @      (@      @       @      $@      3@      6@              @      �?       @      @              @       @      @                                      @                      @      .@      @              �?              �?       @      @      @       @       @                      @       @      @      @       @      @      @      2@              @      �?      �?       @      P@      @      N@      $@      =@      $@       @     �A@      L@      @      3@      @@     �P@     @S@      @      1@      ,@      1@      1@      @@      @     �C@      @      0@      @      @      ,@      =@      @      *@      *@      @@     �H@      @      @      @      @      @      .@       @      2@              �?              @      @      &@               @      @      $@      .@                                      @      1@      @      5@      @      .@      @              @      2@      @      @      "@      6@      A@      @      @      @      @      @      @@              5@      @      *@      @      @      5@      ;@              @      3@      A@      <@       @      &@      @      $@      $@      &@               @       @      @              �?      &@      @              �?      @      @      @              @      @               @      5@              *@      @      "@      @       @      $@      8@              @      0@      =@      5@       @      @      @      $@       @     �B@      4@      O@      "@      &@      $@      <@      8@     �F@      3@      5@     �C@     @P@      M@       @      *@      1@      7@      4@      B@      4@      K@      @      @      @      :@      8@      F@      1@      5@      ?@     @P@      M@              *@       @      6@      2@      4@       @      $@              �?              @      *@      0@      $@       @      $@      <@      ,@              @      @      $@       @      0@      �?      @                              @      $@      *@      @       @      @      (@      (@              �?      @      @      @      @      �?      @              �?              �?      @      @      @              @      0@       @              @      �?      @      @      0@      2@      F@      @      @      @      4@      &@      <@      @      *@      5@     �B@      F@               @      @      (@      $@      @              4@                                      @      @      �?      @      @      $@      @                              @              &@      2@      8@      @      @      @      4@      @      8@      @      $@      2@      ;@     �B@               @      @      @      $@      �?               @      @      @      @       @              �?       @               @                       @              "@      �?       @                      �?               @      �?                      �?                      �?                                      @                      �?              @      @       @       @       @                       @              @                       @              @      �?       @      �?                      @               @       @                                       @                                      @                                      @       @       @                                       @              @                       @                      �?       @     �l@     �F@     @f@      5@      3@       @     �H@     �z@     pz@      D@     �A@     �R@     �v@      m@      @      @@      .@     �D@      5@     @R@      @      J@                              @     `l@     �c@      @      "@      $@     �W@      F@               @              @       @      2@              (@                                      ;@      K@      @      @      �?      6@      $@              �?                              ,@              "@                                      6@     �D@       @      @      �?      @      @              �?                              @              @                                      0@      =@              @              @                                                      �?              @                                      @      4@               @              @                                                      @              @                                      "@      "@               @              @                                                      $@              @                                      @      (@       @              �?              @              �?                              @              �?                                      @      @       @              �?              @              �?                              @               @                                       @      @                                                                                      @              @                                      @      *@      �?      �?              .@      @                                              @                                                              @                              @      �?                                                              @                                      @      $@      �?      �?              $@      @                                                                                                      @       @      �?                      @                                                                      @                                      �?       @              �?              @      @                                             �K@      @      D@                              @      i@     @Z@              @      "@     @R@      A@              �?              @       @      0@              �?                                      P@      $@                              @      �?                              �?              @                                                      D@      @                               @                                                       @                                                      9@       @                               @                                                      �?                                                      .@      �?                                                                                      *@              �?                                      8@      @                              @      �?                              �?              @                                                      2@      @                               @      �?                              �?              @              �?                                      @      �?                              @                                                     �C@      @     �C@                              @      a@     �W@              @      "@     �P@     �@@              �?              @       @      8@       @      *@                              �?      P@      N@              @      @      A@      $@                               @              *@      �?       @                              �?      H@     �I@              @      @      3@       @                                              &@      �?      @                                      0@      "@                      �?      .@       @                               @              .@       @      :@                               @      R@     �A@                      @      @@      7@              �?              �?       @      $@              4@                              �?      P@      8@                      �?      :@      2@                                       @      @       @      @                              �?       @      &@                       @      @      @              �?              �?             �c@     �D@     �_@      5@      3@       @      G@     �h@     �p@     �B@      :@     @P@     �p@     �g@      @      >@      .@     �B@      3@     @`@      4@     �T@      0@       @       @      =@     `e@      k@      4@      ,@      F@     �g@      b@       @      1@      @      :@      (@      Z@      0@     �Q@      "@       @      �?      3@     �b@     @h@      0@      *@     �A@      c@     �Y@      �?      *@      @      4@       @     �@@      @      8@              �?      �?      @      L@      W@      �?      �?       @     �L@     �M@              @      �?      @      @      .@      �?      1@              �?      �?      @      B@     �N@      �?      �?      @      F@      I@              @      �?      @      �?      2@      @      @                              �?      4@      ?@                      �?      *@      "@              @              �?       @     �Q@      "@      G@      "@      @              ,@      W@     �Y@      .@      (@      ;@      X@     �E@      �?      @      @      0@      @      M@      @      C@      "@      @              *@     �O@     �Q@      (@      &@      1@      L@      A@              @      @      $@      @      *@      @       @              @              �?      =@      @@      @      �?      $@      D@      "@      �?                      @              :@      @      (@      @              �?      $@      7@      6@      @      �?      "@      C@      E@      �?      @              @      @       @              @       @              �?      @      .@       @      @      �?      �?      9@      7@              @              @              @              �?       @              �?              $@      @              �?      �?      2@      $@                              @              @              @                              @      @      @      @                      @      *@              @                              2@      @       @      @                      @       @      ,@                       @      *@      3@      �?      �?              �?      @      *@      @      @      @                      @      @       @                      @      @      @              �?              �?       @      @              �?                              �?      @      @                      @      @      (@      �?                               @      :@      5@      F@      @      &@      @      1@      <@      H@      1@      (@      5@     �R@     �F@       @      *@       @      &@      @      :@      3@     �D@      @      &@      @      .@      <@      H@      $@      (@      3@     �R@     �E@       @      *@       @      &@      @      0@      @      3@       @      &@      @       @      0@     �C@      @      "@      *@      M@      ?@       @      "@      @      @      @      ,@      @      ,@       @      @      @      @      "@      2@      @      @      $@     �B@      6@       @      "@      @      @      @       @      @      @              @               @      @      5@              @      @      5@      "@                       @      �?              $@      (@      6@      @                      @      (@      "@      @      @      @      0@      (@              @       @      @      @              @                                      @      @      @      �?              �?       @      @               @      �?      �?      �?      $@      "@      6@      @                      @      @      @       @      @      @      ,@      "@               @      �?      @       @               @      @                       @       @                      @               @               @                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJH-�@hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKuhnh4h7K ��h9��R�(KKu��hu�B�         <                   �7@��5�?��?�	           ��@       !                    �?h*p���?�           h�@                          �1@�x�?P           ��@                          �0@:8�L�w�?�            �t@                           @�T���?G            �]@                           @���Hx�?+             R@������������������������       �VUUUU��?             H@������������������������       ��q�q�?             8@	       
                    @Ya�)��?            �G@������������������������       ���W64<�?             ?@������������������������       �     @�?	             0@                            @c
Gb�F�?�            �j@                           �?t��G0��?_            �c@������������������������       �lv�"��?             5@������������������������       �������?S             a@                           @�0�Qy�?"            �K@������������������������       ���"e���?             ;@������������������������       ��Cc}�?             <@                           @�v7&q��?�           ��@                           @�닿�?�           ��@                          �5@@�ꌅ��?�            �x@������������������������       �S:.����?�            �r@������������������������       �5h0zF�?A            �X@                            @���"��?�            @m@������������������������       ��G�z4�?c             d@������������������������       ��H
����?5            �R@                            @� &�m�?�            �w@                           @��b��?�            `s@������������������������       �<pƵ��?�             j@������������������������       �s	�6�c�?C            �Y@                            �?r����B�?*            @Q@������������������������       ��8��8��?             8@������������������������       �#���[�?            �F@"       1                     @���7���?|           ܕ@#       *                   �0@��+hF�?c           Ѝ@$       '                    @     P�?)             P@%       &                     �?���"͏�?            �B@������������������������       �ϊF�y�?             >@������������������������       �����>4�?             @(       )                     �?j�+$�j�?             ;@������������������������       ��n���?             "@������������������������       �����H�?	             2@+       .                    �?�gP�m�?:           Ћ@,       -                   �6@
�^���?�            �t@������������������������       ���C'7��?�            �r@������������������������       �2���h��?             C@/       0                    �?��M���?b           X�@������������������������       ��������?7            @U@������������������������       �V�4Na��?+           `}@2       5                   �0@��O��?           �{@3       4                    �?�;N��?             =@������������������������       �*D>��?             *@������������������������       �     ��?             0@6       9                    @a��"��?            z@7       8                    �?�CהOn�?�            �l@������������������������       ��(\����?             D@������������������������       �^�����?{            �g@:       ;                   �3@n�x����?r            �g@������������������������       �'޼��'�?.            �R@������������������������       ��x�V��?D            �\@=       Z                   �;@2�ʅ�S�?�           T�@>       K                   �9@����?�           h�@?       D                     @C"�R*��?           �}@@       C                    @�X��c��?�             u@A       B                    �?Q�d����?�            �s@������������������������       �!͎Z��?             E@������������������������       ���HVB�?�            0q@������������������������       �4և����?             5@E       H                    �?��e[��?X            `a@F       G                    �?�;��KM�?             C@������������������������       ������H�?             "@������������������������       �΃�\W�?             =@I       J                    �?��L�n��?<            @Y@������������������������       �`������?             7@������������������������       �A<:�&�?1            �S@L       S                    �?��ʻ��?�             q@M       P                    @}h����?D             \@N       O                    @��KL��?-            �R@������������������������       �n۶m۶�?#             L@������������������������       ������H�?
             2@Q       R                    �?�Q��X�?             C@������������������������       ��)O�?             2@������������������������       �>
ףp=�?             4@T       W                     �?33333��?o             d@U       V                    @�R�Gu�?>            �W@������������������������       ����i�?5            �T@������������������������       �UUUUUU�?	             (@X       Y                   �:@�,�F.�?1            �P@������������������������       �(+�>��?             ?@������������������������       ���yqY��?            �A@[       f                   �<@.��Q��?           �z@\       c                    @�Z�Gs3�?<            @X@]       `                    �?m��7�I�?.            �R@^       _                     �?     ��?             @@������������������������       �t�û��?             7@������������������������       ��2�tk~�?             "@a       b                    �?F?�!��?             E@������������������������       �l�l��?             >@������������������������       �UUUUUU�?             (@d       e                     �?�^|�!�?             7@������������������������       �����X�?             @������������������������       �     @�?             0@g       n                    �?f�j,���?�            pt@h       k                    �?'������?~            `g@i       j                    @	]Xt�?,            �Q@������������������������       ���e Ʊ�?            �E@������������������������       ��Cc}h��?             <@l       m                     �?Ĝ��?R             ]@������������������������       ��V�e�t�?             A@������������������������       ���"�x��?:            �T@o       r                    @�=�����?X            �a@p       q                   @@@C����?7            �U@������������������������       ��D��?'            �L@������������������������       �V4�ͫ�?             >@s       t                    @t������?!            �J@������������������������       �     ��?
             0@������������������������       ���0\K5�?            �B@�t�bh�h4h7K ��h9��R�(KKuKK��h��BxE       @|@      S@     �v@      @@      Q@      8@     �S@     ��@     ��@     �P@     @W@     �d@     ��@     �{@      (@      O@      J@     �`@     �L@     @v@      >@     �k@      (@      =@      @     �C@     @@     @~@      B@      L@     �W@     p{@     �p@      @      B@      2@     �U@      8@     �d@      (@     �V@      @      "@      �?      .@     ps@      q@      *@      6@      D@     `l@     @]@              "@      @      8@      @     �B@      �?      @                              @     �]@     �S@      �?      �?       @      P@      $@                               @              *@               @                                     �I@      @@              �?              3@      �?                                              @              �?                                      8@      7@              �?              .@      �?                                              @              �?                                      5@      "@              �?              $@                                                      �?                                                      @      ,@                              @      �?                                              @              �?                                      ;@      "@                              @                                                       @              �?                                      6@      @                              @                                                      @                                                      @      @                              �?                                                      8@      �?      @                              @      Q@      G@      �?               @     �F@      "@                               @              .@      �?       @                              @      M@      ?@                      @      ?@      @                               @              @              �?                                      @       @                       @      @       @                                               @      �?      �?                              @      K@      =@                      @      <@      @                               @              "@              @                                      $@      .@      �?              �?      ,@       @                                               @               @                                       @      @                      �?      (@      �?                                              @              �?                                       @       @      �?                       @      �?                                              `@      &@      U@      @      "@      �?      &@      h@     @h@      (@      5@      @@     `d@     �Z@              "@      @      6@      @     @X@      $@      M@      @      "@      �?       @     �U@     @\@      @      &@      >@     @Y@     �P@              @       @      1@      @     �I@      @      >@       @      @      �?      @     �O@      V@      �?      @      0@      J@     �F@              @       @      &@      @      A@      @      ,@       @      @      �?      @     �I@     @P@              @      &@      D@     �D@              @              &@      @      1@       @      0@              �?                      (@      7@      �?      �?      @      (@      @               @       @                      G@      @      <@       @      @              @      8@      9@      @      @      ,@     �H@      5@                              @             �D@      @      2@               @              @      ,@      0@      @      @      @     �@@      ,@                               @              @              $@       @      �?                      $@      "@               @       @      0@      @                              @              @@      �?      :@                              @     @Z@     @T@      @      $@       @      O@     �D@               @      �?      @      �?      ;@      �?      .@                                      V@     �S@      @      @       @      J@      >@              �?      �?      @      �?      @      �?      &@                                     �R@     �I@      @       @       @      A@      2@                      �?      @      �?      4@              @                                      ,@      ;@       @      @              2@      (@              �?              �?              @              &@                              @      1@      @       @      @              $@      &@              �?              �?              @               @                                       @                                       @       @                                              �?              @                              @      .@      @       @      @               @      @              �?              �?             �g@      2@     @`@       @      4@      @      8@     �g@     �j@      7@      A@     �K@     �j@      c@      @      ;@      .@      O@      3@      a@      $@     @T@      @      @              3@     �c@     �b@       @      4@     �A@     �a@     �X@              3@      ,@      F@      *@      (@              �?                                      9@      1@                              @       @                                              @              �?                                      @      .@                              @      �?                                              @              �?                                      @      .@                              @                                                      �?                                                       @                                      @      �?                                              @                                                      2@       @                              �?      �?                                              @                                                      @       @                                                                                       @                                                      ,@                                      �?      �?                                              _@      $@      T@      @      @              3@     ``@     �`@       @      4@     �A@     �`@      X@              3@      ,@      F@      *@      K@       @      0@              �?              "@     �O@      N@       @       @      "@      E@      G@              @       @      "@      @      H@      �?      ,@              �?               @     �N@      K@       @       @      "@      >@     �F@              @      �?      @      @      @      �?       @                              �?       @      @                              (@      �?              @      �?      @             �Q@       @      P@      @      @              $@      Q@     @R@      @      (@      :@     �V@      I@              *@      (@     �A@      @      @      �?      2@              @               @      @      @      @      �?      @      3@      @              �?              "@       @     �O@      @      G@      @      @               @      P@     �Q@      @      &@      3@      R@     �F@              (@      (@      :@      @      K@       @     �H@      @      *@      @      @     �@@      O@      .@      ,@      4@      R@      K@      @       @      �?      2@      @      "@      �?      �?                                      @      @                                      @                                               @      �?                                              �?      @                                                                                      �?              �?                                      @      @                                      @                                             �F@      @      H@      @      *@      @      @      ;@     �K@      .@      ,@      4@      R@     �H@      @       @      �?      2@      @      4@      @      7@              "@      @       @      7@     �B@      @      "@      @      G@      6@              @              @      @       @       @                       @                      @      *@      �?              �?       @      �?               @                      �?      2@       @      7@              @      @       @      0@      8@      @      "@      @      C@      5@              @              @      @      9@      @      9@      @      @      �?      @      @      2@       @      @      ,@      :@      ;@      @       @      �?      (@       @      @      �?      @      �?                                      &@      @      �?      @      "@      .@               @      �?      $@       @      2@       @      4@      @      @      �?      @      @      @      @      @       @      1@      (@      @                       @              X@      G@     �a@      4@     �C@      2@      D@     �R@      T@      >@     �B@     �Q@     �c@     �e@       @      :@      A@      G@     �@@      O@      >@      Y@       @      3@      @      =@     �P@      F@      (@      1@      B@     �\@      `@      @      .@      ,@      ?@      ,@      D@      5@     �Q@      @      @       @      6@     �E@      =@       @      .@      7@     �Q@     �V@      @      @      @      (@      @      =@      *@     �L@      @      @       @      (@     �C@      5@      @      (@      &@      J@      K@       @      @       @      &@      �?      =@      *@     �I@      @      @       @      (@      B@      5@      @       @      &@      G@      K@       @      @       @      $@      �?      @      @                                              @       @      �?      @      @      @      @               @               @      �?      :@       @     �I@      @      @       @      (@      ?@      3@      @      @       @      D@     �G@       @      �?       @       @                              @                                      @                      @              @                      �?              �?              &@       @      *@      @       @              $@      @       @      �?      @      (@      2@     �B@       @              @      �?       @      �?      @      @              �?               @      �?      @      �?               @      @      (@                      @               @              �?       @                                              @                              �?                              �?              �?      �?       @      �?              �?               @      �?              �?               @       @      (@                      @              �?      $@      @      $@      @      �?               @      @      @              @      $@      .@      9@       @                      �?              @      @      @       @                      @                                      �?      @      �?                                              @       @      @      �?      �?              @      @      @              @      "@      &@      8@       @                      �?              6@      "@      >@      �?      (@       @      @      7@      .@      @       @      *@     �F@     �B@      �?      &@       @      3@      &@      ,@      @      ,@      �?      @              @      (@      @              �?      @      3@      @              @      @      "@      @      "@       @      ,@              @                      @      @              �?      @      "@      @              @      @       @      �?       @      �?      ,@                                              @              �?      @      @      @              @      @      @      �?      �?      �?                      @                      @      @                               @                                      �?              @       @              �?      �?              @      @                                      $@      @              �?              �?      @      �?      �?              �?                                                                       @       @                              �?      @      @      �?                      �?              @      @                                       @       @              �?                               @      @      0@               @       @      @      &@       @      @      �?      "@      :@      >@      �?      @      @      $@      @      @      @      &@              @      �?      �?      @      @      @      �?      @      6@      (@      �?      @       @      @              @      @      "@              @      �?      �?      @      @      @      �?      @      6@      $@      �?      @       @      @                               @                                      @      �?                       @               @              �?                              @      �?      @              @      �?      @      @      �?      �?              @      @      2@              @       @      @      @                      @              �?              �?      @                              @      @      @              @       @      @      @      @      �?       @              @      �?       @              �?      �?              �?      �?      ,@                               @      @      A@      0@     �E@      (@      4@      ,@      &@      "@      B@      2@      4@     �A@      F@      F@      @      &@      4@      .@      3@      @      @      @      @       @       @      �?      @      *@       @      @      @      0@      "@              �?      @      �?      "@      @      @      @      @       @       @      �?              $@      �?      @      @       @       @              �?      @      �?       @       @      @      @                              �?              @               @      @       @      @                                       @       @      @                                                      @               @      @              @                                       @                      @                              �?               @                               @      �?                                              @              �?      @       @       @                      @      �?      �?      @      @      @              �?      @      �?      @      @                      @       @       @                                      �?       @      @      @              �?              �?      @                      �?                                              @      �?              �?              �?                      @              �?                               @                              @      @      �?       @               @      �?                       @              �?                                                                      �?      �?                      �?      �?                       @              �?                               @                              @       @               @              @                                                      <@      &@     �C@      @      2@      (@      $@      @      7@      0@      .@      <@      <@     �A@      @      $@      ,@      ,@      $@      "@       @      :@      @      $@       @      $@      @      $@      "@      (@      0@      &@      ,@       @      @      *@      @       @      @      @       @              @              @       @      @      @      @      @      "@       @      �?       @       @      �?       @      @      @      @              �?              �?              @      @      @       @       @       @               @              �?      �?                      @               @              @       @      @                      @      @              �?               @              �?      @       @      2@      @      @       @      @      @      @      @       @      $@       @      @      �?      @      &@      @      @      �?       @      @              @      @      �?                              @      @                              @       @      �?      �?      @              *@      @      @      @      @      @      @      @      @      @       @      @      �?              "@       @      @      3@      @      *@       @       @      @              �?      *@      @      @      (@      1@      5@      �?      @      �?      $@       @      (@      @       @       @              @              �?      @      @      @      (@      (@      &@      �?       @      �?      @              @       @      @       @               @              �?      @      @      @      @      @      $@      �?      �?      �?      @              "@      �?      �?                       @                               @              @      @      �?              �?                              @              @               @                              $@                              @      $@              �?              @       @                      @              @                              @                               @      �?                                              @               @              @                              @                              @      "@              �?              @       @�t�bub��     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�5hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKuhnh4h7K ��h9��R�(KKu��hu�B�         <                   �5@]���.��?�	           ��@                           �?V,��b��?A           ��@                           @��]�ֲ�?�           0�@                           �?a�0�U�?'            }@                          �1@���Q��?�            �s@                          �0@�?P����?.            �Q@������������������������       �Dy�5��?             3@������������������������       �Jw���+�?            �I@	       
                     �?f"����?�            �n@������������������������       ��b� I`�?*            �Q@������������������������       �' )x L�?l            �e@                          �3@G<�A+K�?c             c@                           @�H�/��?@            �Y@������������������������       ���"c��?4            �S@������������������������       ��q�q�?             8@                          �4@(~��k	�?#             I@������������������������       �     ��?             @@������������������������       ��q�q�?             2@                           @��=$m��?Z           Ё@                           @�"�n��?>           X�@                           �?�Ҕ|���?�            @w@������������������������       �Ǥf~��?c            �d@������������������������       �g\���?�             j@                           @I��t��?V            �b@������������������������       ��7�A�?0             V@������������������������       �~VC�1��?&            �O@                          �2@��I�J�?            �G@������������������������       ��d��E�?             1@                            �?��2Tv�?             >@������������������������       ��(\����?             $@������������������������       ���(\���?
             4@        -                    �?r���?�           ��@!       (                    �?���2M��?           �{@"       %                     �?2 �a�?[            `b@#       $                    �?�q�q��?             H@������������������������       �      �?
             0@������������������������       �     p�?             @@&       '                   �4@�9�� ��??            �X@������������������������       �[����1�?1            @S@������������������������       ��Z=;n�?             6@)       *                   �0@7�[\�s�?�            `r@������������������������       �����>4�?             ,@+       ,                    @����v�?�            �q@������������������������       �ɖٍi��?M            �^@������������������������       �s������?e            �c@.       5                     �?è�b�]�?�           (�@/       2                   �3@o�y{�e�?�            0x@0       1                    @ء����?�             k@������������������������       ��ޖ	�?�            �h@������������������������       ��u]�u]�?             5@3       4                    �?����?a            @e@������������������������       ��Ezu��?#             O@������������������������       �@�9S˅�?>             [@6       9                   �0@T�s���?�             p@7       8                     @�ങa�?             ?@������������������������       �      �?
             ,@������������������������       ��&5D�?
             1@:       ;                     @/��r�?�            `l@������������������������       ���3L��?N             [@������������������������       �p���-�?W            �]@=       \                   �9@��2>�?a           ��@>       M                    �?lB� ��?�           �@?       F                   �7@i��{�$�?            `|@@       C                    �?jq�%���?�             q@A       B                     @����`��?:            @V@������������������������       ���_Ou�?.            �Q@������������������������       �x�5?,R�?             2@D       E                    @��m{��?q             g@������������������������       ��l����?.            �S@������������������������       �����?C            �Z@G       J                     �?�M�)���?u            �f@H       I                   �8@-s�["�?             G@������������������������       ����y4F�?             3@������������������������       �#����?             ;@K       L                   �8@Ԁ�C`(�?Y            �`@������������������������       �T��Z���?5            @T@������������������������       � ���]�?$            �J@N       U                     @����?p           ��@O       R                    @�,����?�            Px@P       Q                   �8@?��H���?�            �l@������������������������       �t�@��?u            �f@������������������������       ��8��8N�?             H@S       T                     �?b�����?l             d@������������������������       �~Ց�X��?(            �M@������������������������       ��������?D            �Y@V       Y                    @P��P;��?t            @g@W       X                   �7@������?-            @R@������������������������       �o,x���?            �C@������������������������       ��0�!��?             A@Z       [                    @�m�S��?G            @\@������������������������       ��2�o�U�?%            �K@������������������������       �� �f>�?"             M@]       l                    �?�\gh��?�           Ї@^       e                    �?eIG����?�             {@_       b                     �?��"��?`            �c@`       a                     �?����?3            @V@������������������������       �.�T�6�?             J@������������������������       ���0\K5�?            �B@c       d                    @G>&���?-            �Q@������������������������       �ΎZ��5�?             E@������������������������       �$I�$I��?             <@f       i                    @l�����?�            q@g       h                   �>@�I�b�?A            @\@������������������������       �W�q����?5            @V@������������������������       ��8��8��?             8@j       k                     �?\���(\�?]             d@������������������������       �����n�?#            @P@������������������������       �R>��\��?:            �W@m       t                   @A@3�����?�            �t@n       q                    @��J����?�            Ps@o       p                    @�a�z��?}            �i@������������������������       ��X���B�?n            �e@������������������������       �rH��7�?             =@r       s                    �?_������?I            @Z@������������������������       ��fG-B��?             5@������������������������       �����S�?8             U@������������������������       �P&�to@�?             5@�t�bh�h4h7K ��h9��R�(KKuKK��h��BxE       pz@      T@     @t@      ?@     �O@      7@     @W@     x�@     ��@      N@     @V@     �e@     H�@     @{@      $@     �P@      M@     @b@      L@     �p@      1@      c@      @      *@      �?     �B@     �{@      y@      3@     �A@     �U@     `v@      g@              ,@      "@      P@      3@     @\@      @      L@      �?      �?              0@     �p@     �k@       @      ,@      9@     `f@     @T@              $@       @      <@      @      N@      @      8@                              @      V@     �Y@       @      @      1@     �T@     �C@               @              5@      @     �F@      �?      5@                              @     �L@      M@       @      @      @     �L@      ;@               @              *@      @      &@              @                                      :@      *@       @               @       @      @                                               @                                                      @      @                              @      �?                                              "@              @                                      3@       @       @               @      @      @                                              A@      �?      2@                              @      ?@     �F@              @      @     �H@      6@               @              *@      @      $@      �?      @                                      @      0@               @      @      <@      �?                                      �?      8@              .@                              @      9@      =@              @       @      5@      5@               @              *@      @      .@       @      @                                      ?@      F@              �?      $@      :@      (@                               @               @              @                                      ;@      ;@              �?      $@      .@      @                              @               @              @                                      :@      *@              �?      @      *@      @                              @                                                                      �?      ,@                      @       @                                      @              @       @                                              @      1@                              &@       @                              �?              @                                                      @      *@                              @      @                              �?               @       @                                              �?      @                               @      �?                                             �J@      @      @@      �?      �?              $@     �f@     �]@      @      @       @      X@      E@               @       @      @             �H@      @      >@      �?      �?               @     �d@     @]@      @      @       @     �T@     �D@               @       @      @             �A@       @      0@      �?                       @      a@     �T@      �?      @      @      K@      6@                       @      @              @       @      @                              �?      R@      C@               @      @      <@       @                                              <@              $@      �?                      �?     @P@      F@      �?      @      �?      :@      4@                       @      @              ,@      �?      ,@              �?                      >@     �A@       @      �?      �?      =@      3@               @               @              @              @                                      &@      5@              �?      �?      4@      2@                               @              @      �?      @              �?                      3@      ,@       @                      "@      �?               @                              @               @                               @      ,@       @      @                      *@      �?                                               @                                                      &@       @                               @                                                       @               @                               @      @              @                      &@      �?                                              �?               @                               @                      @                       @                                                      �?                                              @      @                                      "@      �?                                              c@      &@     @X@      @      (@      �?      5@     `e@     �f@      &@      5@      O@     `f@      Z@              @      @      B@      *@      M@      @     �J@       @      "@      �?      @     �E@     �L@      $@      0@      @@      P@      H@              �?      �?      9@      @      8@      @      &@              @      �?      @      0@      >@       @      &@       @      ,@      $@                      �?       @              $@              @                              @      �?      1@               @       @      @       @                              �?               @              @                              @      �?       @                               @                                      �?               @                                              �?              .@               @       @       @       @                                              ,@      @      @              @      �?              .@      *@       @      "@      @      $@       @                      �?      �?              &@      @      @              @                      .@      &@              @       @      @      @                              �?              @              �?               @      �?                       @       @       @      @      @      �?                      �?                      A@      �?      E@       @       @              @      ;@      ;@       @      @      8@      I@      C@              �?              7@      @      @              �?                                       @      �?                              �?       @                                              ;@      �?     �D@       @       @              @      9@      :@       @      @      8@     �H@      B@              �?              7@      @      *@      �?      2@       @       @              �?      @      "@      @      �?      @     �A@      6@                              @              ,@              7@                               @      3@      1@      @      @      3@      ,@      ,@              �?              2@      @     �W@      @      F@      �?      @              ,@      `@      _@      �?      @      >@     �\@      L@              @      @      &@      @     �M@       @      5@               @              @      P@     �T@      �?      @      6@     @Q@     �A@              @      @      @      @      @@       @       @                              @     �E@     �H@      �?       @      @      F@      &@              @      @      @      @      ?@       @       @                              @      D@      D@      �?       @      @     �C@      &@              @      @      @      @      �?                                              �?      @      "@                      �?      @                                      �?              ;@              *@               @              @      5@      A@              �?      0@      9@      8@                       @      �?      �?      �?                              �?                      *@      3@                      @      "@      .@                                              :@              *@              �?              @       @      .@              �?      (@      0@      "@                       @      �?      �?     �A@       @      7@      �?      �?              @      P@     �D@               @       @      G@      5@                              @       @                      �?              �?                      3@      @                              @      �?                                                                                                      "@                                      @      �?                                                              �?              �?                      $@      @                               @                                                     �A@       @      6@      �?                      @     �F@      C@               @       @      D@      4@                              @       @      2@              @                               @      >@      4@                              5@      "@                              �?      �?      1@       @      0@      �?                      @      .@      2@               @       @      3@      &@                              @      �?     �c@     �O@     `e@      ;@      I@      6@      L@     �]@     �i@     �D@      K@     @U@     0p@     `o@      $@      J@     �H@     �T@     �B@     �Z@      9@     @Z@      $@      5@      (@      ?@     �U@     �b@      4@     �@@      D@     �b@     �c@      @      0@      ;@      ;@       @      F@       @     �H@              @      @      $@     �E@      V@       @      $@      .@      O@     �S@              @      2@      @      @      ?@      @      =@              @      @      �?      :@     �H@       @      @       @      J@     �C@              @      (@      @              1@      �?      0@               @              �?       @      4@       @      �?      @      .@      "@                                              "@      �?      .@              �?              �?       @      4@       @      �?      @      &@      @                                               @              �?              �?                                                              @      @                                              ,@      @      *@              @      @              8@      =@              @      @     �B@      >@              @      (@      @              @              @                      @              $@       @              �?      �?      .@      ,@              @      (@                      @      @      "@              @      �?              ,@      5@               @      @      6@      0@                              @              *@      @      4@                              "@      1@     �C@              @      @      $@     �C@              @      @      @      @      @      �?       @                              @      �?      (@              �?               @      0@                              @              �?      �?      �?                                      �?      @                                      $@                              �?               @              �?                              @               @              �?               @      @                               @              $@      @      2@                              @      0@      ;@              @      @       @      7@              @      @      �?      @      @      �?      *@                              @      *@      1@               @       @       @      ,@              �?      @              @      @       @      @                                      @      $@              @      @      @      "@               @      @      �?              O@      1@      L@      $@      ,@       @      5@     �E@      O@      2@      7@      9@     @V@     �S@      @      $@      "@      4@      @      J@      "@      B@      @      @      @      1@      =@      A@      0@      2@      2@     �R@      E@      �?      $@      @      .@       @      E@      @      8@      @      �?      @      @      8@      8@      @      @      &@      B@      7@              @      �?      "@      �?     �C@      @      1@      @      �?              �?      2@      7@      @       @      &@      ;@      4@              @      �?      @      �?      @      �?      @                      @      @      @      �?      �?      @              "@      @                              @              $@      @      (@       @       @              $@      @      $@      $@      *@      @      C@      3@      �?      @      @      @      �?      @      @      @       @                      @      @      �?              "@      �?      0@      @              @       @      �?      �?      @      �?      "@               @              @       @      "@      $@      @      @      6@      ,@      �?       @       @      @              $@       @      4@      @      &@      @      @      ,@      <@       @      @      @      .@     �B@      @              @      @      @      @      @       @      @      @      @       @      �?      5@      �?       @      @      @       @                      @      @       @              �?                      @      @              �?      *@      �?       @      �?      @                               @      @       @      @       @       @      @                       @               @                       @      �?       @                      �?                      @      @      2@      �?      @       @       @      *@      @      �?      @      @      $@      =@      @              �?       @      �?      @      @      @              @       @              @      @      �?      �?      @      @      1@       @                                      �?       @      .@      �?       @               @      "@      @               @              @      (@      �?              �?       @      �?      J@      C@     �P@      1@      =@      $@      9@     �@@     �K@      5@      5@     �F@      [@     �W@      @      B@      6@     �K@      =@      <@      6@      B@      0@      6@       @      3@      @      B@      @      1@      >@     �I@      E@      @      9@      0@      9@      6@      5@      .@      .@      @      @              "@      @      0@       @       @       @      =@      ,@              @      @      @      @      "@      *@      @       @                      @      @      &@       @      �?      �?      &@       @              �?      @      @      @      @      @               @                      @               @       @                      &@      @              �?      @      @      @       @      $@      @                               @      @      @              �?      �?              @                      �?      �?      �?      (@       @       @      �?      @              @              @              �?      �?      2@      @              @       @              �?      $@      �?       @              �?                              @              �?      �?      @      @              @      �?                       @      �?              �?      @              @               @                              (@      �?                      �?              �?      @      @      5@      *@      1@       @      $@       @      4@      @      .@      <@      6@      <@      @      3@      $@      3@      1@      �?      �?      @      "@      (@       @      @       @      "@      �?      �?      @      @       @       @      @      @      2@      $@      �?      �?      @      "@      "@      �?      @       @      "@                       @      @      @               @      @      2@      @                      �?              @      �?                              �?      �?      @              @       @      @      @              @      @      @      ,@      @      @      @      @              &@      @      ,@      7@      .@      4@      @      ,@      @      �?      @      @       @              �?       @       @       @              @      �?      "@      @      &@      @              $@                      �?       @      @      ,@      @      @      @       @              @      @      @      1@      @      *@      @      @      @      �?      @      8@      0@      >@      �?      @       @      @      <@      3@      ,@      @      .@     �L@      J@      �?      &@      @      >@      @      8@      ,@      ;@      �?      @       @      @      <@      3@      &@      @      ,@     �L@      F@      �?      $@      @      <@      @      .@      @      &@      �?      @       @      @      6@      ,@      $@       @      @      E@      =@      �?       @       @      7@      @      *@      @       @      �?      @       @       @      3@      $@       @       @      @      E@      9@      �?      @       @      1@      @       @              @              @              �?      @      @       @                              @              �?              @              "@      &@      0@              �?               @      @      @      �?       @      @      .@      .@               @      @      @      @      �?      @                      �?                       @      @                       @      �?       @              �?              �?               @      @      0@                               @      @      �?      �?       @      @      ,@      *@              �?      @      @      @               @      @                              �?                      @              �?               @              �?               @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ,�BhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         <                    �?h瘳�?�	           ��@                          �2@BTaU*�?           ��@                          �1@P�C��?�            �t@       	                    �?�1�Lz�?x            �f@                          �0@|��U�=�?-            �P@������������������������       �ݾ�z�<�?             *@                           @y��G'�?"            �J@������������������������       �      �?             8@������������������������       �@�"s�?             =@
                           �?��0RZV�?K            �\@                            �?s
^N���?             E@������������������������       �*L�9��?             &@������������������������       ������?             ?@                          �0@ʛE��}�?3            @R@������������������������       ��nkK�?             7@������������������������       ���q���?&             I@                           �?�짮���?\            �b@                           �?Hk�����?%            �I@                           @�������?             9@������������������������       �      �?             0@������������������������       �0�����?             "@                           �?��?��?             :@������������������������       �      �?              @������������������������       �Lh/����?             2@                           �?�43&���?7            @X@                           @�m(�9W�?            �E@������������������������       �_B{	�%�?             2@������������������������       �a��+e�?             9@                           @82Y�Qo�?!             K@������������������������       �h�T�B�?            �D@������������������������       �؉�؉��?             *@        /                   �=@�PsMT�?1           ��@!       (                    �?�qXn	�?�           p�@"       %                     �?��r��e�?           0{@#       $                   �3@<��wZ�?R            ``@������������������������       ��q�q�?             (@������������������������       ��	�0�?J            �]@&       '                   �<@^Cy��?�             s@������������������������       �x�b���?�            �q@������������������������       �4%���?
             1@)       ,                     �?+�%m�P�?�           H�@*       +                    �?��4eQ^�?�            �t@������������������������       ��3�9A��?O            @_@������������������������       �Y�Cc�?�            @j@-       .                   �3@�V���?�            �y@������������������������       ���(��(�?             E@������������������������       �v=q��?�             w@0       7                   �@@/`1��?W             a@1       4                    �?�טb���?>            �Y@2       3                   �>@>��^�?             ?@������������������������       �      �?	             (@������������������������       �"P7��?
             3@5       6                    �?ݚ)�?+             R@������������������������       ����Q��?             7@������������������������       �p*�o��?            �H@8       ;                   �A@�.k���?             A@9       :                     @�8��8��?             8@������������������������       �9��8���?	             (@������������������������       �r�q��?	             (@������������������������       �ffffff�?             $@=       X                   �3@܀b��?�           ��@>       K                     @174`?�?I           �@?       D                   �0@*���?�           �@@       C                    @�����R�?U            �`@A       B                    �?��W!�r�?I            �[@������������������������       ���Ӡy��?-            @Q@������������������������       ���&q	��?            �D@������������������������       �����!p�?             6@E       H                   �1@8�V�4�?�           �@F       G                    @��z>׬�?�            �k@������������������������       ��������?|            @j@������������������������       �"���c��?             *@I       J                     �?�I
F�m�?�            �w@������������������������       ���lW+��?�            �p@������������������������       �Ô�*��?M            �\@L       Q                    �?�8��8J�?s             h@M       P                    @����o�?4             W@N       O                    @o�Z<�?)            �R@������������������������       ���Xh��?            �K@������������������������       �{�G�z�?             4@������������������������       ��?�0�!�?             1@R       U                    �?��3���??             Y@S       T                    @�W+J���?            �G@������������������������       ���/��@�?             7@������������������������       ���8��8�?             8@V       W                    @��R�:��?$            �J@������������������������       ��)F�?            �F@������������������������       �      �?              @Y       h                   �;@�L��?^           �@Z       a                    @r#��U��?�           ̑@[       ^                    �?�����b�?�           \�@\       ]                    @~I+��?J           �~@������������������������       �v�����?�            �p@������������������������       ��M�j�e�?�            �k@_       `                   �7@�9����?b           p�@������������������������       �Z�n����?�            �x@������������������������       ��(%LL��?p            �d@b       e                    @]@˜���?:             W@c       d                    @�,y8"q�?            �B@������������������������       ��Q����?             4@������������������������       �U��6���?	             1@f       g                     �?�>��6��?!            �K@������������������������       �q=
ףp�?             4@������������������������       �{�X�o�?            �A@i       p                    �?ظ�, u�?x            �h@j       m                    @���%�?#             J@k       l                     �?tk�
��?             =@������������������������       ��>4և��?             ,@������������������������       ���2Tv�?
             .@n       o                     �?J��LQ�?             7@������������������������       ���!pc�?             &@������������������������       �9��8���?             (@q       t                     �?}A(�x�?U            `b@r       s                    @(x��:�?            �D@������������������������       ��;��KM�?             3@������������������������       ��Ra����?             6@u       v                   @A@Y��l�6�?>            �Z@������������������������       ��)�w�?�?5            @V@������������������������       �/k��\�?	             1@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       }@     �V@     0u@     �@@     �Q@      :@     @W@      �@     ��@     �S@     �V@     @e@     �@     Py@      *@     �Q@     �K@     �`@      N@     �i@     �C@     @d@      (@     �C@      5@      G@     �_@     @g@     �C@     �I@     �W@      n@      g@      @     �B@      A@     @S@      G@      L@      �?      9@      �?      �?              @     �P@     �F@      @      @      "@     �K@      C@               @      �?       @       @      D@      �?      (@              �?              @      E@      2@      @      �?      @      :@      7@              �?      �?      �?       @      *@              @                                      8@      @       @              �?      @      @                                              �?              @                                      @       @                              �?      �?                                              (@              @                                      3@      @       @              �?      @      @                                              @                                                      @       @       @              �?      @      @                                              "@              @                                      (@      @                              �?                                                      ;@      �?      @              �?              @      2@      &@       @      �?      @      4@      1@              �?      �?      �?       @      *@                                                      "@      @       @              @      @       @                              �?              �?                                                      @       @                      @      �?                                                      (@                                                      @      @       @                      @       @                              �?              ,@      �?      @              �?              @      "@      @              �?      �?      *@      .@              �?      �?               @      (@      �?      �?                                      �?      �?                               @      @                                               @              @              �?              @       @      @              �?      �?      &@      $@              �?      �?               @      0@              *@      �?                      @      8@      ;@      @      @      @      =@      .@              �?              @               @              @                                      @      &@              @              &@       @              �?               @               @               @                                      @       @               @              "@      �?              �?              �?               @                                                      @      �?                              @      �?              �?                                               @                                      �?      �?               @               @                                      �?              @              @                                      �?      "@              �?               @      �?                              �?              @                                                      �?      �?                              �?                                      �?               @              @                                               @              �?              �?      �?                                               @              @      �?                      @      2@      0@      @      �?      @      2@      *@                              @              @              �?                              @      *@      @                      @       @      �?                              @              �?              �?                              @      $@                                      �?      �?                                               @                                                      @      @                      @      @                                      @              @              @      �?                              @      "@      @      �?      �?      $@      (@                               @               @              @      �?                               @       @      @      �?      �?      @      $@                               @              @                                                      @      �?                              @       @                                             �b@      C@      a@      &@      C@      5@     �C@      N@     �a@      @@      G@     @U@     @g@     @b@      @     �A@     �@@     @Q@      F@     `a@     �B@      _@      @      :@      *@      @@     �M@      a@      <@      B@     �R@      g@      a@       @      >@      9@      L@      A@      L@       @     �@@      �?      "@      �?      $@      >@      M@      ,@      $@      2@     �W@     �I@               @      @      *@      0@      &@      @      @      �?      @      �?      �?      @      2@              �?      @     �G@      *@                      �?      @      @       @       @                                                                              �?      @      @                                              "@      @      @      �?      @      �?      �?      @      2@              �?      @      F@      "@                      �?      @      @     �F@      @      <@              @              "@      :@      D@      ,@      "@      *@     �G@      C@               @      @      @      "@      F@      @      6@              @              @      :@      C@      *@      "@      *@     �G@      B@               @      @      @       @      �?              @                               @               @      �?                               @                               @      �?     �T@      =@     �V@      @      1@      (@      6@      =@     �S@      ,@      :@     �L@     �V@     �U@       @      6@      4@     �E@      2@     �A@      "@     �F@       @      @              $@      6@      ;@      "@      2@      6@     �B@      A@      �?      (@       @      =@      "@      $@      �?      2@              �?              @       @      *@              "@      @      9@      $@                      @      "@      @      9@       @      ;@       @      @              @      ,@      ,@      "@      "@      1@      (@      8@      �?      (@       @      4@      @      H@      4@      G@      @      &@      (@      (@      @     �I@      @       @     �A@     �J@      J@      �?      $@      (@      ,@      "@               @      @                                      �?       @      �?              @      *@      @                              @              H@      2@      E@      @      &@      (@      (@      @     �E@      @       @      @@      D@     �H@      �?      $@      (@      @      "@      $@      �?      *@      @      (@       @      @      �?      @      @      $@      $@       @      "@      @      @       @      *@      $@      $@      �?      &@      @      @       @      @      �?      @      �?       @      @       @      "@              @      @      (@      @      @                               @               @      �?      @                      @       @      @                       @       @       @                                      �?               @      �?      �?                      �?      �?      �?                       @               @      @                              �?                               @                      @      �?      @                               @              @      �?      &@      @      @       @      @              �?      �?       @                      @              @      @      $@      @      @               @      �?      �?       @      �?                                                       @                       @       @              �?      �?      "@      @       @      @      @              �?      �?       @                       @              @      @       @      @                       @              @              �?              �?      @       @      @                      @       @      �?      �?      @                       @               @                                      @      �?      @                      @       @              �?      @                       @                                                      @      �?      @                              �?              �?                                               @                                                                              @      �?                      @                                      @              �?              �?              �?      �?                                      �?                     @p@     �I@      f@      5@      @@      @     �G@      z@     �y@     �C@     �C@      S@      u@     �k@      @      A@      5@      M@      ,@     �[@      "@      M@       @      @              ,@      q@     �i@      @      @      9@     �`@     @P@              "@      @      @      @     �T@      @      ?@               @              $@     �l@     �e@      @      @      5@     �Z@     �G@              @      @      @      �?      6@              @                                      J@      B@              �?       @      .@                                      �?              $@              @                                     �H@      >@              �?       @      ,@                                      �?              @              �?                                     �A@      3@              �?               @                                                      @               @                                      ,@      &@                       @      @                                      �?              (@                                                      @      @                              �?                                                     �N@      @      <@               @              $@      f@     `a@      @      @      3@     �V@     �G@              @      @      @      �?      3@       @       @                              @      Q@     �I@              �?      $@     �E@      ,@                               @              3@       @       @                              @      N@      I@              �?       @      E@      *@                               @                                                                       @      �?                       @      �?      �?                                              E@      @      4@               @              @     @[@      V@      @      @      "@      H@     �@@              @      @      @      �?     �@@      @      *@                              @     @S@     �H@      �?      @       @      A@      <@              @      @      �?      �?      "@              @               @                      @@     �C@       @              �?      ,@      @                              @              ;@       @      ;@       @      �?              @     �E@      ?@              �?      @      <@      2@               @                       @      .@              "@                               @      >@      $@                      �?      4@      @                                              ,@              @                                      =@      @                      �?      .@       @                                               @              @                                      7@      @                      �?      .@                                                      @              @                                      @      @                                       @                                              �?               @                               @      �?      @                              @      @                                              (@       @      2@       @      �?               @      *@      5@              �?      @       @      *@               @                       @       @              "@      �?                       @      @      @              �?       @      @      "@               @                              @              @      �?                              �?      @              �?       @       @      �?                                              @              @                               @       @                                      �?       @               @                              @       @      "@      �?      �?                      $@      ,@                      �?      @      @                                       @      @       @      "@      �?      �?                      "@       @                      �?      @      @                                       @                                                              �?      @                              �?                                                     �b@      E@     �]@      3@      =@      @     �@@     @b@     �i@      B@     �@@     �I@     �i@     �c@      @      9@      2@     �I@      &@     �`@      7@     �Y@      .@      1@      @      ?@     @a@      h@      7@      >@      B@     `f@     ``@       @      5@      (@      C@      $@     @^@      7@     �U@      &@      &@      @      5@      `@     �g@      6@      :@     �A@     �d@     �_@       @      5@      $@      @@      $@      H@      $@      C@      @       @      �?      @     @P@      \@      "@      .@      *@      U@     �O@              @      @      *@       @      <@      $@      <@      @              �?      @      <@     �N@      @      @      "@      H@      @@               @      �?      @      �?      4@              $@               @                     �B@     �I@      @      &@      @      B@      ?@               @       @      @      �?     @R@      *@     �H@       @      "@      @      1@     �O@     �S@      *@      &@      6@     �T@     �O@       @      1@      @      3@       @      M@       @      <@      @      @              $@     �G@     �G@      @      @      2@      P@      J@              *@      @      ,@      @      .@      @      5@      @      @      @      @      0@      @@      @      @      @      2@      &@       @      @              @      �?      *@              .@      @      @              $@      $@       @      �?      @      �?      *@      @                       @      @              @              @      @                      @      @              �?      @      �?      �?      �?                                              @              �?                              @      @                      @      �?      �?                                                      @              @      @                      �?      �?              �?                              �?                                              @               @              @              @      @       @                              (@      @                       @      @              @              @                                      �?       @                               @       @                       @                       @              �?              @              @      @                                      $@       @                              @              0@      3@      1@      @      (@      �?       @       @      &@      *@      @      .@      9@      9@      @      @      @      *@      �?      �?       @      �?      �?                                      @       @       @      @      $@      @              �?              @      �?      �?              �?      �?                                       @       @       @      @      @      �?              �?              @                              �?                                               @       @      �?      �?      @      �?                               @              �?                      �?                                                      �?      @      @                      �?               @                       @                                                      @                              @      @                              �?      �?                                                                      @                               @      @                                                       @                                                                                      �?      �?                              �?      �?      .@      &@      0@      @      (@      �?       @       @      @      &@      �?       @      .@      2@      @      @      @       @                      @      @              @                      @      �?       @              @              "@               @      @      �?                      @      @                                      �?                              @               @               @      @      �?                               @              @                      @      �?       @                              @                       @                      .@      @      &@      @       @      �?       @      @      @      "@      �?      @      .@      "@      @      �?      �?      @              "@      @       @      @       @      �?       @      @      @      @      �?      @      .@      "@      @      �?      �?      @              @       @      @                                                      @               @                                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��)hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKehnh4h7K ��h9��R�(KKe��hu�B         8                     @��__&��?�	           ��@                           �?	 `j�?�           �@                          �1@?[����?)           �@                           @�DQ:q��?�             n@                           �?�q�?�            �l@                          �0@ϊF��?K             ^@������������������������       ������t�?            �G@������������������������       �
a\�CZ�?,            @R@	       
                    @:�G���?J            �[@������������������������       �p=
ףp�?             D@������������������������       ��!�`�u�?.            �Q@������������������������       �ffffff�?             $@                           @�1�	��?�           (�@                           �?    �V�??            �@                            �?�9�Q�a�?o            �f@������������������������       ��y�#�?*            �O@������������������������       �(}�'}��?E             ^@                          �5@��	z�?�            �t@������������������������       �     �?S             `@������������������������       ��R����?}             i@                          �=@�d"@��?M           P�@                          �8@-�����?B           �@������������������������       � n[�"^�?           �z@������������������������       ���W�3�?2             S@������������������������       ����[���?             2@       )                    �?.*!���?�           �@       "                    @}�v��?           �y@                          �9@�����B�?�             i@                            �?Yc���?o            �c@������������������������       ���^B{	�?1             R@������������������������       �������?>            �U@        !                   �:@ĭ[F�?            �D@������������������������       �~h����?             ,@������������������������       ��L-���?             ;@#       &                    @-֓��|�?�            �j@$       %                     �?X�<ݚ�?c             b@������������������������       ��i��i��?;             U@������������������������       �""""""�?(             N@'       (                     �?��=�/�?,            @Q@������������������������       �9�>� ��?!            �H@������������������������       ����(\��?             4@*       1                   �3@lk}�?�           P�@+       .                     �?_<X�μ�?�             u@,       -                    @�D����?�            �o@������������������������       ���T��?P             ]@������������������������       �I�9߄�?Y             a@/       0                    @����>4�?2             U@������������������������       �r-�T��?             :@������������������������       ����6��?#             M@2       5                   �>@&jā�h�?�           Є@3       4                   �9@��	O�?�           �@������������������������       �P:���?           �z@������������������������       ��@�mM`�?r             g@6       7                    @cT!)��?$            �L@������������������������       ��h$���?             .@������������������������       ������?             E@9       J                    �?��f[��?            �@:       ;                   �0@&���1�?�           @�@������������������������       � �P|��?             ;@<       C                    �?�*�4�?�           h�@=       @                    �?-�N����?�            �q@>       ?                    �?�U�����?4            �P@������������������������       ���M[�?             ;@������������������������       �      �?             D@A       B                    �?�ӇA��?�            `k@������������������������       �*�%q��?!            �K@������������������������       �B�b�?b            �d@D       G                    �?�zZ�@�?           �z@E       F                   �9@^������?I             [@������������������������       ��gB����?@            �W@������������������������       �I�$I�$�?	             ,@H       I                    �?Ћ~,*�?�            0t@������������������������       ��閮�h�?3            �U@������������������������       �z��_��?�            �m@K       Z                    @O%�DI�?,           �}@L       S                    @�������?�            �u@M       P                   �5@:㨾��?n            `f@N       O                   �1@     >�?P             `@������������������������       �=;n,��?             F@������������������������       ��U̠ç�?2             U@Q       R                    @ *4>HR�?            �I@������������������������       �Y2���h�?             C@������������������������       ��]�`��?             *@T       W                    @Q]NR'�?t            �e@U       V                    �?$B`~���?$            �I@������������������������       �      �?             <@������������������������       �K����?             7@X       Y                   �5@���9d\�?P            @^@������������������������       �`����x�?&             M@������������������������       ����h%��?*            �O@[       `                   �5@     ��?J             `@\       _                   �4@��ڬ���?*            �S@]       ^                   �0@~]y�Q��?#            @P@������������������������       ��9����?             &@������������������������       �Ĺ��3�?             K@������������������������       �ݾ�z�<�?             *@a       b                   �6@	�c��?              I@������������������������       ��Cc}�?	             ,@c       d                    @Lh/����?             B@������������������������       ��h$���?	             .@������������������������       �lv�"��?             5@�t�bh�h4h7K ��h9��R�(KKeKK��h��B�;       �y@      W@     `u@     �A@     �S@      7@     �S@     x�@     �@     �M@      W@     �e@     ��@     |@      2@      P@     �K@      e@      E@     Pq@     �L@     �k@      3@     �E@      @      L@     �z@      }@      E@      N@     @]@     y@     �q@       @     �C@      C@     @[@      :@     �a@      :@      U@      �?      *@              3@     �n@     �p@      1@      >@     �@@     �i@     ``@              $@      $@      >@      $@      >@       @      @                              @     �Y@     �J@               @      @      A@       @                                              ;@       @      @                              @     �X@     �J@               @       @      @@       @                                              .@       @      �?                                     �I@      5@               @       @      4@      @                                              @              �?                                      =@       @               @              @                                                      &@       @                                              6@      *@                       @      1@      @                                              (@               @                              @     �G@      @@                              (@       @                                              @              �?                                      *@      2@                              @                                                      @              �?                              @      A@      ,@                              "@       @                                              @                                                      @                              �?       @                                                     �[@      8@     @T@      �?      *@              .@      b@     �j@      1@      <@      >@     �e@     �^@              $@      $@      >@      $@     �L@      .@     �K@              @              $@     �B@     �U@      @      .@      2@     @W@     @Q@              "@      $@      3@      @      .@      @      1@              �?              @      0@      I@      @      @      @      @@      3@              �?       @       @              "@              @                               @      @      4@                       @      2@      @                       @                      @      @      *@              �?               @      *@      >@      @      @      �?      ,@      0@              �?               @              E@       @      C@              @              @      5@      B@      @      $@      .@     �N@      I@               @       @      &@      @      8@               @               @                      ,@      2@      �?      �?      @      A@      &@              @              @              2@       @      >@              @              @      @      2@      @      "@      "@      ;@     �C@              @       @      @      @     �J@      "@      :@      �?      @              @      [@      `@      $@      *@      (@      T@      K@              �?              &@      @      J@      "@      9@      �?      @              @      [@      `@      "@      *@      (@      T@     �E@                              &@       @      H@      @      6@              �?              @     �Y@      ]@      @      @      @     �O@     �B@                              $@       @      @      @      @      �?      @                      @      (@       @       @      @      1@      @                              �?              �?              �?                                                      �?                              &@              �?                      @      a@      ?@      a@      2@      >@      @     �B@     �f@     �h@      9@      >@      U@     @h@     @c@       @      =@      <@     �S@      0@      F@      @      8@      �?      @       @      (@      R@      T@      @      "@      1@      H@     �M@              @      @      1@      @      8@      �?      ,@      �?      @              "@      4@      C@       @      @      "@      6@     �A@               @       @      (@       @      6@      �?      *@                              @      4@     �A@       @      �?       @      4@      8@               @       @      @       @      ,@              @                              @      @      .@       @              @       @      @               @       @      @      �?       @      �?      @                                      .@      4@              �?      @      (@      2@                                      �?       @              �?      �?      @              @              @               @      �?       @      &@                               @              �?                                                                                                      @                              @              �?              �?      �?      @              @              @               @      �?       @      @                               @              4@      @      $@               @       @      @      J@      E@       @      @       @      :@      8@               @      @      @      @      &@      @      @              �?       @      �?      E@     �@@      �?      @      @      0@      &@                       @       @              @              @              �?                      6@      5@      �?      @      @      $@       @                               @              @      @      �?                       @      �?      4@      (@                      @      @      @                       @                      "@              @              �?               @      $@      "@      �?              �?      $@      *@               @      �?      @      @      @               @              �?               @      @      "@                      �?      @      &@               @      �?      @              @               @                                      @              �?                      @       @                                      @     @W@      ;@      \@      1@      8@      @      9@     �[@     @]@      5@      5@     �P@     @b@     �W@       @      9@      7@      O@      &@      =@      @      =@              @              @     �P@     �P@      @      @      4@      K@      =@              @      @      0@              8@      @      *@               @              @     �F@      G@      @      @      1@      G@      8@              @      @      (@              3@      @       @               @               @      5@      .@      �?      @      @      :@      @              �?              @              @              @                               @      8@      ?@      @      �?      ,@      4@      2@               @      @      @              @              0@              �?                      5@      5@                      @       @      @                              @              �?              *@              �?                       @      @                       @       @      �?                                              @              @                                      3@      1@                      �?      @      @                              @              P@      7@     �T@      1@      5@      @      5@     �F@      I@      1@      1@     �G@      W@     �P@       @      6@      3@      G@      &@      P@      5@     �S@      ,@      4@       @      5@     �F@     �F@      ,@      0@      @@     �V@     �M@       @      5@      ,@     �D@      $@      H@      .@      I@      &@      &@      �?      2@     �D@     �A@      @      ,@      7@     @Q@     �C@              @      @      ;@       @      0@      @      <@      @      "@      �?      @      @      $@      @       @      "@      5@      4@       @      ,@      @      ,@       @               @      @      @      �?      �?                      @      @      �?      .@       @      @              �?      @      @      �?               @                                                               @              @              @              �?                                              @      @      �?      �?                      @      �?      �?      $@       @       @                      @      @      �?     �`@     �A@     �^@      0@      B@      2@      6@     @X@     �a@      1@      @@     �K@     `i@     �d@      0@      9@      1@     �M@      0@     �U@      :@     @Q@      &@      =@      *@      &@     �D@     @U@      (@      7@      A@     �X@      [@      &@      4@      0@     �@@      0@      ,@      �?       @                                      @                                       @      �?                                             @R@      9@     �P@      &@      =@      *@      &@      A@     @U@      (@      7@      A@     @X@     �Z@      &@      4@      0@     �@@      0@      B@      $@      4@       @      @      �?      @      5@      C@      �?      @      *@     �K@      @@      @      "@       @      *@       @      @      @       @                                      &@      (@      �?      �?      @      .@      @              @               @      �?      @      @       @                                      @       @      �?      �?       @       @       @               @                                                                                      @      $@                      �?      *@      @              �?               @      �?      ?@      @      2@       @      @      �?      @      $@      :@              @      $@      D@      9@      @      @       @      &@      @      1@       @      �?                                       @       @                              (@      @      �?                      @      �?      ,@      @      1@       @      @      �?      @       @      2@              @      $@      <@      4@       @      @       @      @      @     �B@      .@     �G@      "@      6@      (@      @      *@     �G@      &@      3@      5@      E@     �R@       @      &@       @      4@       @      2@      @      @              @                       @      &@       @      @      @      *@      1@              @      @      "@      @      2@      �?      @              @                      @      &@       @      @      @      *@      (@                      @       @      @               @      �?                                      �?                                              @              @      �?      �?              3@      (@     �D@      "@      3@      (@      @      @      B@      "@      .@      2@      =@      M@       @       @      @      &@      @      $@      @      *@      @      .@       @               @      *@              �?      @       @      @              @      �?      �?              "@      "@      <@      @      @      $@      @      @      7@      "@      ,@      .@      5@     �I@       @      @      @      $@      @     �F@      "@     �J@      @      @      @      &@      L@      L@      @      "@      5@      Z@      L@      @      @      �?      :@              B@      @      D@       @      @      @      @      H@      F@       @      @      *@      U@      C@      @      @              &@              5@      @      &@       @       @      @      �?      7@      8@      �?       @       @     �J@      3@      �?                      @              *@      �?      $@                      @      �?      1@      1@              �?      @      I@      "@                               @              @              @                                      @      $@              �?      @      &@       @                                              "@      �?      @                      @      �?      $@      @                             �C@      @                               @               @      @      �?       @       @                      @      @      �?      �?      @      @      $@      �?                       @               @      @      �?       @       @                      @      @      �?      �?      @              @      �?                       @                                                                       @      @                              @      @                                              .@       @      =@              �?       @      @      9@      4@      �?      @      @      ?@      3@      @      @              @              �?              4@                                      $@      @               @       @      @      @                              �?                              0@                                       @      @                              @      @                                              �?              @                                       @      �?               @       @      @      �?                              �?              ,@       @      "@              �?       @      @      .@      0@      �?      �?      @      8@      .@      @      @              @              @              @                              �?      *@       @              �?              @      $@              @               @              @       @      @              �?       @      @       @       @      �?              @      2@      @      @      �?              @              "@      @      *@      @      @              @       @      (@      @      @       @      4@      2@      �?              �?      .@               @              @      @       @              @      @      "@      @      @      @      *@      @                      �?      &@              @              @      @       @               @      @      "@       @      @      @       @      @                              &@               @                               @                      @       @                              �?      �?                                              @              @      @                       @              @       @      @      @      @       @                              &@               @                                              @      �?              �?                      @                              �?                      �?      @       @               @              �?      @      @                      �?      @      .@      �?                      @                              �?              �?                      �?      @                                      @                              @              �?      @      @              �?              �?      @                              �?      @      $@      �?                      �?                              @              �?                       @                              �?              @                              �?              �?      @      @                              �?      �?                                      @      @      �?                                �t�bub��      hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���LhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKmhnh4h7K ��h9��R�(KKm��hu�B�         4                    �?���K��?�	           ��@                          �4@2y�)%%�?           �@                           @S6cTe4�?�           p�@                            @�Z��f&�?n           ��@                            �?ˊ�ǣ�?�            �s@                           �?���,d�?k             g@������������������������       ��f��?0             S@������������������������       �����?;             [@	       
                   �0@nN,�4�?[             `@������������������������       ��$I�$I�?
             ,@������������������������       �74(���?Q            �\@                          �3@l;���k�?�            Pp@                           @+��k�P�?{            �f@������������������������       ��_�!p�?Y            �`@������������������������       ����ҧ�?"            �H@                           �?�HSw��?-            �S@������������������������       ��E��ӭ�?
             2@������������������������       ��{+H��?#            �N@                           �?�qǱ�?             H@                          �2@��@����?             9@������������������������       �r�q��?	             (@������������������������       ��5��?             *@                           �?J��LQ�?             7@������������������������       ��G�z��?             $@������������������������       ��θ�?	             *@       )                   �=@�8C'�r�?�           X�@       "                    �?K��x�3�?2           `�@                          �;@��
͵��?�            `q@                           �?FC�����?�             n@������������������������       ���f�?D            �]@������������������������       ����?J<�?F            �^@        !                    �?V������?            �B@������������������������       ��Q����?             4@������������������������       �Iє�?             1@#       &                   �8@P1o��#�?�           ��@$       %                   �6@L�<��	�?�            �v@������������������������       ��!pc��?o             f@������������������������       �6?��?x             g@'       (                    �?vna� �?�            �p@������������������������       ��;��1X�?:            �U@������������������������       ���8!&D�?p            �f@*       /                    @��
���?]            @a@+       .                     @r�q�?@             X@,       -                    �?zk&{��?$            �H@������������������������       �������?             *@������������������������       ����^B{�?             B@������������������������       ��d�����?            �G@0       3                   @A@Dc}h��?             E@1       2                    @ܶm۶m�?             <@������������������������       �     ��?             0@������������������������       ��8��8��?	             (@������������������������       �^N��)x�?             ,@5       T                   �5@ղ�S��?�           ��@6       E                   �1@T���?}           �@7       >                    @������?           �y@8       ;                   �0@d�6h��?�            `q@9       :                     �?��Ph���?A            @X@������������������������       ��-��?)             O@������������������������       ��	B�~�?            �A@<       =                     @w��lY��?s            �f@������������������������       ����ߠ��?Z            �`@������������������������       ��q���?             H@?       B                     �?c���E�?Y             a@@       A                    @���?            �D@������������������������       ��?�(��?             :@������������������������       ��.�?�P�?
             .@C       D                    @I/=ө]�?>            �W@������������������������       �R�}e�.�?             :@������������������������       �T#G�h�?.            @Q@F       M                    �?�E�f�?p           8�@G       J                   �3@�F�yu�?4            ~@H       I                    @�]���?�?�            q@������������������������       �Wr!�m�?s            @g@������������������������       ��p�j�A�?3            �U@K       L                     @*�&�o_�?�            �i@������������������������       ����`d�?q            �d@������������������������       ��p=
ף�?             D@N       Q                    @�њ��?<           8�@O       P                    @BC����?�            `x@������������������������       ���|Zc�?Q             `@������������������������       ��4@��}�?�            Pp@R       S                   �2@��`b��?M             `@������������������������       ��*f����?             E@������������������������       �(~�[�?6            �U@U       `                    �?�B�����?            �@V       [                    @ɼ9�=�?�            �v@W       Z                   �=@    ���?�             p@X       Y                   �8@��#ӱ��?�            �m@������������������������       �M���3��?\            @a@������������������������       ������?>            �X@������������������������       �H�z�G�?
             4@\       _                   �=@WZX�?G            �[@]       ^                     �?�8EGr��??             Y@������������������������       �;�;��?$             J@������������������������       ��8��8��?             H@������������������������       ��������?             $@a       h                    @u0F,#�?            }@b       e                     �?^6wJ��?�            �y@c       d                    �?ߗ���?9            @W@������������������������       �c��gS~�?             =@������������������������       �     @�?)             P@f       g                    @�|)����?�            �s@������������������������       ��k����?7             V@������������������������       �	�GHZ��?�            �l@i       l                   �=@˕6�#��?!            �K@j       k                   �6@�Q����?             D@������������������������       �VUUUUU�?             "@������������������������       ��� =�	�?             ?@������������������������       �$߼�x�?             .@�t�bh�h4h7K ��h9��R�(KKmKK��h��B�@       �{@     �V@     �r@      =@     �W@     �@@     @S@     H�@     ��@     �R@     @T@     �c@      �@      {@      *@     �P@     �I@      `@      J@     �g@     �B@     `c@      .@     @P@      8@      D@     �]@      h@      @@     �K@     �U@      p@     �i@      $@     �B@      A@      S@     �C@     �X@      @     �H@      @      @              @     @R@     �V@      @      ,@      <@     �\@     �P@              @      @     �A@      "@     �T@      @     �G@      @      @              @     �Q@     @T@      @      &@      :@     @\@      P@              @      @      A@      @      H@       @      :@      @       @              @     �H@     �J@      �?      �?      .@      P@      7@              @              0@      @      >@       @      ,@      @                       @      4@      :@      �?      �?      "@      H@      &@              @              *@      �?      ,@              @                              �?      $@      *@                      @      9@                                       @      �?      0@       @      "@      @                      �?      $@      *@      �?      �?      @      7@      &@              @              &@              2@              (@               @              �?      =@      ;@                      @      0@      (@              �?              @       @                                                              @       @                               @                                                      2@              (@               @              �?      9@      3@                      @      ,@      (@              �?              @       @     �A@      @      5@       @      @               @      5@      <@      @      $@      &@     �H@     �D@              @      @      2@      @      8@      @      &@       @       @               @      0@      9@      �?      @       @      <@     �@@              @       @      0@      @      6@      @      "@       @       @               @      *@      ,@      �?      @      �?      5@      5@              @               @      @       @               @                                      @      &@                      �?      @      (@                       @       @      �?      &@              $@              �?                      @      @       @      @      "@      5@       @                      @       @              @                                                      @               @                      @      �?                      @                      @              $@              �?                       @      @              @      "@      1@      @                               @              .@               @               @                      @      $@      @      @       @       @      @                              �?       @      @                               @                              $@       @      �?      �?       @      �?                              �?              @                                                              �?       @      �?      �?       @                                      �?              �?                               @                              "@                                      �?                                              $@               @                                      @              �?       @      �?               @                                       @      @               @                                      �?                       @      �?                                                              @                                                       @              �?                               @                                       @     @W@      >@     �Z@      $@      M@      8@     �A@      G@     @Y@      9@     �D@     �M@     �a@      a@      $@      >@      =@     �D@      >@     �U@      =@     �X@      @     �B@      2@      ?@      F@     �W@      4@      <@      I@     �`@     �_@      @      6@      3@      ?@      7@      D@      &@      2@       @      "@      @      @      &@      F@      @      &@      @      E@     �@@      @      @      @      "@      "@      B@      $@      0@       @      @      @      @      &@     �@@      @       @      @      D@      :@      @      @      @      "@       @      7@      �?      &@              �?              @       @      3@       @                      3@      *@      @      @      �?      @      @      *@      "@      @       @      @      @              @      ,@      @       @      @      5@      *@       @      @      @      @      @      @      �?       @              @               @              &@              @               @      @                                      �?      @      �?      �?              @                              @              �?                      @                                                              �?                               @              @               @               @       @                                      �?     �G@      2@      T@      @      <@      (@      9@     �@@     �I@      .@      1@     �G@     @W@     �W@      �?      .@      *@      6@      ,@      >@      &@     �F@      @      *@      "@      &@      ;@     �@@      @      0@      4@     �G@      N@              @      $@      ,@       @      *@      @      2@       @      @      @       @      *@      $@      @      @      "@      A@      ;@              �?      @      &@      �?      1@      @      ;@      �?      "@      @      @      ,@      7@       @      *@      &@      *@     �@@              @      @      @      �?      1@      @     �A@       @      .@      @      ,@      @      2@      "@      �?      ;@      G@      A@      �?      &@      @       @      (@       @      �?      1@                              @      �?      &@      �?      �?      @      4@      ,@               @      @      �?      @      .@      @      2@       @      .@      @      $@      @      @       @              7@      :@      4@      �?      "@              @       @      @      �?       @      @      5@      @      @       @      @      @      *@      "@      @      $@      @       @      $@      $@      @      @      �?      @      @      3@      @      @              @      @      (@      @      @      "@              @      @       @      @       @      �?      @              .@               @              @       @      @      @      �?      �?              @      @       @      �?      �?                              �?               @              @      �?       @              �?                                      �?      �?      �?      �?      @              ,@                                      �?       @      @              �?              @      @      �?              �?              �?      @      @      @      �?               @      @       @      �?      @       @               @       @              @      @               @               @       @      �?       @      �?              �?      @      �?      �?      @      @      @       @      @      @                              �?       @      �?       @                      �?      �?      �?      �?              @      @       @              @                                                                                      �?      �?                      @       @      @                                              �?       @      �?       @                      �?                      �?                       @       @                               @              �?                              �?                      @                      @                              @     @o@      K@     `b@      ,@      =@      "@     �B@      {@      {@     �E@      :@      R@      v@     �l@      @      >@      1@     �J@      *@      d@      *@      S@      @      @      �?      :@     �u@     @t@      3@      (@      B@      j@      a@              &@      "@      6@      @     �D@      @      (@                              @     �a@     @Z@      @      @      $@     �M@      :@              �?               @              2@      @      $@                              �?     @\@     �Q@              @      @      C@      *@                               @              @               @                                     �G@      6@               @              1@      �?                                              @              �?                                      :@      5@               @              "@                                                      @              �?                                      5@      �?                               @      �?                                              (@      @       @                              �?     �P@      H@              @      @      5@      (@                               @              "@      @       @                              �?     �K@     �@@              �?      �?      1@      "@                               @              @              @                                      &@      .@               @      @      @      @                                              7@               @                              @      >@     �A@      @              @      5@      *@              �?                              �?                                              @      @      6@                      �?      @       @                                                                                              @      @      2@                              �?                                                      �?                                                      @      @                      �?      @       @                                              6@               @                                      7@      *@      @              @      0@      &@              �?                              @              �?                                       @      "@      @                      @       @                                              0@              �?                                      5@      @                      @      *@      "@              �?                             �]@      $@      P@      @      @      �?      6@      i@     `k@      0@      @      :@     �b@     �[@              $@      "@      4@      @      N@      �?      9@       @                      @     �[@     �_@      "@       @       @      N@      N@               @       @       @              @@              1@       @                      �?     �R@     @P@      @      �?      @      <@     �B@              �?              @              2@              ,@       @                              F@      H@      �?      �?      @      5@      <@              �?              @              ,@              @                              �?      ?@      1@       @              �?      @      "@                               @              <@      �?       @                              @     �A@      O@      @      �?       @      @@      7@              �?       @      @              5@      �?       @                              @      ;@     �N@      @               @      6@      1@              �?                              @                                                       @      �?       @      �?              $@      @                       @      @             �M@      "@     �C@       @      @      �?      2@     �V@      W@      @      @      2@     �V@      I@               @      @      (@      @     �F@      @      B@      �?      @      �?      @     �R@      Q@      @      @      $@      S@      B@              �?      @      @      @      ,@      @       @              @      �?      @      3@      =@       @       @              9@      0@                       @                      ?@      @      <@      �?                       @      L@     �C@      @      @      $@     �I@      4@              �?       @      @      @      ,@      @      @      �?      �?              &@      0@      8@                       @      ,@      ,@              @      @       @       @       @                                              @      @      @                      �?      @       @              @       @      @              (@      @      @      �?      �?               @      "@      3@                      @      @      (@              �?      �?      �?       @     �V@     �D@     �Q@      $@      9@       @      &@     �V@      [@      8@      ,@      B@     �a@     �W@      @      3@       @      ?@      @     �D@      4@      @@              &@              �?      L@     �L@      @      @      "@     @P@      D@              @       @       @      @      8@      $@      6@               @                      C@     �I@      @      @       @     �F@      @@              @      �?       @      @      4@      $@      6@              @                      C@     �I@      @      @       @     �A@      @@              @      �?       @      @      $@       @      ,@              @                      <@     �B@      �?               @      4@      2@                      �?               @      $@       @       @              �?                      $@      ,@      @      @      @      .@      ,@              @               @      �?      @                              @                                              �?              $@                      �?                              1@      $@      $@              @              �?      2@      @       @      @      �?      4@       @               @      �?      @       @      0@      $@      $@               @              �?      2@      @              @      �?      3@      @               @      �?      @              0@      @      �?                              �?      @      @              @              @      @              �?      �?      @                      @      "@               @                      &@      �?                      �?      ,@      �?              �?               @              �?                              �?                                       @                      �?      @                                       @     �H@      5@     �C@      $@      ,@       @      $@      A@     �I@      2@      @      ;@     �S@      K@      @      *@      @      7@      �?     �E@      5@      <@      "@      @       @       @      <@     �I@      2@      @      :@     @R@     �F@      @      *@      @      4@              @      �?      @      @      �?       @      @      *@      "@       @               @      1@      @              @      @      @               @               @                               @      @       @                              "@      @                                              @      �?      @      @      �?       @      �?      @      @       @               @       @      �?              @      @      @             �B@      4@      5@      @      @      @      @      .@      E@      0@      @      2@      L@     �C@      @      "@      @      ,@              $@               @      @              @      @      @      .@      $@              @      "@      $@       @      �?              $@              ;@      4@      3@      �?      @      @       @      &@      ;@      @      @      (@     �G@      =@      �?       @      @      @              @              &@      �?      $@               @      @                              �?      @      "@                              @      �?      @              @      �?      @              �?      @                              �?      @      @                               @      �?                      @              �?                                                      �?      @                                                      @              �?      �?      @              �?      @                                       @      @                               @      �?                      @              @              �?                                                       @                              �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��bvhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKqhnh4h7K ��h9��R�(KKq��hu�B�         8                   �2@U��"̅�?�	           ��@                           �?��>�m��?�           ؐ@                            @��Cȃ��?            �y@                           �?����U�?�            Ps@                           �?6�80\��?/             S@                            �?����D��?            �@@������������������������       �     @�?             0@������������������������       ���'s�	�?             1@	       
                     �?k�F	��?            �E@������������������������       �*L�9��?             6@������������������������       �"�����?             5@                          �0@���x�?�             m@                            �?�w^�V�?$            �H@������������������������       �ԍx��?             C@������������������������       ��C��2(�?	             &@                           �?I� ��?r             g@������������������������       ���{�b��?D            @\@������������������������       �f "` �?.            �Q@                          �1@�$��C�?;             Y@                           @�E��Y��?%             O@                           �?�(\����?             D@������������������������       �������?             *@������������������������       �������?             ;@������������������������       ��4_�g�?             6@                           �?UH�� �?             C@������������������������       �،A��_�?	             1@������������������������       ��U̠ç�?             5@       )                    �?^;:Q�?�           �@       "                   �0@��/ �?�            �r@                           �?�>�\��?+             O@������������������������       �b�r���?	             .@        !                     @��Lp�?"            �G@������������������������       ��x?r���?            �@@������������������������       �$I�$I��?             ,@#       &                    @�>a0�D�?�            @m@$       %                    �?v�����?F             [@������������������������       �>�ؑ�J�?.            @R@������������������������       ��mTM�?            �A@'       (                    @��N8�?K            �_@������������������������       �     ��?             0@������������������������       ��bX�h�?D            �[@*       1                   �0@}�����?�            Pw@+       .                    @�d� ��?*            �P@,       -                    @B�0�~��?             F@������������������������       ��g���u�?             ;@������������������������       ��d��E�?
             1@/       0                     �?�r��_�?             7@������������������������       ��T�x?r�?	             &@������������������������       ���8��8�?             (@2       5                    @����?�             s@3       4                   �1@J�I�3�?|            @j@������������������������       ������?>            �X@������������������������       ���>�y�?>            �[@6       7                    �?�q�1�?;             X@������������������������       �t�E]t�?             &@������������������������       �{�/��>�?4            @U@9       R                    �?y,w\���?           &�@:       I                     �?*��c:4�?%           ��@;       B                   �8@YyN��?%           �|@<       ?                    �?�X���?�            Pv@=       >                    @��3� ��?t            `h@������������������������       �	j*D�?A             Z@������������������������       �\�ڔ��?3            �V@@       A                   �5@��I�?j            @d@������������������������       ��8��8��??             X@������������������������       ���rW��?+            �P@C       F                   �<@�T�6|��?G             Z@D       E                     �?�.�{B��?4            �S@������������������������       �
ףp=
�?             D@������������������������       �mvq`���?             C@G       H                    �?�h��9�?             :@������������������������       ��2�tk~�?             "@������������������������       �Iє�?             1@J       Q                   �>@i)F��?            px@K       N                   �7@D�����?�            `w@L       M                    �?:g����?�            �o@������������������������       �*.c!�?X            �a@������������������������       ���sG��?N            @\@O       P                    @�~ɖ���?O            �]@������������������������       ��g���e�?;             V@������������������������       ��QNZ���?             ?@������������������������       �J,�ѳ�?             1@S       b                   �7@��5���?�           ��@T       [                    �?������?�           ��@U       X                    �?�P�`�S�?2             W@V       W                   �5@�fG-B��?             5@������������������������       ��������?             (@������������������������       ��<ݚ�?             "@Y       Z                    �?����7�?$            �Q@������������������������       ���)x9�?             <@������������������������       ��hZ_�?            �E@\       _                    @�gV��~�?�           P�@]       ^                    �?�w`*�}�?B           h�@������������������������       ��ƭ���?�            x@������������������������       �W������?L           `�@`       a                     �?DEM���?Y            �`@������������������������       �L�w�Z��?            �A@������������������������       �H�}8g�?A             Y@c       j                    �?�"�f�?           x�@d       g                    @r�x�'|�?           p|@e       f                   �<@n[_}P��?�            @m@������������������������       ��Wg:�?�?g            �c@������������������������       ��˦1i�?.            �S@h       i                    �?7�8����?�            �k@������������������������       �8��;��?2             U@������������������������       �u����?X             a@k       n                   �:@��鲲��?�            �x@l       m                    @g�Y�X\�?�            �l@������������������������       �z)[IPo�?:            �X@������������������������       �o�)�Ư�?Q            @`@o       p                    @r��tq'�?l            �d@������������������������       �چ=	�?/            �R@������������������������       �����kE�?=            @V@�t�bh�h4h7K ��h9��R�(KKqKK��h��BC       @z@     �S@     �u@      :@     �T@      5@     �Q@     p�@     ��@      Q@     �T@     �c@     �@     �y@      *@      N@      J@      `@     �Q@     �_@       @     �U@              @              $@     `r@     �k@      @       @      5@     �e@     @R@              &@      @      7@      "@     �H@       @      =@               @              @     @a@     �T@      �?       @       @     �N@      0@              @              @      @     �@@              "@                               @     �]@     �R@               @      @     �E@      (@              @               @      @      ,@              �?                                      3@      3@                      @      *@      @                              �?       @      @              �?                                      ,@      @                      �?      @      @                                              @              �?                                      @      @                              @      �?                                               @                                                      "@                              �?      @       @                                              "@                                                      @      0@                      @      @                                      �?       @      @                                                       @      "@                      @       @                                      �?              @                                                      @      @                              @                                               @      3@               @                               @      Y@     �K@               @              >@      "@              @              �?       @      @              @                                      <@      @              �?              @                                                      @              @                                      2@      @              �?              @                                                      �?                                                      $@                                                                                              .@              @                               @      R@     �H@              �?              7@      "@              @              �?       @      @              @                                     �F@      B@                              ,@       @                                               @               @                               @      ;@      *@              �?              "@      �?              @              �?       @      0@       @      4@               @              �?      3@      "@      �?              @      2@      @                              @              (@       @       @               @                      0@      @      �?              @      (@      @                                              "@       @                       @                      @      @      �?               @      "@      @                                              @                                                      @              �?              �?      @                                                      @       @                       @                       @      @                      �?      @      @                                              @               @                                      $@       @                       @      @                                                      @              2@                              �?      @       @                              @                                      @               @              "@                                                                               @                                      @               @              "@                              �?      @       @                              @                                                     @S@      @      M@               @              @     �c@     �a@      @      @      *@     �[@     �L@              @      @      1@      @      C@      @      1@                               @      X@     �R@                       @      H@      *@              �?               @              "@               @                                      1@      7@                              $@      �?                                                               @                                      @      @                                      �?                                              "@                                                      &@      1@                              $@                                                      @                                                      &@      ,@                              @                                                      @                                                              @                              @                                                      =@      @      .@                               @     �S@     �I@                       @      C@      (@              �?               @              ,@      �?      @                                      9@      ?@                      �?      7@      @              �?               @               @      �?      @                                      4@      .@                              4@      @              �?              �?              @              �?                                      @      0@                      �?      @       @                              �?              .@       @      $@                               @      K@      4@                      �?      .@      @                                               @              @                                      "@                                       @                                                      *@       @      @                               @     �F@      4@                      �?      *@      @                                             �C@      @     �D@               @              @      N@     �P@      @      @      &@     �O@      F@              @      @      .@      @      *@               @                                      (@      0@                       @       @      @                              �?              "@              @                                      @      .@                              @      �?                                              @              @                                      @      @                              @      �?                                               @               @                                       @      &@                                                                                      @              @                                      @      �?                       @      �?      @                              �?              @                                                       @      �?                       @      �?      �?                              �?              �?              @                                      @                                              @                                              :@      @     �@@               @              @      H@      I@      @      @      "@     �K@     �B@              @      @      ,@      @      1@       @      >@               @              @      3@      >@      @      @      @      C@     �@@               @       @      $@      @      @      �?      .@               @               @      &@      0@      �?      @      @      ,@      $@               @       @      @      @      $@      �?      .@                              �?       @      ,@      @      @      @      8@      7@                              @      �?      "@      �?      @                               @      =@      4@                       @      1@      @              @      �?      @      �?      @      �?      �?                                                                               @                                                       @               @                               @      =@      4@                       @      .@      @              @      �?      @      �?     `r@     �Q@     0p@      :@     �S@      5@      N@     �p@     y@      O@     �R@      a@     p}@     @u@      *@     �H@     �H@     �Z@     �N@     �[@      9@      L@      @      ,@      @      ,@     @U@      d@      .@      3@      ?@      c@     �Y@              *@      &@      3@      0@     �G@      @      8@      �?      @              $@      E@     �Y@      $@      &@      5@     �W@     @P@              @      @      $@      $@      @@              0@               @              @      @@     @W@      @      @      2@     �T@     �I@              @      @       @      $@      .@              "@              �?              �?      1@     �I@      �?      @      *@     �M@      3@                                      @       @              @              �?              �?      @      @@              @      (@      9@      @                                      @      @              @                                      *@      3@      �?              �?      A@      *@                                              1@              @              �?              @      .@      E@      @      �?      @      8@      @@              @      @       @      @      $@              @              �?               @       @      ?@              �?      @       @      6@              �?      �?               @      @              �?                              �?      @      &@      @               @      0@      $@               @       @       @       @      .@      @       @      �?      �?              @      $@      "@      @      @      @      (@      ,@              �?               @              $@      �?       @      �?      �?              �?      $@      @      @      @      @      (@      @              �?              @              @              �?      �?      �?              �?      @      @      �?              @       @      @              �?              @              @      �?      @                                      @       @       @      @              @      @                              �?              @       @                                      @              @      @                              @                              �?              @       @                                      �?               @                                      �?                                               @                                              @              �?      @                              @                              �?              P@      6@      @@       @      &@      @      @     �E@     �M@      @       @      $@      M@      C@              "@       @      "@      @      P@      6@      @@      �?      &@       @      @     �E@     �M@      @      @      "@     �H@      C@               @      @      "@      @     �G@      @      1@      �?       @      �?       @      D@     �G@      @      @      @      A@      8@              @      @      @      @      <@       @      @               @                      =@      :@              @      �?      8@      *@              �?              @      �?      3@      @      &@      �?      @      �?       @      &@      5@      @      �?      @      $@      &@              @      @      �?       @      1@      1@      .@              @      �?       @      @      (@      �?       @      @      .@      ,@              @      @       @      @      *@      @      .@              @      �?               @      "@               @      @      *@      (@              @       @      �?       @      @      (@                                       @      �?      @      �?              �?       @       @                      �?      �?      �?                              �?              �?                                       @      �?      "@                      �?       @                     �f@      G@     `i@      7@      P@      2@      G@     `f@      n@     �G@     �K@     @Z@     �s@     �m@      *@      B@      C@     �U@     �F@      `@      4@      W@      "@      3@      @      4@     �a@     �d@      6@     �@@      J@      j@     �^@              0@      .@      M@      "@      9@              @              �?              @       @      @       @      @       @      2@      $@              @       @       @               @              @              �?              �?              �?       @      @       @      @                                                       @              @                              �?              �?              �?       @       @                                                                                      �?                                       @       @              @                                                      7@                                              @       @      @                              (@      $@              @       @       @              &@                                                      �?      @                                      "@                       @       @              (@                                              @      @       @                              (@      �?              @                              Z@      4@     @V@      "@      2@      @      ,@     �`@     �c@      4@      >@      I@     �g@      \@              (@      *@      L@      "@     �W@      4@     �P@      "@      .@       @      $@     �^@     �a@      ,@      ;@     �D@     �c@     �Y@              (@      &@      J@      "@     �F@      &@      A@       @      "@       @      @      >@      @@      @      .@      7@      Q@      L@              @      $@      :@      @      I@      "@     �@@      @      @              @     @W@      [@      @      (@      2@     �V@     �G@              @      �?      :@      @      "@              6@              @       @      @      &@      3@      @      @      "@      @@      "@                       @      @              @              &@                                      @      @              �?      �?      $@                                                      @              &@              @       @      @       @      ,@      @       @       @      6@      "@                       @      @              K@      :@     �[@      ,@     �F@      ,@      :@     �B@     �R@      9@      6@     �J@     @[@     �\@      *@      4@      7@      =@      B@      7@      2@      Q@      @      >@      (@      ,@      &@     �@@      &@      ,@      B@     �E@      L@       @      (@      .@      &@      A@       @      @      G@       @      4@      @       @       @      *@      @      @      .@      5@      E@      @      @       @      @      (@      @      @      5@              0@      @              @      (@       @      @      $@      2@     �B@              �?       @      @      @      @      @      9@       @      @               @      �?      �?      @      @      @      @      @      @      @               @      "@      .@      &@      6@      @      $@      @      (@      @      4@      @       @      5@      6@      ,@      @       @      @      @      6@       @      �?       @              @      �?      @       @      &@                      @      *@      @      @              @      �?      &@      @      $@      ,@      @      @      @      @      �?      "@      @       @      2@      "@      "@       @       @       @      @      &@      ?@       @     �E@       @      .@       @      (@      :@      E@      ,@       @      1@     �P@     �M@      @       @       @      2@       @      3@       @      7@      @      @               @      8@     �A@      �?      @      $@     �C@     �B@      @       @              @      �?      ,@              (@      @      @              @      @      "@              @      @      3@      (@                              @      �?      @       @      &@      �?      @              @      3@      :@      �?      �?      @      4@      9@      @       @              @              (@      @      4@      @       @       @      @       @      @      *@      @      @      ;@      6@       @      @       @      &@      �?      @       @      ,@       @      �?      �?              �?      @       @       @      @      @      @       @      @      @      @              @      @      @      �?      @      �?      @      �?      @      @      �?      @      4@      1@               @      �?      @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJL��nhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�         @                    �?<ҹ)v��?�	           ��@       !                    �?��T��	�?)           ��@                           �?�:�N��?;           0~@                            @��h'<�?|            �g@                          �2@촠S��?S            ``@                           �?A�m�1�?             A@������������������������       ��U̠ç�?             5@������������������������       �����W�?
             *@	       
                   �<@����H��?<            @X@������������������������       �6\�҇��?4            �U@������������������������       ��ˠT�?             &@                           �?bΊx��?)             M@                          �7@)\���(�?            �A@������������������������       ��T'"7�?             ;@������������������������       �      �?              @                          �3@��Moz��?             7@������������������������       ����>4��?             ,@������������������������       �0�����?             "@                          �4@!N�x;��?�            `r@                          �1@ C��ڔ�?O            �^@                           �?"���V�?            �A@������������������������       �������?             ,@������������������������       �Z�eY�e�?             5@                            @L�9���?9             V@������������������������       ��;��1X�?            �E@������������������������       �˪Qj��?            �F@                          �;@��Eb_��?p            `e@                            �?|�o��?X            �`@������������������������       �u�t��?            �B@������������������������       �L���O5�?@            �X@                            �?3�tk~X�?             B@������������������������       ��h$���?             .@������������������������       �W�7�L�?             5@"       1                   �4@z�'-�"�?�           H�@#       *                   �0@����ї�?           `|@$       '                     �?н��9q�?$            �L@%       &                    @��D���?             5@������������������������       ��G�z��?             $@������������������������       ���!pc�?             &@(       )                     �?�"e����?             B@������������������������       ��"e����?             2@������������������������       ��"e����?             2@+       .                     @H��"W"�?�            �x@,       -                   �3@}�!�Z�?�            �s@������������������������       �G�DX��?�            @m@������������������������       �^�"R��?,            �S@/       0                    �?��U���?5            @U@������������������������       ��E����?             B@������������������������       �1�&�}��?            �H@2       9                    �?�X0��"�?�            0t@3       6                     @v����?q            �d@4       5                   �6@�g�z��?]             a@������������������������       �     ��?*             P@������������������������       ���69	@�?3            @R@7       8                   �7@�P�a�r�?             >@������������������������       �UUUUUU�?	             (@������������������������       ��E��ӭ�?             2@:       =                    @T�C,���?f            �c@;       <                    @RC4%�?+             Q@������������������������       �R���Q�?             D@������������������������       �����X�?             <@>       ?                   �8@�|���?;             V@������������������������       �*x9/��?$             L@������������������������       �     0�?             @@A       `                    �?�q�Y��?�           ��@B       Q                   �6@-�qj�<�?�           `�@C       J                    �?�#IP�o�?z           ��@D       G                   �2@��WV/�?�             j@E       F                    �?C|��'a�?:            @U@������������������������       ���yqY��?            �A@������������������������       �-C��6�?#             I@H       I                   �4@�b��"�?T            �^@������������������������       �lz�c�u�?-            �O@������������������������       �!Ce����?'             N@K       N                    �?�Kz��?�            @v@L       M                      @�	"P7��?             3@������������������������       ��2�tk~�?             "@������������������������       ��(\����?             $@O       P                   �2@��=ȟ�?�            u@������������������������       �K�DSue�?V            �_@������������������������       �y2FЋ��?�            `j@R       Y                   �=@B��m|n�?|            �@S       V                     �?�`�}7��?,           �}@T       U                   �;@)O���?a             b@������������������������       �D��{�?L            �\@������������������������       ��� Ce��?             >@W       X                     @ˀ0��?�            �t@������������������������       �z|���?P            @^@������������������������       �\D��K��?{            @j@Z       ]                     �?�c4O��?P             a@[       \                    @xvJ;��?            �F@������������������������       ����Kϟ�?             =@������������������������       �     @�?	             0@^       _                    �?��H�~Z�?6             W@������������������������       �
ףp=
�?             4@������������������������       �����K�?*             R@a       p                   �3@}il�>F�?�           �@b       i                    @�#w����?o           �@c       f                     �?�1�	���?�            �m@d       e                   �0@�6E��?1            @R@������������������������       ��)O�?             2@������������������������       �M�.���?%            �K@g       h                    �?��m�=�?j            �d@������������������������       ���(\���?             $@������������������������       ��1�g\ �?d            `c@j       m                    �?X3�Ƣ�?�            @u@k       l                    �?���ލL�?             ;@������������������������       ��ˠT�?	             &@������������������������       �      �?	             0@n       o                    @���O��?�            �s@������������������������       �ʑªS��?�            @k@������������������������       �i��S��??            �W@q       x                    �?�v�T��?B           �@r       u                    @?���2��?�            @w@s       t                    @hОτ�?i            �b@������������������������       �Z4���?_            �`@������������������������       ��@�m�?
             1@v       w                   �<@^ 꼆��?�            �k@������������������������       ��/��>��?�            �i@������������������������       �P�|�@�?             1@y       |                    @1U:L��?E           x�@z       {                   �;@!�����?F            �\@������������������������       �������?:             X@������������������������       �&���^B�?             2@}       ~                    @��҈��?�            �y@������������������������       �[1N��?�            �r@������������������������       ��\����?G            �\@�t�bh�h4h7K ��h9��R�(KKKK��h��BhK       |@     �U@      u@      F@      R@      C@     �P@     ؀@     H�@     �P@      U@     @c@     Ȃ@     �z@      1@     �T@     �P@      b@      H@     �c@      7@     �U@      @      5@      @      0@     `m@     �m@      5@      0@      =@     �e@     �_@       @      ;@      2@     �C@      2@     �R@      "@     �E@       @      .@       @      @      F@     �R@      $@      $@      $@     �L@      M@       @      (@      .@      =@      $@      :@      @      $@               @               @      1@     �F@      @       @      @      6@      2@              @      @      @      @      3@      @       @              �?               @      "@      D@              @       @      .@      ,@              �?      @      @      @      (@               @                                       @       @                               @      �?                              �?              @               @                                      @      @                                      �?                                              @                                                      @      �?                               @                                      �?              @      @      @              �?               @      �?      @@              @       @      *@      *@              �?      @      @      @      @              @                              �?      �?      =@              @       @      *@      $@              �?      @      @      @              @                      �?              �?              @                                      @                                              @               @              �?                       @      @      @      @       @      @      @              @       @      @       @      @               @                                      @      @      @               @       @       @              @              @              @              �?                                      @      �?      @              �?               @              @              @              �?              �?                                              @                      �?       @                                                                                      �?                      @      �?      �?      @              @       @               @       @               @                                      �?                       @                      @              @                       @                                                                                      �?      �?      �?                               @                       @               @      H@      @     �@@       @      *@       @      @      ;@      >@      @       @      @     �A@      D@       @      @       @      6@      @      4@      �?      @              @                      6@      0@                      @      5@      2@                              $@              @                               @                       @      @                              &@      @                                              �?                                                      @                                      @      �?                                              @                               @                      �?      @                              @      @                                              .@      �?      @              @                      ,@      &@                      @      $@      ,@                              $@              @              @                                      $@      @                       @      @      @                              @              $@      �?      @              @                      @      @                      �?      @       @                              @              <@      @      :@       @       @       @      @      @      ,@      @       @      @      ,@      6@       @      @       @      (@      @      4@      @      8@              @       @      @      @      $@      @       @      @      ,@      6@       @       @      @       @       @      $@               @               @                              @       @              �?       @      @      �?                      @              $@      @      6@               @       @      @      @      @      �?       @       @      (@      1@      �?       @      @       @       @       @      �?       @       @      @              �?              @       @                                              @      @      @       @      @      �?                       @                              @                                                      @                               @               @       @       @              �?              �?       @                                                      @      @       @      U@      ,@      F@      @      @      @      $@     �g@     `d@      &@      @      3@     @]@     @Q@              .@      @      $@       @     �J@      �?      0@      @      �?              @     `c@     @W@      �?      �?      &@     �P@      >@              "@       @       @      @      @                                                     �@@      $@              �?              @                                                       @                                                      @       @              �?              @                                                       @                                                       @      @              �?              �?                                                                                                              @      @                               @                                                      @                                                      :@       @                              @                                                       @                                                      *@      �?                               @                                                       @                                                      *@      �?                               @                                                     �G@      �?      0@      @      �?              @     �^@     �T@      �?              &@     �M@      >@              "@       @       @      @      A@      �?      @              �?              @     �Z@     @Q@      �?              @     �G@      6@              @       @       @      @      ;@      �?      @                              @     @R@     �K@      �?              @     �A@      .@              @       @       @      @      @              �?              �?                      A@      ,@                      �?      (@      @              �?                              *@              $@      @                      �?      .@      ,@                      @      (@       @              @                       @      @              @                                      "@      @                               @       @                                              @              @      @                      �?      @      @                      @      @      @              @                       @      ?@      *@      <@              @      @      @      B@     �Q@      $@      @       @     �I@     �C@              @      �?       @      @      0@      @      2@               @               @      1@      F@       @      @       @      @@      3@               @               @              (@      @      1@                               @      .@     �D@       @      @       @      9@      *@                                               @      @      @                              �?      @      :@               @      �?      *@      @                                              $@      �?      *@                              �?      "@      .@       @      �?      �?      (@       @                                              @      �?      �?               @                       @      @                              @      @               @               @              @                               @                              �?                               @      �?                               @                      �?      �?                                       @       @                              @      @               @                              .@      @      $@              @      @      @      3@      :@       @       @      @      3@      4@              @      �?      @      @      @      �?      "@              �?      @      �?      @      @      @               @      .@      $@              �?              �?              @      �?      @                      @      �?      @      @       @              �?       @      @              �?              �?               @              @              �?                      �?              @              �?      @      @                                               @      @      �?               @               @      (@      7@       @       @      @      @      $@              @      �?      @      @       @      @      �?                                      @      5@                       @      @      @               @               @      �?              @                       @               @      @       @       @       @       @      �?      @              �?      �?      @       @     0r@     �O@     `o@     �C@     �I@      @@     �I@      s@     �u@     �F@      Q@     @_@     �z@      s@      .@      L@      H@     �Z@      >@     �[@     �B@      b@      2@      <@      =@      8@     �R@      [@      8@      F@     @Q@     �d@      d@      @     �B@      =@     �F@      7@      Q@       @      O@      "@      @      @      @     �O@     �P@      $@      3@      7@     �[@     @P@              $@      @      =@      @      9@      �?      ,@              �?       @              B@     �@@              @      $@      K@      ,@              @      �?      @       @      @      �?      @                                      0@      6@                      @      4@      @              �?              @               @              �?                                      @       @                      @      &@      �?                              @              @      �?      @                                      &@      ,@                      �?      "@      @              �?              �?              4@               @              �?       @              4@      &@              @      @      A@      "@               @      �?       @       @      *@              �?              �?                      (@      @              @      @      (@      @               @              �?       @      @              @                       @               @      @              �?       @      6@      @                      �?      �?             �E@      @      H@      "@       @      @      @      ;@      A@      $@      *@      *@      L@     �I@              @       @      7@      �?      �?       @      @                                              �?      @      @               @                                                      �?               @                                              �?       @      @                                                                               @      @                                                      �?       @               @                                                      E@      @     �E@      "@       @      @      @      ;@     �@@      @       @      *@      K@     �I@              @       @      7@      �?      8@              1@      �?      �?              �?      3@      5@               @      @      4@      ,@              �?               @              2@      @      :@       @      �?      @      @       @      (@      @      @      $@      A@     �B@              @       @      5@      �?      E@      =@     �T@      "@      9@      8@      1@      &@     �D@      ,@      9@      G@      L@     �W@      @      ;@      :@      0@      4@     �D@      7@     @Q@      @      1@      4@      &@      $@      @@      $@      (@      =@      K@     �U@      �?      (@      0@      &@      ,@      .@      1@      5@      �?       @      @      �?      �?      @      �?      @      @      4@      2@              "@      �?       @      @       @      1@      5@              @      @      �?      �?      @      �?      @      @      &@      2@              @               @       @      @                      �?      @                                                              "@                      @      �?              @      :@      @      H@      @      "@      0@      $@      "@      ;@      "@      @      7@      A@     @Q@      �?      @      .@      "@      @      *@      �?      1@       @       @               @      @      @      @       @      @      (@     �A@                      @      @      @      *@      @      ?@      @      @      0@       @      @      6@      @      @      4@      6@      A@      �?      @       @      @      @      �?      @      ,@      @       @      @      @      �?      "@      @      *@      1@       @       @      @      .@      $@      @      @              @       @                      @      @              @              @      @              @              @       @      @       @              @       @                       @      �?              @              @      �?              �?              @              �?      �?                                              �?      @                              �?      @              @                       @       @      �?      �?      �?      (@      @       @      �?       @      �?      @      @      @      *@       @      @      @      $@       @       @      @              �?      @               @                      �?      @                      @       @      �?                      �?                      �?               @      @      @      �?       @               @      @      @       @              @      @      $@      @       @      @     �f@      :@     �Z@      5@      7@      @      ;@     �l@     �m@      5@      8@      L@     Pp@      b@      "@      3@      3@     �N@      @     @Q@      @      ;@      @      @              @      b@      `@      @      @      *@     �W@      I@              @       @      ,@       @      <@      �?      ,@      @      @               @      G@     �P@              @      @     �D@      3@                      �?      @               @              �?      �?                      �?      (@     �A@                      �?      $@       @                               @                                                                      �?      ,@                              @                                                       @              �?      �?                      �?      &@      5@                      �?      @       @                               @              4@      �?      *@       @      @              �?      A@      @@              @      @      ?@      1@                      �?      @                              �?              �?                      �?                       @              @                                                      4@      �?      (@       @       @              �?     �@@      @@              �?      @      :@      1@                      �?      @             �D@      @      *@       @                      @     �X@     �N@      @      @       @     �J@      ?@              @      �?      "@       @      *@                                                      @      @                              @      @                                              �?                                                       @      @                               @       @                                              (@                                                      �?      �?                              �?      �?                                              <@      @      *@       @                      @      X@      L@      @      @       @      I@      <@              @      �?      "@       @      3@               @                               @     @S@     �@@      @      �?      @      D@      5@                              @       @      "@      @      @       @                      @      3@      7@              @      �?      $@      @              @      �?      @              \@      5@     �S@      0@      4@      @      4@     @U@     �[@      2@      1@     �E@     �d@     �W@      "@      .@      1@     �G@      @      G@      @      9@      �?      @              @      J@      K@      @      (@      @      T@     �E@              @      @      5@       @      9@      @      @      �?      @              �?      (@      1@       @      @      @      D@      2@                      �?      "@      �?      5@      @      @      �?      @              �?      $@      0@      �?      �?      @     �C@      0@                      �?      "@      �?      @                              �?                       @      �?      �?      @      �?      �?       @                                              5@       @      3@              @               @      D@     �B@      @      @              D@      9@              @      @      (@      �?      2@       @      (@              @               @     �C@     �B@      @      @              D@      7@              �?      @      (@      �?      @              @                                      �?                                               @              @                             �P@      0@      K@      .@      *@      @      1@     �@@     �L@      (@      @     �B@     �U@     �I@      "@      $@      *@      :@      @      8@              7@      "@               @      @      "@       @      @              @      ,@      "@              �?      @                      7@              6@       @                      @      "@      @       @               @      &@       @              �?                              �?              �?      �?               @                      �?      �?               @      @      �?                      @                      E@      0@      ?@      @      *@      �?      ,@      8@     �H@      "@      @     �@@     @R@      E@      "@      "@       @      :@      @      ?@      @      5@      @      "@              "@      5@      F@      "@      @      3@     �M@      8@      @       @       @      4@       @      &@      "@      $@       @      @      �?      @      @      @                      ,@      ,@      2@      @      �?      @      @      �?�t�bub��     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJo�vhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmK]hnh4h7K ��h9��R�(KK]��hu�BX         6                    �?�{��ؙ�?�	           ��@                           @2��TP��?Y           L�@                           �?L���N�?M           `�@                           �?[����~�?�             s@                          �2@f4I��N�?;            �V@                          �1@
^N��)�?             <@������������������������       �/k��\�?             1@������������������������       �F]t�E�?             &@	       
                     �?��A���?'            �O@������������������������       ���\���?
             1@������������������������       �UA�>�)�?             G@                            @������?�            �j@                           �?�\�����?Z            @_@������������������������       �;�;��?(             J@������������������������       �L���?2            @R@                          �:@�����|�?6             V@������������������������       �̥-����?-            �R@������������������������       �؉�؉��?	             *@                          �3@�X�֌�?�           ��@                           @��� ]�?�            �h@                           �?�+.�k�?z            �f@������������������������       ��q�q�?$             H@������������������������       �E������?V            �`@������������������������       �     ��?	             0@                            @Zyv�7��?�            Py@                            �?�`�:k��?�            `m@������������������������       �6��`�?G            �]@������������������������       ��7+���?J            @]@                           �?�{E٢�?n            @e@������������������������       ��M,�7��?            �A@������������������������       ������?W            �`@        )                   �1@����P��?           8�@!       (                    @�M��t~�?o             g@"       %                    @n��Q�?i            �e@#       $                    @t��kl�?L             _@������������������������       �9%�R�@�?!             K@������������������������       �����L�?+            �Q@&       '                     �?NMM�?            �H@������������������������       ��$�_�?             3@������������������������       ��������?             >@������������������������       �9��8���?             (@*       1                   �8@�t�>g�?�           p�@+       .                    @�6WM���?P           ��@,       -                    @����F��?6           0~@������������������������       �����+O�?�             j@������������������������       ���E�?�             q@/       0                     @��2Tv�?            �F@������������������������       �a��V{q�?             ?@������������������������       �
^N��)�?             ,@2       5                   �=@�¿��?M            �_@3       4                    �?��D����?B            �Z@������������������������       �;U��j�?             =@������������������������       �*�z4:�?0            @S@������������������������       ��Q����?             4@7       J                   �5@~Gq�R��?G           �@8       G                    @���,�?�           ,�@9       @                   �1@$��N/$�?�           А@:       =                     �?`!�2���?�            �q@;       <                    �?R�=�U��?1            �T@������������������������       ����Դ�?             3@������������������������       �     ��?%             P@>       ?                    �?����z
�?�            �h@������������������������       �3�R�f�?2             S@������������������������       ��/�K.��?Y            �^@A       D                    @�w�e�?�           Ј@B       C                    �?�)G/��?5           `@������������������������       �5]���?�            @l@������������������������       �=b����?�            @q@E       F                    �?{G0�ˡ�?�            @r@������������������������       �lykl���?L            �\@������������������������       �d���3�?n            @f@H       I                     �?K����?             7@������������������������       ���"e���?             "@������������������������       ��)x9/�?             ,@K       Z                    @�B6W�?�           ��@L       S                    @��	jP�?�           \�@M       P                     �?��<���?�           (�@N       O                    �?�Žf�@�?�            @y@������������������������       ����6�?Q            @b@������������������������       ���n�H��?�             p@Q       R                   �@@݇�s�?�            s@������������������������       �1rq�RW�?�            `r@������������������������       �b���i��?             &@T       W                    @8����x�?�             u@U       V                    �?_��+��?b            �d@������������������������       ���s�؟�??            @Z@������������������������       �J��8���?#             O@X       Y                    @K�W#&�?u            `e@������������������������       �~")d�?0            @T@������������������������       ���M1j��?E            �V@[       \                     �?{�G�z�?             4@������������������������       �9��8���?             (@������������������������       �      �?              @�t�bh�h4h7K ��h9��R�(KK]KK��h��B87        }@     �S@     pt@     �H@     �S@      ?@      X@     @�@      �@      Q@     �Q@     �b@     ��@     `{@      "@     �P@     �F@     @^@     �P@     �i@      @@     �]@      &@      3@      "@     �C@     �u@     0u@      9@      7@     �L@     0q@     �d@       @      8@      (@      >@      2@     �^@      .@     �R@      "@      $@      "@      8@     �]@      b@      &@      &@     �C@     �d@     �U@       @      4@      "@      1@      1@     �L@      @      1@              �?              @      @@     �O@      @      @      .@      M@      ;@      �?      @      �?      @      @      .@       @      @                                       @      ?@       @      �?      @      &@      @              �?      �?      �?       @      (@              @                                      @      @      �?              �?               @              �?                              @               @                                      @       @      �?              �?              �?                                              @              �?                                      �?       @                                      �?              �?                              @       @       @                                      @      ;@      �?      �?      @      &@      @                      �?      �?       @                                                                      $@                              @                              �?                      @       @       @                                      @      1@      �?      �?      @      @      @                              �?       @      E@      @      (@              �?              @      8@      @@      �?       @      $@     �G@      5@      �?      @              @       @      7@       @      "@              �?              @      3@      2@      �?       @      "@      8@      @               @               @              $@              @              �?              @      @       @              �?      @      (@      @               @               @              *@       @      @                                      *@      0@      �?      �?      @      (@      @                                              3@       @      @                                      @      ,@                      �?      7@      ,@      �?       @               @       @      ,@              �?                                      @      ,@                      �?      6@      *@      �?                       @       @      @       @       @                                                                              �?      �?               @                             �P@      "@      M@      "@      "@      "@      2@     �U@     �T@       @       @      8@     @[@     �M@      �?      .@       @      (@      *@      =@      �?      @                              �?      I@     �E@      @              @     �C@      (@               @               @      @      =@      �?      @                              �?      I@      C@       @              @      A@      (@                               @      @      @              �?                                      *@      "@       @               @      $@      @                                              9@      �?      @                              �?     �B@      =@                       @      8@      @                               @      @                      �?                                              @      �?               @      @                       @                             �B@       @     �I@      "@      "@      "@      1@     �B@     �C@      @       @      2@     �Q@     �G@      �?      *@       @      $@      "@      ?@      @      B@              @              $@      ;@      ,@      @      @      @      B@      9@              "@      @       @      @      3@      @      2@                              @      @      @       @      @       @      6@      (@              @               @       @      (@       @      2@              @              @      6@       @      @      @      @      ,@      *@              @      @              @      @      �?      .@      "@      @      "@      @      $@      9@              �?      &@      A@      6@      �?      @      @       @      @                      �?                      @      �?      @      "@                      �?       @       @              �?      �?               @      @      �?      ,@      "@      @      @      @      @      0@              �?      $@      :@      4@      �?      @      @       @       @     �T@      1@     �E@       @      "@              .@     @l@     @h@      ,@      (@      2@      [@     �S@              @      @      *@      �?      2@      �?      @                               @     �T@      I@                      @      4@       @                                              *@      �?      @                               @     �S@      I@                      @      1@       @                                              @      �?      @                                      O@      >@                      @      0@                                                      @      �?      @                                      3@      .@                       @      "@                                                      �?              @                                     �E@      .@                      �?      @                                                      @                                               @      1@      4@                              �?       @                                                                                               @      @      (@                              �?                                                      @                                                      *@       @                                       @                                              @                                                      @                                      @                                                      P@      0@     �B@       @      "@              *@     �a@      b@      ,@      (@      .@      V@      S@              @      @      *@      �?      H@      @      =@              @              "@     �^@     �_@      (@      @      $@     �Q@     @Q@              @      @      $@             �F@      @      ;@              @              @      Z@      ^@      &@      @      $@     �O@     @Q@              @       @      $@              3@      @      2@                              @      E@     �F@      @      @      "@     �B@      4@                      �?      �?              :@       @      "@              @                      O@     �R@      @       @      �?      :@     �H@              @      �?      "@              @               @                              @      2@      @      �?                       @                              �?                      @              �?                                      .@      @      �?                      @                              �?                                      �?                              @      @       @                              @                                                      0@      $@       @       @      @              @      5@      1@       @      @      @      1@      @                              @      �?      (@      $@      @       @      @              @      5@      0@      �?      @      @      &@      @                              @      �?      @      �?                                      @      @      &@              �?       @      �?       @                                               @      "@      @       @      @                      2@      @      �?      @      @      $@       @                              @      �?      @              @               @                              �?      �?                      @      @                                             Pp@      G@      j@      C@     �M@      6@     �L@     �i@     �p@     �E@      H@      W@      t@      q@      @      E@     �@@     �V@      H@     �c@      0@     @Z@      $@      *@      �?      6@      d@     �h@      @      0@     �C@     �b@     @`@               @      &@     �D@      1@      c@      0@     �Y@      $@      *@      �?      3@     �c@     �h@      @      0@     �C@     `b@     �^@               @      &@     �D@      ,@     �B@       @      .@              @               @     �O@      R@              @      "@     �B@      9@                       @      @      @       @      �?      �?                               @      2@      <@               @      @      $@      @                                      �?                                                       @      @      @                       @      @       @                                               @      �?      �?                                      *@      9@               @      @      @      @                                      �?      =@      �?      ,@              @                     �F@      F@              @      @      ;@      2@                       @      @       @      3@      �?      @              �?                      @      .@              �?      @      "@      @                       @      @       @      $@              @               @                      C@      =@              @      �?      2@      (@                              @              ]@      ,@      V@      $@      $@      �?      1@      X@     @_@      @      $@      >@     �[@     �X@               @      "@     �A@      &@     @U@       @      I@      @      @      �?      ,@     �P@     @R@      @      @      (@     �R@     �R@              @      @       @      @      A@      @      9@      @      @      �?      @      0@      B@              @       @      =@      F@              �?      @      @             �I@      �?      9@       @      @              "@     �I@     �B@      @       @      @      G@      >@              @       @      �?      @      ?@      @      C@      @      @              @      =@      J@      @      @      2@     �A@      8@              @      @      ;@      @      1@      �?      ;@              �?               @      @      &@       @      �?      &@      0@      @                       @      &@      @      ,@      @      &@      @       @              �?      :@     �D@      �?      @      @      3@      2@              @       @      0@       @      @               @                              @      �?                                       @      @                                      @                       @                                      �?                                              @                                      @      @                                              @                                               @      @                                             �Y@      >@      Z@      <@      G@      5@     �A@     �G@      R@     �B@      @@     �J@     `e@      b@      @      A@      6@      I@      ?@     �X@      >@     �X@      6@      G@      5@     �A@      G@      R@     �B@      >@     �J@     `e@      b@      @     �@@      6@      I@      ?@     @P@      3@      O@      1@      E@      5@      ;@      :@      D@      :@      8@     �B@     �W@     �Y@      @      9@      0@      =@      =@     �E@       @     �C@      @      3@      $@      5@      0@      (@      .@      1@      1@     @R@     �G@      @      .@      (@      3@      *@      .@      @      (@              $@      �?      &@       @      @       @      @      @     �C@      *@              @       @      @      @      <@      @      ;@      @      "@      "@      $@       @      @      *@      &@      (@      A@      A@      @      (@      $@      .@      @      6@      &@      7@      (@      7@      &@      @      $@      <@      &@      @      4@      6@     �K@      @      $@      @      $@      0@      6@      &@      6@      (@      7@      &@      @      $@      <@      $@      @      3@      6@     �K@              $@      @      $@      (@                      �?                                                      �?              �?                      @                              @      A@      &@      B@      @      @               @      4@      @@      &@      @      0@      S@      E@               @      @      5@       @      7@      @      6@      @      �?              �?      $@      5@       @      @      @      5@      6@               @      @      @      �?      3@      @      @              �?              �?      @      ,@      @      @      @      (@      0@              @      @       @      �?      @       @      0@      @                              @      @       @                      "@      @              @      �?      @              &@      @      ,@      �?      @              @      $@      &@      @       @      &@     �K@      4@                       @      0@      �?      �?      @      @      �?                      �?      @      @      @       @      @     �@@      @                              "@              $@      �?      "@              @              @      @      @                      @      6@      *@                       @      @      �?      @              @      @                              �?                       @                                      �?                               @              @      @                              �?                      �?                                      �?                               @               @      @                                                      �?                                                                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��1QhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmK}hnh4h7K ��h9��R�(KK}��hu�BX         >                   �3@��~�я�?�	           ��@                           @�.�I���?\           @�@                            @�@���?�           ��@                           �?gȧ�0�?�            �w@                          �0@Iy��	:�?p            @e@                            �?����S�?             <@������������������������       ��h$���?
             .@������������������������       ��	j*D�?             *@	       
                    @�_���?^            �a@������������������������       �K`ݞ��?J            @\@������������������������       �΃�\W�?             =@                           �?@0��>�?�            @j@                            �?��paR�?W             a@������������������������       ��?*             Q@������������������������       �=[y���?-             Q@                           @�^���B�?.            �R@������������������������       ��BR�8�?             C@������������������������       �6?,R��?             B@                           �?���n��?�            �o@                          �2@`��6��?I            �\@                          �1@��5�X�??            �Y@������������������������       �IPS!���?              J@������������������������       ��&�W�?             I@������������������������       ��������?
             (@                           @��P�Y�?_            @a@                          �2@Z��Z���?)            @P@������������������������       �k�w��#�?             I@������������������������       �hE#߼�?             .@                           @�2��	a�?6            @R@������������������������       ��#��Z=�?             6@������������������������       ���X���?$            �I@        /                    @�]�ط�?�           ��@!       (                     @��H��?D           h�@"       %                    @ڃ����?           �z@#       $                    @8�RY�l�?�            �k@������������������������       �7�3��?E             [@������������������������       �6��|r�?A            �\@&       '                   �0@�kd#���?~            �i@������������������������       �Cu��?             E@������������������������       �OK���V�?e            `d@)       ,                    @���ˈ�?@            �X@*       +                   �2@M=ֱ߹�?$            �L@������������������������       ��I��k��?            �F@������������������������       �r�q��?             (@-       .                   �2@�&q	�X�?            �D@������������������������       �R����?            �@@������������������������       �      �?              @0       7                     �?����	�?{            `i@1       4                   �1@�~�u�7�?1            �U@2       3                    �?      �?             B@������������������������       �䃞ͪ��?             9@������������������������       ���!pc�?             &@5       6                    �?�t.��?            �I@������������������������       ���>4և�?             ,@������������������������       ���0\K5�?            �B@8       ;                    �?[-��p�?J             ]@9       :                     @����I��?$            �K@������������������������       �̄���?            �D@������������������������       �������?	             ,@<       =                    �?�x/^���?&            �N@������������������������       �J��LQ�?             7@������������������������       ����Դ�?             C@?       ^                    �?e~Ѡ�?5           �@@       O                    �?U%��-X�?�           ��@A       H                    �?���Ǜ�?�            �t@B       E                   �9@�P�7���?M            �_@C       D                    �?�w��&��?5            �T@������������������������       �(&ޏ��?             F@������������������������       �������?            �C@F       G                     �?V#��?            �E@������������������������       �����X�?             ,@������������������������       �:2��h�?             =@I       L                     @ƵHPS��?�             j@J       K                     �?��e]��?H            �Z@������������������������       ��D�M��?&            �K@������������������������       �|���t��?"             J@M       N                   �4@B=�����?@            @Y@������������������������       ��zv��?             6@������������������������       �k�*��?3            �S@P       W                    �?[���mV�?           ��@Q       T                    �?Kz^4���?�            0u@R       S                    @������?F            @Z@������������������������       ����!pc�?             6@������������������������       ���c�6�?9            �T@U       V                    @�%�u��?�            @m@������������������������       ���0\K5�?            �B@������������������������       �������?|            �h@X       [                   �?@��4�!z�?F            �@Y       Z                   �4@Ae6#P9�?'           �|@������������������������       ���?�(�?              J@������������������������       �����f�?           �y@\       ]                   @A@���s��?            �K@������������������������       �#>�֕�?            �A@������������������������       ���(\���?             4@_       n                    @�$2Hw�?C           P�@`       g                    �?)�`�J:�?�            �w@a       d                   �5@����_��?b             d@b       c                    �?��>4և�?              L@������������������������       �     ��?             @@������������������������       ��q�q�?             8@e       f                     �?���y�F�?B            @Z@������������������������       �     ��?             @@������������������������       �*c����?/            @R@h       k                    @ �t�Vl�?�            @k@i       j                     �?U$	��$�?{            �h@������������������������       ���Moz��?*            @Q@������������������������       ����G��?Q             `@l       m                   �7@��Q���?             4@������������������������       ���"e���?             "@������������������������       �j�V���?             &@o       v                   �8@�tN�m�?X           Ȏ@p       s                     @������?�           �@q       r                    �?X/se���?g           P�@������������������������       �V�Z��?�            0q@������������������������       ��0	�\�?�            ps@t       u                    �?O�b����?H            �\@������������������������       ��k��(A�?%            �M@������������������������       ��$I�$I�?#             L@w       z                   �9@������?�            �q@x       y                    @
�~�n[�?'            @P@������������������������       ���Er��?             A@������������������������       �N�s�-�?             ?@{       |                    @�J�5� �?�            `k@������������������������       ��z�G��?F             ^@������������������������       ���M=-�?<            �X@�t�bh�h4h7K ��h9��R�(KK}KK��h��B8J       Py@     �W@     v@      9@     @R@      :@     @T@     �@     ��@     @S@      V@     �d@     H�@     �y@      1@     �P@      L@     @[@      J@      d@      1@      U@      @      @              (@     �u@     pp@      0@      *@     �C@     �n@     �Z@              "@      @      <@       @     @V@      "@     �E@       @      @              @      Z@      [@      "@      @      8@     �`@      L@              @      @      5@       @      M@      �?      9@      �?       @              @     �R@      U@      @      @      0@      Q@      :@               @      �?      @      @      =@      �?      $@                                      G@      D@       @      @      @      5@      @                              @      �?      �?                                                      "@      ,@               @               @                                                      �?                                                      @      @               @               @                                                                                                              @      "@                                                                                      <@      �?      $@                                     �B@      :@       @       @      @      3@      @                              @      �?      2@      �?       @                                      @@      5@              �?      @      .@      @                              @      �?      $@               @                                      @      @       @      �?              @                                                      =@              .@      �?       @              @      =@      F@       @              $@     �G@      3@               @      �?      @      @      6@              @      �?       @               @      *@      9@       @              $@     �@@      *@              �?              @      @      (@              @      �?                      �?       @      "@                      @      5@      $@                                              $@              @               @              �?      @      0@       @              @      (@      @              �?              @      @      @              "@                              �?      0@      3@                              ,@      @              �?      �?                       @              @                              �?      $@       @                              (@      @              �?                              @              @                                      @      1@                               @                              �?                      ?@       @      2@      �?      @               @      =@      8@      @       @       @     @P@      >@              @       @      .@      @      0@       @      @                               @      3@      &@      @              @      A@      *@              �?              @      �?      0@       @       @                               @      1@      $@      @              �?      @@      &@              �?              @              $@               @                                      "@      @      @              �?      0@      @                                              @       @                                       @       @      @                              0@      @              �?              @                              �?                                       @      �?                      @       @       @                                      �?      .@      @      .@      �?      @                      $@      *@       @       @      @      ?@      1@               @       @      $@      @      @      @       @              @                      @      @              �?      @      6@       @              �?              �?              @      @      @               @                      @      @                      @      4@      �?                                               @              @              @                                              �?               @      �?              �?              �?              "@       @      @      �?                              @      @       @      �?      �?      "@      .@              �?       @      "@      @      @      �?      @      �?                              @       @              �?              �?      @                                              @      �?      @                                      �?      @       @              �?       @      &@              �?       @      "@      @      R@       @     �D@       @                      @      n@     `c@      @      @      .@      \@      I@              @      �?      @              E@      @      <@      �?                      @      h@      \@      @      @      $@      U@     �@@                               @              ?@      @      &@                               @      f@      X@      @      @      @     �O@      9@                               @              3@      @      @                                     @[@      E@      @      �?      @      7@      (@                                              ,@      @       @                                      E@      5@      @      �?              *@      @                                              @              @                                     �P@      5@                      @      $@      @                                              (@              @                               @     �P@      K@      @      @      �?      D@      *@                               @              @                                                      5@      &@                              @      �?                                              @              @                               @      G@     �E@      @      @      �?      B@      (@                               @              &@              1@      �?                      �?      0@      0@              �?      @      5@       @                                               @              ,@      �?                      �?      @      "@                       @      1@      @                                               @              ,@                              �?      @      @                       @      0@                                                                              �?                               @       @                              �?      @                                              "@              @                                      &@      @              �?      @      @       @                                              "@              �?                                      &@      @                      �?      @       @                                                               @                                               @              �?      @                                                              >@      @      *@      �?                      @      H@     �E@              �?      @      <@      1@              @      �?      @              $@      @      @      �?                      @      3@      0@                      @      2@      @                      �?      @              @              �?                                      $@      @                      @      *@                                                                      �?                                       @       @                      @      &@                                                      @                                                       @      �?                               @                                                      @      @      @      �?                      @      "@      *@                      �?      @      @                      �?      @               @                                              @              @                                      @                                               @      @      @      �?                              "@      @                      �?      @                              �?      @              4@              @                              �?      =@      ;@              �?      �?      $@      ,@              @               @              @              @                                      4@      (@              �?              @      "@                                              @              �?                                      1@      &@                               @      @                                                               @                                      @      �?              �?              �?      @                                              *@              @                              �?      "@      .@                      �?      @      @              @               @              "@              @                                      @      �?                              @       @                                              @                                              �?      @      ,@                      �?      @      @              @               @             �n@     @S@     �p@      5@     �P@      :@     @Q@     �l@     �t@     �N@     �R@     �_@     @y@     �r@      1@     �L@      J@     @T@      F@     �]@      E@     `b@      "@      I@      5@     �A@     �J@     �[@      B@      G@     @P@     `c@     `c@      @     �@@      A@     �C@      A@     �K@      $@      A@      �?      2@      @      @      ,@     �E@      @      ,@      2@      C@     �B@       @      (@      "@      @      @      *@      @      @               @              �?      @      :@      @      (@      @      0@      (@              @      @      �?      @      "@      @      @                                      @      8@      @      @      @      $@      @              @      �?      �?      @      @      @       @                                       @      .@       @      �?              @      �?              @              �?      @      @               @                                      @      "@      �?      @      @      @       @                      �?              �?      @      @       @               @              �?               @               @              @      "@              @       @                      @                              �?                               @              @              @                               @                      �?      @       @              �?              �?                              @              @      "@              @                              E@      @      <@      �?      0@      @      @       @      1@      @       @      &@      6@      9@       @      @      @      @       @      <@      �?      0@              @              @      @      @       @      �?      @       @      0@       @               @      @              *@              @               @                       @      @      �?              @      @      "@       @               @      @              .@      �?      "@              �?              @      @       @      �?      �?      @       @      @                                              ,@       @      (@      �?      *@      @              �?      $@      �?      �?      @      ,@      "@              @      @       @       @      @      �?                      @                      �?                                      @      @                                              $@      �?      (@      �?      @      @                      $@      �?      �?      @      $@      @              @      @       @       @     �O@      @@     @\@       @      @@      .@      >@     �C@      Q@      >@      @@     �G@     @]@     �]@      @      5@      9@     �@@      <@      :@       @     �D@       @      &@      @      &@      7@     �@@      @      "@      2@     �M@      H@              @      (@      *@      (@      $@              &@               @      �?       @      $@      &@      @       @      @      6@      *@               @       @      @      @      �?               @                                       @      �?      @               @      @                      �?                              "@              @               @      �?       @       @      $@               @      @      2@      *@              �?       @      @      @      0@       @      >@       @      "@       @      "@      *@      6@              @      &@     �B@     �A@              @      $@      $@       @      @              @                               @       @       @                      @              "@              @              @              *@       @      8@       @      "@       @      @      &@      4@              @      @     �B@      :@               @      $@      @       @     �B@      8@      R@      @      5@      (@      3@      0@     �A@      ;@      7@      =@      M@     �Q@      @      ,@      *@      4@      0@      B@      8@     @Q@      @      2@      @      3@      0@      ?@      3@      5@      1@      M@      Q@              *@      (@      2@      &@      @              &@                                       @      @                       @      3@      @                              �?       @      ?@      8@      M@      @      2@      @      3@      ,@      <@      3@      5@      .@     �C@     �N@              *@      (@      1@      "@      �?              @       @      @      @                      @       @       @      (@               @      @      �?      �?       @      @      �?              @      �?      @      @                               @              @               @              �?      �?       @      �?                              �?                                      @               @      @                      @                              @     �_@     �A@     �^@      (@      0@      @      A@      f@     �k@      9@      =@     �N@      o@     `b@      &@      8@      2@      E@      $@      ?@      .@      =@      @      @      @      *@      8@     @R@       @      @      ,@     @R@      K@      �?      @              (@      @      3@       @      *@       @                      �?      1@      B@      �?      @      @      >@      5@              @                              @      @       @                                      @      4@                              .@      @                                              @      @                                              @      1@                              @       @                                              @               @                                      @      @                              &@      �?                                              (@      @      &@       @                      �?      &@      0@      �?      @      @      .@      2@              @                              �?      @      @                              �?      @      $@              �?       @      @       @                                              &@       @       @       @                              @      @      �?       @      @      $@      0@              @                              (@      @      0@       @      @      @      (@      @     �B@      @      @       @     �E@     �@@      �?       @              (@      @      $@      @      (@       @      @      @      $@      @     �B@      @      @       @      D@      @@      �?                      &@      @      @              "@      �?              �?      @      @      "@      �?      @       @      2@      @                              @       @      @      @      @      �?      @      @      @      @      <@      @              @      6@      9@      �?                      @       @       @              @              @               @                              �?              @      �?               @              �?                              @               @              �?                                              @                                                       @              �?               @              �?                              �?                      �?               @              �?             �W@      4@     @W@       @      "@      �?      5@      c@     �b@      1@      6@     �G@      f@     @W@      $@      2@      2@      >@      @     �S@      @      K@      @      @              $@      _@     �]@      @      $@      A@     @_@     �Q@      "@      &@      "@      7@      @     �O@      @      F@      @       @              $@      \@     �Z@      @      "@      <@     �X@     �J@      @      &@      @      3@      @      >@      �?      1@                              @      O@     �P@      @      @      @     �C@      <@              @      �?      @             �@@       @      ;@      @       @              @      I@      D@      �?      @      6@      N@      9@      @       @      @      (@      @      0@      �?      $@              �?                      (@      (@      �?      �?      @      :@      1@      @               @      @               @              @                                      $@      @      �?      �?              3@       @                       @      @              ,@      �?      @              �?                       @      @                      @      @      "@      @                                      0@      0@     �C@      �?      @      �?      &@      <@      >@      &@      (@      *@     �I@      7@      �?      @      "@      @       @      @      @      @                              @      @      @      @      @      @      5@       @               @      �?       @               @              @                              @      �?      @      @      @      �?      @                       @      �?       @              �?      @      �?                              �?      @                               @      1@       @                                              *@      (@      A@      �?      @      �?      @      8@      ;@      @      @      $@      >@      5@      �?      @       @      @       @      @      $@      9@              �?      �?      @      *@       @      @      @      @      ,@      @      �?      @       @      @       @      @       @      "@      �?      @              @      &@      3@       @      @      @      0@      .@                              �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�
hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         :                   �3@Om�}Ǧ�?�	           ��@                           �?h�"�?           P�@                          �1@�7'�K�?�           h�@                           @��	"P7�?�             s@                            @k8�{F�?�            q@                           �?��Dp2h�?�            �i@������������������������       ��c�1��?             ?@������������������������       ���x���?s            �e@	       
                    �?"�O�|�?-             Q@������������������������       �
���?            �@@������������������������       �ۨ:�.�?            �A@������������������������       ��d�ۇ��?             ?@                           @�����?�            �w@                            @�ejd��?k            @f@                           @HɶZ���?<            �X@������������������������       ����t�?"            �M@������������������������       �>
ףp=�?             D@                           �?���8��?/            �S@������������������������       ��^��T�?             =@������������������������       ���|?5^�?             I@                            �?��P��?~            `i@                          �2@@�'�@��?             C@������������������������       �{�G�z�?             4@������������������������       ������H�?             2@                          �2@���R���?d            �d@������������������������       ��|Z
���?1            �W@������������������������       �RMw���?3            �Q@       +                    @nHF�6��?�           8�@       $                    @n3����?#           @}@       !                   �2@�{�I���?�            �t@                           �0@{�p�]�?�            `m@������������������������       ���Q0�x�?            �E@������������������������       �UUUUU��?y             h@"       #                    @ށ����?<            �X@������������������������       �`�Q��?1            �R@������������������������       �J��LQ�?             7@%       (                     @�&�co��?X            �`@&       '                   �0@=��G��?8            �T@������������������������       �������?             ,@������������������������       �� =[y�?0             Q@)       *                   �2@�+ Wd�?             �J@������������������������       �f��E�?            �B@������������������������       �     ��?
             0@,       3                    @b9���n�?�            0q@-       0                    @X��W��?w            @g@.       /                     @d_� H�?Z            �`@������������������������       ���ښ��?G            @Z@������������������������       �[�[��?             >@1       2                   �1@��X�w�?            �I@������������������������       ��Q�}e�?             :@������������������������       ���JY�8�?             9@4       7                    @%L���x�?8            @V@5       6                   �2@N�zv�?            �@@������������������������       �<ݚ�?
             2@������������������������       �t�@�t�?             .@8       9                    @s
^N���?#             L@������������������������       �P7�Z�?             C@������������������������       �<ݚ�?
             2@;       T                   �7@�&��h�?           j�@<       K                    @�{7s�?>           ��@=       D                    �?��GJh�?�           ��@>       A                     �?��c����?o           p�@?       @                   �4@�an�D�?�            `u@������������������������       �"n����?>            @Z@������������������������       � ���B�?�            �m@B       C                   �6@� ����?�             o@������������������������       �Tc�W��?            `i@������������������������       �!����?!            �F@E       H                    �?���'��?�           ��@F       G                   �4@�"����?�            �j@������������������������       �z$�J0c�?*            @P@������������������������       �(\A��?`            �b@I       J                   �4@ܮ����?�            �y@������������������������       �     ��?P             `@������������������������       �B����#�?�            �q@L       S                    !@S�f��?K            �\@M       P                    @��+�J-�?E            �Y@N       O                   �5@[�[��?.            �R@������������������������       ����J�?             F@������������������������       ��η���?             ?@Q       R                   �4@T�r
^N�?             <@������������������������       ��������?	             (@������������������������       �      �?             0@������������������������       ��zv��?             &@U       d                    @1��v�?�           �@V       ]                     @�� ��?�           ��@W       Z                   �?@����Π�?8           p~@X       Y                    �?��m����?            {@������������������������       ��4����?V            ``@������������������������       �H�]aZ��?�            �r@[       \                    �?�:��R�?#            �J@������������������������       �s
^N���?             ,@������������������������       �y�*3��?            �C@^       a                    �?mvq`��?�             s@_       `                   �8@�ۏ��?G            �^@������������������������       �(N:!���?            �A@������������������������       ���a��Y�?5            �U@b       c                    @ٝ�����?v            �f@������������������������       �X��|�`�?l             e@������������������������       ���>4և�?
             ,@e       l                    @L�f���?�            �v@f       i                    @� �����?\            �c@g       h                     �?I��M�z�?<            �Y@������������������������       �x�����?!             M@������������������������       �
�d�j��?            �F@j       k                     @�b-����?             �J@������������������������       �"�O�|�?             A@������������������������       ��}�+r��?
             3@m       p                   �?@0-��l�?�            @j@n       o                    @UUUUUI�?w             h@������������������������       �;h�r�?c            �c@������������������������       �]�l� �?             A@q       r                    @�E��ӭ�?             2@������������������������       �������?             @������������������������       �*L�9��?             &@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       |@     �X@     0u@     �@@     �S@      =@     @U@     ��@     �@      S@     �T@     �d@     P�@     0{@      @      O@     �K@     �`@      I@     `d@      1@      Y@      @      @              1@      v@     �q@      &@      4@      D@     �k@     @_@              .@      @      C@      @      T@      @     �@@      �?                      @     �k@     �`@      @      @      4@     �X@      J@              @              0@       @      C@      @      *@                              �?     �]@      R@      @       @      "@     �B@      @                                             �B@      @      (@                              �?      Z@     �P@      @       @      @     �@@      @                                              ;@      @      @                              �?     �U@     �I@               @      @      6@      @                                              @              @                                      $@      "@                      �?      @      �?                                              8@      @       @                              �?      S@      E@               @      @      3@       @                                              $@              @                                      2@      0@      @              �?      &@      @                                              @              @                                      (@      @       @              �?      �?      �?                                              @               @                                      @      $@      �?                      $@       @                                              �?              �?                                      .@      @                      @      @      �?                                              E@      @      4@      �?                      @     @Y@      O@      @      @      &@     �N@     �F@              @              0@       @      :@      @      @                                      B@      :@               @       @      =@      6@              @              *@       @      4@      �?      @                                      7@      .@               @      @      0@      @                               @               @      �?      @                                      .@      ,@               @       @      &@      @                              @              2@                                                       @      �?                       @      @       @                              @              @      @      �?                                      *@      &@                      @      *@      0@              @              @       @      @      @                                                      @                              �?       @              @              @              �?              �?                                      *@      @                      @      (@       @               @              �?       @      0@              .@      �?                      @     @P@      B@      @      @      @      @@      7@                              @              @                      �?                              @      *@      �?              �?      $@      @                                              �?                                                       @      &@                              @      @                                               @                      �?                               @       @      �?              �?      @       @                                              *@              .@                              @     �N@      7@       @      @       @      6@      2@                              @              @              $@                                     �F@      (@      �?                      *@      $@                                              "@              @                              @      0@      &@      �?      @       @      "@       @                              @             �T@      $@     �P@      @      @              *@     �`@     �b@      @      *@      4@     �^@     @R@              $@      @      6@      @     �M@      @      H@      @      @               @      N@      S@      @      (@      (@      V@     �M@              @      @      0@      @      G@      @      ;@       @      @              @      H@     �H@      @      &@      &@     @R@     �B@              @       @      @       @      >@      @      .@               @              @      @@     �A@      @      @      "@      O@      8@              �?       @      @      �?      (@      �?                                              @      @                              ,@      @                                              2@      @      .@               @              @      :@      <@      @      @      "@      H@      5@              �?       @      @      �?      0@              (@       @      �?                      0@      ,@              @       @      &@      *@               @              @      �?      &@              (@       @      �?                      ,@      @               @       @      @      *@               @              @      �?      @                                                       @       @              @              @                                                      *@              5@      �?      @              @      (@      ;@       @      �?      �?      .@      6@                      �?      $@      �?      @              .@              �?              @      $@      8@      �?              �?      $@      @                               @      �?      �?                                                      �?      &@                              �?                                                      @              .@              �?              @      "@      *@      �?              �?      "@      @                               @      �?       @              @      �?       @                       @      @      �?      �?              @      .@                      �?       @              @              @               @                       @      �?              �?               @      &@                              @              �?                      �?                                       @      �?                      @      @                      �?      @              8@      @      3@      @                      @     �R@      R@              �?       @      A@      ,@              @      @      @      �?      6@       @      *@                              @      J@     �J@                              9@      "@              @      �?                      4@       @      &@                              @     �B@      @@                              .@      "@              @      �?                      .@       @      @                              �?     �A@      >@                              "@      @               @      �?                      @              @                              @       @       @                              @      @               @                               @               @                              �?      .@      5@                              $@                                                       @              �?                                      @      *@                              @                                                                      �?                              �?      $@       @                              @                                                       @      �?      @      @                              6@      3@              �?       @      "@      @              @      @      @      �?              �?      @      @                              @      @              �?      @      @                       @              �?      �?                                                              @       @                      @      @                       @                      �?              �?      @      @                              �?      @              �?              �?                                      �?               @               @                                      2@      ,@                       @      @      @              �?      @      @               @               @                                      ,@       @                              @       @              �?      @      @                                                                      @      @                       @      �?      @                               @             �q@     �T@     �m@      :@     @R@      =@      Q@     �f@     �t@     @P@     �O@     @_@     �v@     `s@      @     �G@      H@      X@      F@     �g@      4@     @^@       @      :@      *@      9@      a@      j@      0@      @@     �M@      l@      c@      �?      4@      0@     �H@      (@     �e@      4@     �V@      @      7@      &@      7@     ``@     �h@      ,@      ;@      K@     �i@      b@              4@      0@     �F@      (@     �V@      @     �C@      �?      @      @       @     �Q@     @]@      �?      "@      9@      \@     @P@              $@      @      1@      @     �N@      @      ;@              �?              @      8@     @T@              @      &@     @P@     �@@               @       @      $@      @      3@              @                                      (@      >@              @       @      0@      @              @              @       @      E@      @      7@              �?              @      (@     �I@              @      "@     �H@      :@              �?       @      @      �?      >@       @      (@      �?      @      @      �?      G@      B@      �?      @      ,@     �G@      @@               @      @      @      �?      5@      �?      "@      �?      @      @      �?     �D@      <@               @      @      D@      @@               @      @      @      �?      "@      �?      @                                      @       @      �?      �?      "@      @                                      �?             �T@      .@      J@      @      1@       @      .@     �N@      T@      *@      2@      =@      W@      T@              $@      "@      <@       @      ;@      @      $@       @      "@      @      @      >@     �A@       @      @      &@      7@      @@              @      @      "@       @      "@                       @      @              �?      ,@      &@              �?      @      $@       @                                              2@      @      $@              @      @       @      0@      8@       @      @      @      *@      8@              @      @      "@       @      L@      (@      E@      @       @      @      (@      ?@     �F@      &@      ,@      2@     @Q@      H@              @      @      3@      @      3@              $@      �?                      �?      ,@      *@      �?              "@      <@      3@              �?      �?      $@      �?     �B@      (@      @@      @       @      @      &@      1@      @@      $@      ,@      "@     �D@      =@              @      @      "@      @      ,@              >@      �?      @       @       @      @      (@       @      @      @      4@       @      �?                      @              &@              <@      �?               @       @      @      (@              @      @      4@      @      �?                      @               @              6@      �?               @       @       @      (@              @      @      $@      @                               @              @              1@                               @              @              @      @      @      �?                               @              @              @      �?               @               @      "@              �?      �?      @      @                                              @              @                                      @                              �?      $@       @      �?                       @              @               @                                                                              @       @                                                              @                                      @                              �?      @              �?                       @              @               @              @                                       @                              �?                                             �X@      O@     �]@      2@     �G@      0@     �E@      G@      ^@     �H@      ?@     �P@     �a@     �c@      @      ;@      @@     �G@      @@      P@      C@     @U@      .@      C@      *@      9@      3@     �P@     �A@      4@     �I@      U@     �\@      @      9@      ?@      B@      =@     �B@      ;@      H@       @      7@      @      0@      2@      I@      >@      (@      5@      J@      N@              5@      ,@      ;@      2@     �A@      ;@     �F@      @      4@      @      .@      1@      I@      1@      &@      .@      G@     �K@              2@      *@      7@      1@      "@      ,@      $@              @       @      @      @      3@       @      @      @      5@      (@               @       @      @       @      :@      *@     �A@      @      0@       @      "@      *@      ?@      .@       @      "@      9@     �E@              0@      &@      0@      "@       @              @       @      @      �?      �?      �?              *@      �?      @      @      @              @      �?      @      �?      �?               @                                                       @                      @      @                               @              �?              �?       @      @      �?      �?      �?              &@      �?      @       @       @              @      �?       @      �?      ;@      &@     �B@      @      .@       @      "@      �?      0@      @       @      >@      @@      K@      @      @      1@      "@      &@      "@      @      0@      @      @       @      @               @              �?      (@      3@      $@              @      *@              @               @       @      �?               @                      @                      &@              @              �?       @                      "@      @      ,@      @      @              @              @              �?      �?      3@      @              @      @              @      2@      @      5@       @       @      @      @      �?       @      @      @      2@      *@      F@      @              @      "@      @      &@      @      5@      �?      @      @      @      �?       @      @      @      2@      *@      E@      @              @       @      @      @      �?              �?      �?              �?                                                       @                              �?              A@      8@     �@@      @      "@      @      2@      ;@      K@      ,@      &@      .@      M@     �E@      @       @      �?      &@      @      *@      3@      *@      �?      @      @      @      0@      <@      *@      @       @      1@      "@              �?              @              @      ,@      &@      �?      @      @       @      *@      3@       @      @       @      ,@      @              �?              @              @       @      @              @               @       @      0@       @      @              @       @                              @              �?      (@      @      �?              @              @      @              �?       @      $@      �?              �?                               @      @       @              �?              @      @      "@      &@                      @      @                              �?               @               @                                      @      @      "@                       @      @                                                      @                      �?              @              @       @                      �?                                      �?              5@      @      4@       @      @              (@      &@      :@      �?      @      *@     �D@      A@      @      �?      �?      @      @      2@      @      ,@       @      @              &@      &@      8@      �?      @      $@     �D@      @@      @      �?      �?      @       @      0@      @      (@       @       @              @      @      8@      �?      @      $@      B@      8@      @      �?      �?      @               @               @              @              @      @                                      @       @                              �?       @      @              @                              �?               @                      @               @                                      �?      �?               @                                               @                                       @                                               @              @                              �?                                      @                                                      �?�t�bub��     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�5<{hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKqhnh4h7K ��h9��R�(KKq��hu�B�         6                    �?z�b�͓�?�	           ��@                          �4@N�°��?"           X�@                            �?H�����?�           �@       	                   �1@V����?z            @h@                          �0@=����?&            �K@������������������������       ��Cc}�?
             ,@                           �?���.}*�?            �D@������������������������       ���8��8�?
             (@������������������������       �x�-�?             =@
                          �3@iH?��?T            `a@                          �2@�F0b��?4            �T@������������������������       �������?            �G@������������������������       ����:���?            �A@                           �?M=ֱ߹�?             �L@������������������������       �@��Z��?             7@������������������������       �RC4%�?             A@                            @?O:!I
�?           |@                          �2@��$��3�?p             e@                           �?^}����?E             [@������������������������       ��f�l+��?            �C@������������������������       ��*��?+            @Q@                           �?� �Lˍ�?+            �N@������������������������       �����>4�?             <@������������������������       �Ȭ�@�S�?            �@@                          �0@����X�?�            �q@                           @ffffff�?             4@������������������������       �t�E]t�?             &@������������������������       ��2�tk~�?             "@                           �?s�O�+�?�            @p@������������������������       �l�Ӑ���?6            �U@������������������������       ����ѻ*�?i            �e@        -                   �?@�Ĩ��[�?�           L�@!       (                    �?��W�3�?X           8�@"       %                    �?�����?�            �t@#       $                    �?�J,jˈ�?<            �Z@������������������������       �\���(\�?             D@������������������������       ��n(T��?!            �P@&       '                    �?gz���?�            �l@������������������������       �      �?	             0@������������������������       �e��c��?�            �j@)       ,                   �>@��,~|E�?�           ��@*       +                    �?���7�?�           P�@������������������������       ����&�?�            �o@������������������������       ����zf�?�            �v@������������������������       �^N��)x�?	             ,@.       /                    �?�d�����?2             S@������������������������       ��m۶m��?	             ,@0       3                    @aS��/�?)             O@1       2                   �@@T�
�	�?             ?@������������������������       �.�袋.�?             6@������������������������       ���"e���?             "@4       5                    @l+�2���?             ?@������������������������       �      �?              @������������������������       �K����?             7@7       R                    @�D)QK��?�           f�@8       E                     �?]�=�R�?i           �@9       @                    @��W�M��?]           H�@:       =                    �?+m5ۂ�?�            @w@;       <                   �2@fl �&�?y             g@������������������������       �L�6�#��?%             O@������������������������       � ��i��?T            �^@>       ?                    �?������?�            �g@������������������������       ���LL=l�?3            @Q@������������������������       ������?R            �]@A       B                   �0@��i1�?_            �b@������������������������       �        
             (@C       D                     �?@Åar��?U             a@������������������������       ��zhr���?#            �L@������������������������       �     @�?2             T@F       K                    �?����a@�?           @{@G       J                   �9@G�6'�?h            �e@H       I                    �?�n���?Z            �a@������������������������       ��~3*�?1            �Q@������������������������       �����[�?)             R@������������������������       �8^s]e�?             =@L       O                   �6@2�,�F�?�            �p@M       N                   �1@A�@���?h            �e@������������������������       ��Wt����?#            �M@������������������������       ������?E            @\@P       Q                    @Ĭ뉳��?<             W@������������������������       �����X�?	             ,@������������������������       �|���?3            �S@S       b                    @fm�뙸�?+           ؓ@T       [                    @��d���?�           X�@U       X                   �1@��t���?�            �v@V       W                     �?0��b�/�?.            �R@������������������������       �T�r
^N�?	             ,@������������������������       �����N�?%            �N@Y       Z                   �2@&���^�?�             r@������������������������       �PV�}(h�?$             O@������������������������       �Y,�Z��?�            @l@\       _                     @��ճC��?�             v@]       ^                    �?SK�;	�?�             t@������������������������       �{���T�?U            �\@������������������������       ��(mA�t�?�            �i@`       a                    �?N贁N�?             >@������������������������       �
^N��)�?	             ,@������������������������       �      �?
             0@c       j                     @���|�?[           X�@d       g                   �3@\U��b�?           �z@e       f                   �1@Rh�W��?e             c@������������������������       ��ޚ����?'            �K@������������������������       �(F.[��?>            �X@h       i                     �?�;���?�             q@������������������������       �C��t���?}            @i@������������������������       �
�%����?,             R@k       n                   �6@     %�?M             `@l       m                   �5@S���Ą�?+            �R@������������������������       �hE#߼�?%             N@������������������������       ���X��?             ,@o       p                    �?�x�zrJ�?"             K@������������������������       �      �?             0@������������������������       ��F<�A+�?             C@�t�bh�h4h7K ��h9��R�(KKqKK��h��BC       0}@     @R@     pt@      @@      T@      =@      U@     ��@      �@     �L@     @V@      f@     ��@     @z@      ,@     �R@      J@      `@      F@      j@      :@     `d@      ,@     �F@      7@     �H@     �^@     �j@      ?@     �K@     @Y@     �n@     `i@       @      D@      B@     @R@      >@     �Y@       @     �H@       @      @              @     @V@     �Z@      @      3@      A@     @[@     @P@               @       @      @@      "@      ?@       @      ,@      �?                       @      7@      8@              "@      @     �H@      1@               @              $@      @      @              @                              �?      0@      @              @      �?      ,@      @                                      �?      @              @                                      @                                      �?       @                                               @              �?                              �?      (@      @              @      �?      *@       @                                      �?      �?              �?                                      @      �?                      �?      @       @                                              �?                                              �?      "@      @              @              $@                                              �?      9@       @      $@      �?                      �?      @      3@              @      @     �A@      *@               @              $@      @      1@       @      @      �?                              @      .@              @       @      *@      "@                              @       @      "@      �?      @                                      @      "@                      �?      $@      @                              @               @      �?              �?                              @      @              @      �?      @      @                              @       @       @              @                              �?      �?      @              @       @      6@      @               @              @       @      @                                                      �?       @              @       @      @                       @                               @              @                              �?               @                              .@      @                              @       @     �Q@             �A@      �?      @              @     �P@     �T@      @      $@      =@      N@      H@              @       @      6@      @      :@              (@              @              �?     �C@      C@      �?      @      &@      ,@      &@               @              @       @      0@              @               @              �?      9@      ?@              @       @      ,@      �?                                              @               @                                      ,@      @                       @      @      �?                                              "@              @               @              �?      &@      8@              @      @       @                                                      $@              @               @                      ,@      @      �?              @              $@               @              @       @      @               @               @                      @      @      �?                              @                                      �?      @              @                                      @       @                      @              @               @              @      �?     �F@              7@      �?                       @      ;@     �F@      @      @      2@      G@     �B@              @       @      1@       @      "@              �?                                      @                                       @      @                                              @                                                       @                                      �?      �?                                               @              �?                                      @                                      �?       @                                              B@              6@      �?                       @      6@     �F@      @      @      2@      F@      A@              @       @      1@       @      (@              @                                      @      3@       @       @      @      &@      *@              @      �?      @              8@              .@      �?                       @      .@      :@       @      @      *@     �@@      5@              �?      �?      (@       @     �Z@      8@     �\@      (@     �D@      7@      F@      A@     �Z@      :@      B@     �P@     �`@     @a@       @      @@      A@     �D@      5@     �Y@      8@     @[@      $@      ;@      6@      E@      A@     �Z@      7@      ?@     �K@     �`@     ``@      @      ;@      ;@     �C@      3@      D@      @      =@              "@      @      ,@      .@     �K@      @      0@      *@     �M@     �A@              @      @      2@      @      $@      @      @                              @      �?      ?@      �?      $@      @      ,@       @              @      �?       @      @      @      @      @                                      �?      *@              @              @      �?                               @      �?      @              @                              @              2@      �?      @      @      $@      @              @      �?              @      >@      @      6@              "@      @      "@      ,@      8@      @      @       @     �F@      ;@               @      @      0@      @      @              @                               @                       @                                                              @              :@      @      2@              "@      @      @      ,@      8@      @      @       @     �F@      ;@               @      @      (@      @     �O@      2@      T@      $@      2@      3@      <@      3@     �I@      1@      .@      E@      S@      X@      @      5@      7@      5@      (@     �O@      1@      T@      $@      0@      2@      :@      3@      G@      1@      .@      E@      S@      X@      @      4@      7@      5@      $@      C@      @      >@       @      @      @      &@      @      9@              �?      (@      K@     �A@               @      .@      @      @      9@      &@      I@       @      *@      ,@      .@      (@      5@      1@      ,@      >@      6@     �N@      @      2@       @      0@      @              �?                       @      �?       @              @                                                      �?                       @      @              @       @      ,@      �?       @              �?      @      @      (@              @      @      @      @       @       @      �?              �?              @                              �?                      @                              �?                               @              @       @       @      �?       @                      @      @       @              @      @      @      @       @       @       @               @       @      �?                                      �?      @       @              @      @      @               @               @              �?       @                                              �?      @                      @              @               @                              �?              �?                                                       @                      @      �?                                               @              @      �?       @                       @      �?      @                      �?              @               @                      �?                              �?                              �?                                              @                                      �?              @      �?      �?                       @              @                      �?               @               @     0p@     �G@     �d@      2@     �A@      @     �A@     �y@     �z@      :@      A@     �R@      v@      k@      @      A@      0@     �K@      ,@      \@      2@     �Q@      &@      2@      @      .@      a@     �f@      *@      1@     �C@     @d@     @]@      �?      (@      @      6@      @      P@      @     �D@       @       @      @      "@     �R@     �^@       @      "@      ,@     @Q@     @R@              @      �?      ,@       @     �J@       @      ;@      �?       @      @      @     @P@     �S@      @      @      &@     �F@     �L@              �?      �?      @       @      ?@              @              �?              @      E@     �I@       @      �?      @      0@      7@              �?              @              @                                                      <@      3@              �?       @      @      �?                              �?              9@              @              �?              @      ,@      @@       @               @      (@      6@              �?               @              6@       @      5@      �?      �?      @       @      7@      ;@      @      @      @      =@      A@                      �?      @       @       @              @      �?      �?               @      *@      &@      �?      @              &@      ,@                      �?               @      4@       @      ,@                      @              $@      0@      @       @      @      2@      4@                              @              &@      @      ,@      �?                      @      $@      F@      �?      @      @      8@      0@              @               @                                                                              (@                                                                                      &@      @      ,@      �?                      @      $@      @@      �?      @      @      8@      0@              @               @              @       @      @      �?                              @      ,@              @      @      @       @              @              �?              @      @      &@                              @      @      2@      �?                      2@       @              �?              @              H@      &@      =@      "@      0@      �?      @      O@      M@      @       @      9@     @W@      F@      �?      @       @       @      @      9@      $@      @      @      @      �?              5@      2@              @      ,@      D@      ,@              @              @       @      9@      $@      @       @       @      �?              3@      1@              @      "@     �A@       @              @              @       @      0@      @                      �?      �?              &@      (@                      @      *@      @                               @              "@      @      @       @      �?                       @      @              @      @      6@      @              @              �?       @                              @      �?                       @      �?                      @      @      @              @               @              7@      �?      9@      @      *@              @     �D@      D@      @      @      &@     �J@      >@      �?               @      @       @      0@              ,@      �?                      @      >@     �B@      �?      @      @     �C@      3@                       @       @              @              @                                      2@      ,@      �?                      @      "@                              �?              $@              &@      �?                      @      (@      7@              @      @      @@      $@                       @      �?              @      �?      &@       @      *@              @      &@      @      @       @      @      ,@      &@      �?                      �?       @                      �?       @                               @                              �?      @      @      �?                                      @      �?      $@              *@              @      "@      @      @       @      @      $@       @                              �?       @     `b@      =@     �W@      @      1@       @      4@     �p@     �n@      *@      1@      B@     �g@      Y@      @      6@      *@     �@@       @     �Q@      0@     �M@              @       @      @     @h@     �b@      @       @      1@     @Z@     �I@      �?      @      @      @      @     �B@       @      D@              @       @      @     �Q@     �S@      @      @      "@      L@      9@      �?      @      @      @       @      @                                              �?      A@      5@                      @      "@      �?                                              �?                                                      @       @                                                                                      @                                              �?      =@      *@                      @      "@      �?                                              ?@       @      D@              @       @       @     �B@      M@      @      @      @     �G@      8@      �?      @      @      @       @      &@              2@                                      .@      @                              "@      @                                              4@       @      6@              @       @       @      6@     �J@      @      @      @      C@      4@      �?      @      @      @       @      A@       @      3@              �?              @     �^@     �Q@      @       @       @     �H@      :@              �?      �?       @      �?      ;@      @      0@              �?               @     �]@      Q@      @       @      @      H@      5@              �?      �?       @      �?      @              @                              �?     �M@      :@               @      �?      ,@      @                                              7@      @      *@              �?              �?     �M@      E@      @              @      A@      0@              �?      �?       @      �?      @      @      @                              �?      @      @                       @      �?      @                                              @               @                                      �?      @                                      @                                              @      @      �?                              �?      @                               @      �?                                                      S@      *@     �A@      @      &@              ,@     @S@      X@      @      "@      3@     @U@     �H@      @      0@      @      :@      @      P@      $@      9@      @      @               @      O@     @T@      @       @      2@      L@      ?@              (@      @      6@      @      3@      @      @       @                      @      ?@      G@                      @      .@      $@              @      �?      @              *@                                                      "@      2@                      �?      $@      �?                              @              @      @      @       @                      @      6@      <@                      @      @      "@              @      �?       @             �F@      @      4@      @      @              @      ?@     �A@      @       @      (@     �D@      5@              @      @      1@      @      :@              ,@      @      @              @      8@      @@       @      @      (@      A@      .@              @      @       @      @      3@      @      @              @                      @      @       @       @              @      @               @              "@              (@      @      $@              @              @      .@      .@       @      �?      �?      =@      2@      @      @              @              @              @              @                      ,@      @      �?      �?              7@      $@              @              @              @              @                                      ,@      @      �?      �?              0@      @              @              @                                              @                                                              @      @                                              @      @      @              �?              @      �?      $@      �?              �?      @       @      @                      �?              �?      @      �?                                      �?      @      �?                      @                                      �?              @              @              �?              @              @                      �?      �?       @      @                                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�ahG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKqhnh4h7K ��h9��R�(KKq��hu�B�         8                    �?�V<�͔�?�	           ��@                           �?�=��*�?)           ��@                          �2@+�Y�T��?�           ��@       	                   �1@��M���?]            �_@                           @�Q�g���?1            @Q@                            �?��$�4��?'            �L@������������������������       �4�����?             ?@������������������������       ���?��?             :@������������������������       ���8��8�?
             (@
                           �?DO��O��?,            �L@                           �?��i��i�?             5@������������������������       �r�q��?	             (@������������������������       �0�����?             "@                            �?2�tk~X�?             B@������������������������       �����>4�?             @������������������������       �B�<x�u�?             =@                            �?q�K%���?'           p}@                           �?ӤJ���?W            �`@                           �?��WV��?&             J@������������������������       �      �?             0@������������������������       �X�<ݚ�?             B@                           �?WI)���?1            �T@������������������������       �6�h$��?	             .@������������������������       ���'s�	�?(             Q@                          �?@,�P&��?�             u@                            �?�8�4���?�            `t@������������������������       ��z&/��?]            �b@������������������������       �|�HH���?m             f@������������������������       �ffffff�?             $@       +                   �3@�q��/M�?�           @�@       &                    @)W����?�            @q@        #                    @ł�<��?�             k@!       "                     �?$Vn\1��?p             g@������������������������       ��g:b߱�?            �F@������������������������       �����?W            `a@$       %                    �?���'�?            �@@������������������������       ���ˠ�?             &@������������������������       ��9����?             6@'       *                   �2@���9�?%            �M@(       )                    @_�yܰ��?            �F@������������������������       �     ��?             @@������������������������       �ƵHPS!�?	             *@������������������������       �I�$I�$�?             ,@,       3                   �=@�W�~|�?�           ��@-       0                    �?t䮪^@�?�           x�@.       /                    �?,o���?�            �t@������������������������       �+�-UP��?N            �`@������������������������       �{s�"���?u             h@1       2                   �7@£��R`�?�            px@������������������������       ���N��P�?�            `k@������������������������       �FH��N��?v            �e@4       5                    �?� �H��?C            @[@������������������������       �������?
             .@6       7                   �@@*�6(���?9            �W@������������������������       ����.��?)            �P@������������������������       �����>�?             <@9       X                   �2@��|���?|           H�@:       I                     @���L�?�           H�@;       B                    �?a��zj�?R           p�@<       ?                     �?�"����?�            @k@=       >                    �?�A���?.            �R@������������������������       ������D�?            �C@������������������������       �|"����?            �A@@       A                   �0@����HY�?X             b@������������������������       ���*ʤ��?            �@@������������������������       �(�3
u�?E            �[@C       F                     �?a�y�3�?�            @u@D       E                   �0@rhˀ_��?�             m@������������������������       ���+	��?%            �P@������������������������       �OO@¶�?i            �d@G       H                   �0@�g:,v��?>            �Z@������������������������       �Zo��b�?             ?@������������������������       �����k�?.             S@J       Q                    �?I�!�9�?S            �^@K       N                   �1@�Ep�7�?             �H@L       M                    �?Dc}h��?             <@������������������������       �<ݚ)�?             2@������������������������       ��G�z��?             $@O       P                    @0�w¹��?             5@������������������������       �0�����?             @������������������������       �T�r
^N�?	             ,@R       U                    @�s��W#�?3            �R@S       T                   �0@*�)����?#            �H@������������������������       ���Q��?	             $@������������������������       �8��,�?            �C@V       W                    @`�Q��?             9@������������������������       ����S�r�?             ,@������������������������       �*L�9��?             &@Y       h                   �8@���VS�?�           �@Z       a                    @0�)���?�           t�@[       ^                   �5@�f��?�           0�@\       ]                    @� �=�e�?�           h�@������������������������       ��%)���?'            |@������������������������       ��fO�
�?q            `e@_       `                     @��76���?           �y@������������������������       ���(a�?�            u@������������������������       �z��z���?,            �S@b       e                    @6�ẗ��?<            @T@c       d                   �4@�GN��?0            �P@������������������������       �gE<j���?             =@������������������������       ��,b+���?            �B@f       g                    �?[�[��?             .@������������������������       �������?             @������������������������       �      �?              @i       p                   @A@^�DB,�?�            �y@j       m                    @9l��v�?�            �x@k       l                    @��J���?�            �u@������������������������       �Or;�}��?n             f@������������������������       �B��*$�?g            �d@n       o                   �<@r�q�?             H@������������������������       ������?             A@������������������������       �������?
             ,@������������������������       ��zv�X�?             6@�t�bh�h4h7K ��h9��R�(KKqKK��h��BC        {@     @S@     �t@     �F@     @P@      ?@      M@     h�@     P�@     �R@     �S@     `c@     p�@      z@      4@     �S@      P@     @_@     �N@     �h@      ?@     �d@      6@      E@      7@     �@@      a@      h@     �A@      N@     �R@     �n@     �j@      (@     �J@      I@     �P@     �F@     �Q@      "@      H@              $@       @      "@     �M@     �T@      "@      7@      B@     �[@     �N@              ,@      1@      5@      0@      2@      �?      @                              �?      :@      @@       @       @      &@      1@      @              �?              @      �?      "@              @                                      5@      ,@       @               @      $@      �?                              �?              @               @                                      5@      &@      �?              @      @      �?                                              @              �?                                      (@      "@                       @      �?                                                      �?              �?                                      "@       @      �?              @      @      �?                                               @              �?                                              @      �?              �?      @                                      �?              "@      �?      @                              �?      @      2@               @      @      @      @              �?              @      �?      @      �?      �?                                      @       @                               @       @              �?               @              @                                                       @       @                              �?      �?              �?              �?              @      �?      �?                                      �?                                      �?      �?                              �?               @               @                              �?       @      0@               @      @      @      �?                              �?      �?                       @                                      �?                              �?      @                                                       @                                              �?      �?      0@               @       @       @      �?                              �?      �?      J@       @      E@              $@       @       @     �@@     �I@      @      5@      9@     @W@     �L@              *@      1@      1@      .@      *@      @      *@              @               @      @      (@      �?      @      @     �D@      &@              @      @      @      @      @      �?      @                                       @      "@      �?       @      �?      *@      @              @      �?      @               @              �?                                              @                              @                              �?                      �?      �?       @                                       @       @      �?       @      �?       @      @              @              @              $@      @      $@              @               @      @      @               @       @      <@      @              �?       @      @      @                       @               @               @      �?      �?               @                      �?                      �?      @              $@      @       @              @                       @       @                       @      <@      @              �?      �?      �?      @     �C@      @      =@              @       @      @      <@     �C@      @      1@      6@      J@      G@              @      ,@      $@      &@     �B@      @      =@              �?       @      @      <@     �C@      @      0@      3@      J@      G@              @      ,@      $@      &@      5@      @      (@              �?              @      @      3@      @       @      @      3@      9@              @              @      @      0@      �?      1@                       @              6@      4@       @       @      (@     �@@      5@               @      ,@      @      @       @                              @                                              �?      @                                                             �_@      6@     �]@      6@      @@      5@      8@     @S@     @[@      :@     �B@     �C@      a@     @c@      (@     �C@     �@@     �F@      =@     �E@       @      7@      �?       @               @      G@     �B@      �?      @      @      J@      @@              @       @      &@      @      ?@       @      2@      �?       @               @      >@     �@@      �?      @      @     �E@      8@               @       @      &@      @      >@       @      0@      �?       @               @      <@      9@      �?      @      @     �@@      5@                               @      @      &@              �?                                      @      "@      �?       @              *@       @                                      @      3@       @      .@      �?       @               @      9@      0@              @      @      4@      3@                               @       @      �?               @                                       @       @                              $@      @               @       @      @              �?              �?                                       @      �?                              @                                                                      �?                                              @                              @      @               @       @      @              (@              @                                      0@      @                       @      "@       @               @                      �?      $@              @                                      .@      @                              @      @               @                      �?       @              �?                                      *@      @                               @      @                                               @              @                                       @                                      @                       @                      �?       @              �?                                      �?                               @      @      @                                              U@      4@      X@      5@      >@      5@      6@      ?@      R@      9@      >@      A@     @U@     �^@      (@     �A@      ?@      A@      7@     �R@      4@     @W@      .@      :@      *@      4@      ?@     �P@      0@      7@      @@     �T@     �[@      @      7@      7@      :@      1@     �C@       @      G@      @      (@      @      &@      (@      A@              @      $@     �I@     �F@      @      &@      1@      @       @      9@      @      5@      �?      @              @      @      @               @       @      8@      5@      @      �?              @       @      ,@      @      9@      @       @      @      @      @      ;@              @       @      ;@      8@              $@      1@              @     �A@      (@     �G@      &@      ,@      $@      "@      3@      @@      0@      1@      6@      @@     �P@       @      (@      @      4@      "@      9@      @      5@      @      @       @      @      *@      9@       @      "@      @      3@     �@@              @      @      1@      @      $@      @      :@      @      "@       @      @      @      @       @       @      0@      *@     �@@       @      @              @      @      $@              @      @      @       @       @              @      "@      @       @       @      &@      @      (@       @       @      @      @              �?      �?                                       @       @                                              �?      �?      �?              @               @      @      @       @       @              @      @      @       @       @      &@      @      &@      @      @      @       @               @      @      @       @      �?               @      @      @               @      &@               @      @      @      �?       @                                              �?               @      @      �?       @                      @      @      �?      @      @     �m@      G@     �d@      7@      7@       @      9@     Pz@     �|@     �C@      3@      T@     pu@     `i@       @      :@      ,@     �M@      0@      M@      @     �@@                              @     �l@     �d@      @      @      1@      X@     �D@              @      �?       @      @     �D@      @      1@                              @     @j@     `b@      @      @      (@      Q@     �A@              @      �?      @      �?      .@              @                              �?     �Y@      H@      �?      @       @      ;@      $@              �?              �?      �?      @              �?                                      ;@      5@              @      �?      *@      �?              �?                      �?      @              �?                                      1@      @              @               @                                                      �?                                                      $@      .@                      �?      @      �?              �?                      �?      $@              @                              �?      S@      ;@      �?              �?      ,@      "@                              �?              @              �?                                      6@      �?                              @                                                      @              @                              �?      K@      :@      �?              �?      "@      "@                              �?              :@      @      (@                              @     �Z@     �X@       @              $@     �D@      9@              @      �?      @              5@      @      @                              @      M@      R@       @              @     �A@      3@              @      �?      @              @                                                      3@      ?@                              @      @                                              ,@      @      @                              @     �C@     �D@       @              @      =@      0@              @      �?      @              @               @                                     �H@      ;@                      @      @      @                                                                                                      4@       @                              �?       @                                              @               @                                      =@      3@                      @      @      @                                              1@              0@                               @      5@      4@              �?      @      <@      @              �?               @      @      @              (@                               @      @      @              �?       @      1@                                                      @               @                                      @      @              �?       @      $@                                                                       @                                      �?      @                              $@                                                      @                                                       @      �?              �?       @                                                              �?              $@                               @      �?                                      @                                                      �?              �?                                                                              @                                                                      "@                               @      �?                                       @                                                      (@              @                                      1@      ,@                      @      &@      @              �?               @      @      $@               @                                      ,@      "@                       @      @      @                                              �?                                                      @       @                                       @                                              "@               @                                      "@      @                       @      @      @                                               @               @                                      @      @                      �?      @      �?              �?               @      @       @               @                                       @       @                                      �?              �?                      @                                                              �?      @                      �?      @                                       @             `f@     �D@     ``@      7@      7@       @      3@     �g@     0r@      B@      .@     �O@     �n@     @d@       @      4@      *@     �I@      &@     �c@      5@     �S@      0@      $@      @       @     �d@      m@      *@      (@      @@     `g@     �\@      @      ,@      @     �B@      @      b@      5@     �Q@      *@       @      @      @     �c@      l@      &@      &@      =@     �d@     �[@      @      (@      @      A@      @     @U@       @     �C@       @      @      @       @      \@      a@      @       @      .@     �Z@      K@              @      @      7@      @     �L@      @      ;@      @      �?      @      �?     �U@     �Z@      @      @      @     �T@     �@@              �?       @      4@      �?      <@      �?      (@      @      @              �?      9@      >@               @      "@      8@      5@              @      �?      @      @      N@      *@      @@      @      @              @     �G@     �U@       @      @      ,@     �L@     �L@      @      @       @      &@       @      J@      "@      >@      @       @              @     �@@     �R@       @      @      ,@      G@     �A@      @      @       @       @       @       @      @       @              �?                      ,@      (@                              &@      6@      �?                      @              (@              @      @       @              @      @      "@       @      �?      @      7@      @      �?       @              @              (@              @               @              �?      @      "@              �?      @      4@      @      �?                      @              @              �?                                      �?      @                              ,@      @                              �?               @              @               @              �?      @      @              �?      @      @              �?                       @                              �?      @                       @       @               @                      @                       @                                                                              �?                       @                       @                       @                                              �?      @                      �?       @                                      �?                                                      6@      4@     �J@      @      *@      @      &@      8@      M@      7@      @      ?@      N@      H@      @      @       @      ,@      @      5@      4@      E@      @      *@       @       @      8@     �L@      5@      @      ?@      N@     �G@      @      @       @      ,@      @      2@      2@     �B@      @       @       @      @      4@      K@      4@      @      ?@      L@     �C@      @      @       @      (@      @      (@       @      "@      @       @       @       @       @      4@      $@       @      1@      >@      =@      @      @       @      @      @      @      $@      <@       @                       @      (@      A@      $@      �?      ,@      :@      $@              �?      @      @              @       @      @              &@              @      @      @      �?                      @       @                               @      �?      @       @       @              @              @      @       @      �?                      @       @                                                              @              @                              �?                              �?                                       @      �?      �?              &@                      @      @              �?       @                              �?                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��LhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKehnh4h7K ��h9��R�(KKe��hu�B         2                    �?���(ل�?�	           ��@                            @������?�           d�@                           @{�]�e�?B           ؔ@                           @�9
i�&�?}            �@                          �2@h)�) �?g           ؁@                           �?�E����?W            �a@������������������������       �{�m<��?            �F@������������������������       ��*��G�?;            �W@	       
                   �8@�?�A`��?           �z@������������������������       �8	��W��?�             s@������������������������       ��s�� �?W            �_@������������������������       �"sLj�'�?            �D@                          �8@Hf�9w�?�           ��@                           @�d�g��?�            �@                          �1@FѬB�?Q            @a@������������������������       ���
I��?             ;@������������������������       ��`{g��?>            �[@                           @���u��?0           �}@������������������������       ��:�π��?           �{@������������������������       ��S�r
^�?             <@                           @0�3$v�?D            �[@                          �9@     ��?             @@������������������������       �������?	             *@������������������������       �窷uJ��?             3@                           @�7���?-            �S@������������������������       ������?             7@������������������������       �˕6�#��?             �K@       +                    @�@�N�m�?@           0~@       $                   �6@�o��u�?�            �v@       !                    �?�D��3��?�            `o@                           �2@�'ls��?I            �Z@������������������������       ����
�?            �B@������������������������       ���{��?.            �Q@"       #                    �?��^B{I�?]             b@������������������������       �R���Q�?             >@������������������������       ��|�i��?J            �\@%       (                    �?��*���?P            �\@&       '                    �?T�r
^N�?             <@������������������������       ��z�G��?	             $@������������������������       ��q�q�?             2@)       *                   �9@:El���??            �U@������������������������       ��R_�y�?            �F@������������������������       �7T�{�?             �D@,       1                    @gl��G��?J            �]@-       .                   �1@}������?B            �Z@������������������������       �j�V���?             &@/       0                    @
2���?<            �W@������������������������       ��5$``�?5            @T@������������������������       ���>4և�?             ,@������������������������       �r�q��?             (@3       H                    �?�v�x��?A           `�@4       ?                     @`�!�,��?�           ��@5       :                    @7V>��;�?           �z@6       9                   �9@�v��t�?�            @j@7       8                    �?h~�8�$�?p            �e@������������������������       �M�#:9�?L             ]@������������������������       ��Cc}�?$             L@������������������������       ��_�;���?             C@;       <                   �0@&�9�%�?�            �j@������������������������       �R���Q�?	             4@=       >                   �:@��<ʷ��?�            @h@������������������������       �*��r,�?t            �e@������������������������       �/�s��?             3@@       E                    @�B� ��?r            `e@A       D                   �=@�0��!��?d            @b@B       C                    �?���6c�?^             a@������������������������       ��"w����?             3@������������������������       �����W2�?N            @]@������������������������       �ffffff�?             $@F       G                   �7@p_�Q�?             9@������������������������       �l�l��?             .@������������������������       ��(\����?             $@I       X                   �7@c�4��?�           t�@J       Q                    @P��T�?Y           P�@K       N                    �?b0ݡ�?`           ��@L       M                     �?T�S�M�?�            �n@������������������������       �qX���?%             O@������������������������       �B��G�N�?k             g@O       P                   �2@4n`��?�            �s@������������������������       ��~VC�1�?O            �_@������������������������       ��q���?�             h@R       U                     @D��-s�?�            Pw@S       T                    �?�JfM�?�            �n@������������������������       �����P�?            �A@������������������������       ��QJ:H�?�             j@V       W                    @�M<�@��?S             `@������������������������       ����m�?J            �\@������������������������       ��h$���?	             .@Y       ^                    �?c�Y��?b           ��@Z       ]                   �=@��|���?             F@[       \                   �8@p��N�?             ?@������������������������       �"���c��?
             *@������������������������       �)O���?             2@������������������������       �pƵHP�?             *@_       b                   @@@!u�cA��?E           8�@`       a                     @+F�|��?$           @}@������������������������       �9��yo��?�            u@������������������������       �Ɩ��#��?S            ``@c       d                   �@@�a ߝ�?!            �I@������������������������       ��K8��?             *@������������������������       �kN¾�?             C@�t�bh�h4h7K ��h9��R�(KKeKK��h��B�;       `}@      T@     v@      B@     �R@      ;@      U@     (�@     ��@      N@      V@     `d@     ��@     �y@      @      J@     �K@     �\@      I@     �l@      5@     �_@      @      7@      @      >@     t@      w@      ,@     �D@     �O@     �r@     �e@              0@      .@      F@      7@     �f@      .@     @U@      @      .@              4@     pp@     `r@      "@      ?@     �C@     �i@     �]@              $@      @      <@      (@      Y@      *@     �H@      �?      $@              (@     @W@     �Z@       @      0@      5@     �V@      K@               @      @      4@      (@     �U@      *@      G@      �?       @              $@     �V@      Y@       @      $@      5@     �U@     �I@               @      @      4@      (@      <@       @      @                                      K@      <@                       @      1@      @                                              *@              @                                      "@      "@                       @      @       @                                              .@       @       @                                     �F@      3@                              &@      �?                                              M@      &@      D@      �?       @              $@     �B@      R@       @      $@      3@     �Q@      H@               @      @      4@      (@     �H@      @      ?@              @              @      >@     �L@      �?       @      0@      L@      ;@               @               @      @      "@      @      "@      �?      �?              @      @      .@      �?       @      @      ,@      5@              @      @      (@      "@      ,@              @               @               @       @      @              @              @      @                                              T@       @      B@       @      @               @     @e@     �g@      @      .@      2@     �\@     @P@               @      �?       @             @P@       @     �@@      �?                      @     �c@      f@      @       @      "@     �W@     �I@                      �?      @              5@      �?       @      �?                      @      9@     �L@      �?              @      *@      "@                                               @                                              �?      &@      (@                              �?                                                      3@      �?       @      �?                      @      ,@     �F@      �?              @      (@      "@                                              F@      �?      ?@                               @     �`@     �]@       @       @      @     @T@      E@                      �?      @             �@@      �?      ?@                               @     @_@      ]@       @       @      @      S@      E@                      �?      @              &@                                                      "@      @                              @                                                      .@              @      �?      @              �?      &@      (@      @      @      "@      5@      ,@               @              @              @                                                      @       @               @      @      @       @                              @               @                                                              @               @      @      �?                                                       @                                                      @      @                               @       @                              @              &@              @      �?      @              �?      @      @      @      @      @      2@      (@               @               @               @              �?              @                              �?              @      @      @       @               @                              "@               @      �?       @              �?      @      @      @      �?      @      *@      $@                               @             �I@      @     �D@       @       @      @      $@      M@     �R@      @      $@      8@      W@     �K@              @      "@      0@      &@      F@      @      >@       @      @      @      @      J@      J@      @       @      0@      O@      F@              @      @      "@      &@      @@      �?      0@       @      @      @       @      H@      ;@      �?      @      $@     �I@      A@              @              "@       @      2@      �?      @              @       @              &@      *@      �?               @      7@      3@               @               @      �?      &@      �?       @                                       @      @      �?               @      $@      �?              �?              @              @              �?              @       @              "@      $@                              *@      2@              �?              @      �?      ,@              *@       @              �?       @     �B@      ,@              @       @      <@      .@               @              �?      �?                      @                                      (@      @                      �?      @      @              �?                              ,@              $@       @              �?       @      9@      $@              @      @      6@      (@              �?              �?      �?      (@      @      ,@              @       @      @      @      9@       @       @      @      &@      $@              �?      @              "@      �?      �?      @                       @                      &@      �?      �?       @      �?      �?                                       @      �?      �?      �?                                              @      �?      �?      �?      �?                                                                      @                       @                       @                      �?              �?                                       @      &@      @      "@              @              @      @      ,@      �?      �?      @      $@      "@              �?      @              @       @      �?      @               @               @      @      "@      �?               @      @      @                      @              @      "@       @      @               @               @              @              �?       @      @       @              �?                      @      @      �?      &@              �?              @      @      6@       @       @       @      >@      &@              �?      @      @              @      �?      "@              �?              @      @      5@       @       @      @      8@      &@              �?      @      @              �?               @                                               @                                                                                      @      �?      @              �?              @      @      *@       @       @      @      8@      &@              �?      @      @              @      �?      @              �?              @      @      *@               @      @      2@      &@              �?      @      @                                                              �?      �?               @                      @                                      @              �?               @                                              �?                       @      @                                                     �m@     �M@     `l@      ?@      J@      6@      K@     �l@     �p@      G@     �G@      Y@     0s@     �m@      @      B@      D@     �Q@      ;@     �Q@      .@      H@      @      (@      "@      *@     �W@     �U@       @       @      8@     �R@     @S@              &@      "@      2@      "@      M@       @      ?@       @      @       @      &@     �U@     �L@       @      @      .@      F@      M@               @      @      .@      @      A@      @      6@       @      �?      �?      @      6@      7@      @      �?      $@      9@      B@               @       @      $@      @      ?@      @      4@                      �?      @      6@      4@      �?      �?      "@      5@      ;@               @       @      @      @      6@      @      *@                              �?      &@      &@      �?      �?      @      .@      3@              �?       @      @      @      "@              @                      �?       @      &@      "@                       @      @       @              �?                              @               @       @      �?              @              @      @              �?      @      "@                              @              8@      @      "@              @      �?      @      P@      A@      @      @      @      3@      6@              @      �?      @       @                                                              1@      @                                                                                      8@      @      "@              @      �?      @     �G@      ?@      @      @      @      3@      6@              @      �?      @       @      8@      �?       @              @              @      G@      ?@       @      @      @      3@      5@              @              �?      �?              @      �?                      �?              �?               @       @      �?              �?                      �?      @      �?      (@      @      1@      @      @      @       @      "@      >@               @      "@      ?@      3@              @      @      @       @      "@      @      1@      @      @      @      �?      "@      <@               @      @      8@      *@              @      @      @       @       @      @      0@      @      @       @      �?      "@      <@               @      @      8@      *@              @      @      @       @                                                              @       @              �?      �?      @      @               @      �?                       @      @      0@      @      @       @      �?      @      :@              �?      @      4@       @              �?      @      @       @      �?              �?              �?      @                                              �?                                      �?                      @      �?                      �?              �?               @                      @      @      @                      �?                      @                                                               @                              @      @                                                      �?                      �?              �?                                      @      @                              �?                      e@      F@     `f@      8@      D@      *@     �D@     �`@     �f@      C@     �C@      S@      m@      d@      @      9@      ?@     �J@      2@     @`@      5@      Z@      .@      *@      �?      2@     �[@      a@      *@      3@     �@@     �e@     �U@              .@      &@      <@      @     �X@      2@      K@       @      @              (@      Q@     �R@       @      $@      0@     @\@     �H@              @       @      *@      @      F@      @      ;@      @      @              @      *@      ;@      @      @      &@      H@      <@              @      @       @       @      @       @      @       @                      @      @       @      �?      @              3@      "@                               @             �B@      @      5@      @      @              @      @      9@      @      @      &@      =@      3@              @      @      @       @     �K@      &@      ;@       @       @              @     �K@     �G@      @      @      @     @P@      5@              @      @      @      �?      *@      @      @                              @      ?@      6@       @              �?      A@      @              �?       @      �?              E@      @      6@       @       @              @      8@      9@       @      @      @      ?@      1@               @      @      @      �?      ?@      @      I@      @       @      �?      @     �E@     �O@      @      "@      1@      O@      C@               @      @      .@      @      5@      �?      9@      @      @              @     �@@     �H@              @      *@      G@      3@               @       @       @      �?      �?                                              �?              $@                      @      1@      �?              �?                              4@      �?      9@      @      @              @     �@@     �C@              @      "@      =@      2@              @       @       @      �?      $@       @      9@      @      @      �?       @      $@      ,@      @      @      @      0@      3@                      �?      @      @      "@       @      9@      @      �?      �?       @      $@      "@      @      @      @      0@      ,@                      �?      @      @      �?                               @                              @                                      @                               @             �C@      7@     �R@      "@      ;@      (@      7@      6@      F@      9@      4@     �E@     �L@     @R@      @      $@      4@      9@      &@              �?      "@      �?              �?                      @       @                      @      *@      �?               @                              �?      "@      �?              �?                      @      �?                      @      "@                      �?                                      �?      �?                                       @                              �?       @                                                      �?       @                      �?                      @      �?                       @      �?                      �?                                                                                              @                              @      �?              �?                     �C@      6@     �P@       @      ;@      &@      7@      6@     �C@      1@      4@     �E@      K@      N@      @      $@      2@      9@      &@      B@      1@      N@      @      ;@      "@      7@      6@      B@      .@      2@      @@      J@      N@      @      $@      (@      6@       @      =@      *@     �C@      @      3@       @      *@      0@      =@      .@      &@      6@      F@     �@@              @      (@      1@      @      @      @      5@      @       @      �?      $@      @      @              @      $@       @      ;@      @      @              @      �?      @      @      @       @               @                      @       @       @      &@       @              �?              @      @      @      �?      @      �?      �?                                      �?      �?                                                      @       @               @       @      @      �?               @                       @      �?       @      &@       @              �?              @      �?      @�t�bub��     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�wthG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKehnh4h7K ��h9��R�(KKe��hu�B         0                    �?����&��?�	           ��@                          �5@P���?           H�@                           @Q:��s�?�           0�@                           �?!jo�#
�?�           ��@                          �1@�}R0)�?�            �u@                           @���R�?2            @T@������������������������       �ajgH��?#            �K@������������������������       ���1G���?             :@	       
                     �?����,E�?�            �p@������������������������       �^���� �?N            �^@������������������������       ���̼���?T             b@                           �?(���Pw�?�            �w@                            @W:��>�?Z            `a@������������������������       �^�T���?8            �T@������������������������       ���o+>�?"            �L@                            �?��.��?�             n@������������������������       �#e�����?/             R@������������������������       �r��n��?u             e@                            @�x���?             G@                           @�>4և��?             <@������������������������       ��
t�F��?             1@������������������������       �b���i��?             &@������������������������       ���"e���?	             2@       !                    �?������?           `�@                           �>@tXfgM��?�            �p@                           �?e��@���?�            �o@                            @a�ıI2�?B            �Y@������������������������       �4ܪ'z�?+            �O@������������������������       �>
ףp=�?             D@                          �7@/�s��?b             c@������������������������       ��c���+�?!             J@������������������������       ��~�:p��?A             Y@������������������������       ��m۶m��?             ,@"       )                    �?��R2��?f           ��@#       &                     �?r&����?Z            @a@$       %                   �8@90\�Uo�?             C@������������������������       �t�@�t�?             .@������������������������       �J��LQ�?             7@'       (                     �?�L�J��?A             Y@������������������������       ��V�D.(�?             =@������������������������       �B������?,            �Q@*       -                   �>@1�XC	��?           P{@+       ,                     @��3B5�?�            `w@������������������������       ���[ �Q�?�            �i@������������������������       �щ��sX�?`            �d@.       /                    @F��1{��?)            �O@������������������������       ������?            �@@������������������������       �� Ce���?             >@1       P                     @�R�J��?�           �@2       A                    @h���:��?�           ��@3       :                   �5@�D��m�?           �|@4       7                   �3@ �*����?�            �p@5       6                   �2@�-s|A�?m            `e@������������������������       ���L��"�?N            �^@������������������������       ��X����?            �H@8       9                    �?�~֌p��?8            �X@������������������������       �| /h�}�?            �C@������������������������       ����*�?&             N@;       >                     �?�W�>�?v            �g@<       =                     �?��w3��?]            @b@������������������������       �� ��V�?2            �S@������������������������       ��������?+             Q@?       @                    �?
x�¶�?            �E@������������������������       ���"e���?             "@������������������������       �� =[y�?             A@B       I                    �?ж'�l��?t           X�@C       F                     �?c�b�]�?0           @D       E                   �0@��1�8�?�            �t@������������������������       �     ��?             @@������������������������       �:%��`��?�            �r@G       H                    @Ew���-�?h            �d@������������������������       �٢��{�?M            �^@������������������������       ��3_<X�?             E@J       M                    �?TZk�?D           (�@K       L                   �>@; �P��?           �z@������������������������       ��Jn���?�            Py@������������������������       ��ˠT��?             6@N       O                   �3@����q�?=           �@������������������������       �;�4��`�?o            `f@������������������������       ���{����?�            pt@Q       Z                    �?�H���?           `y@R       Y                   �:@q5܀���?~            `g@S       V                    @!�K�[�?s            `e@T       U                    �?b3����?*            �P@������������������������       �"�����?             ?@������������������������       ������H�?             B@W       X                    @F��
ц�?I             Z@������������������������       ��l	H��?8            �S@������������������������       �xɃg\�?             :@������������������������       �     ��?             0@[       `                    @ه��V��?�            `k@\       ]                   �0@Ө*��?g            @c@������������������������       �     ��?             0@^       _                    @��t{H�?a            @a@������������������������       �R,K�H�?1            �R@������������������������       �     h�?0             P@a       b                   �3@��E)�?,            @P@������������������������       �     @�?
             0@c       d                    @�q��/��?"            �H@������������������������       �     p�?             @@������������������������       �|�l�]�?
             1@�t�bh�h4h7K ��h9��R�(KKeKK��h��B�;       0|@     @V@     �s@     �A@     �N@      ;@      V@     ��@     ��@      O@     @U@      c@     ȃ@      |@      "@     �K@     �J@      `@     �H@     @i@      F@     @d@      1@     �A@      6@     �G@     @^@     `f@      B@     �I@     �S@     �n@     �h@      @      @@     �@@     �P@     �C@     �`@      $@     �P@      @      @       @      "@      X@     �Y@      (@      0@      >@     `b@     �T@              "@      @      @@      (@      _@      $@      L@      @      @       @      "@     �W@     �X@      $@      .@      >@     �a@     @R@              "@      @      @@      $@     �Q@      @      .@                               @     �P@     �G@       @      @       @     �R@      =@              @              .@      @      6@              @                                      5@      2@                       @       @      @                                              0@               @                                      1@      @                       @       @      @                                              @              @                                      @      (@                                                                                      H@      @      "@                               @     �F@      =@       @      @      @     �P@      9@              @              .@      @      9@       @      @                              �?      7@      2@       @              @      B@      @               @              �?       @      7@       @      @                              �?      6@      &@              @      @      >@      4@              @              ,@      @      K@      @     �D@      @      @       @      @      <@      J@       @       @      6@     @Q@      F@              @      @      1@      @      4@      �?      (@                               @      &@      5@      @      @      &@      <@      (@              �?      �?       @      @      "@      �?      $@                              �?      $@      1@               @      "@      *@      @              �?              @       @      &@               @                              �?      �?      @      @      �?       @      .@       @                      �?      @       @      A@      @      =@      @      @       @      @      1@      ?@      @      @      &@     �D@      @@              @      @      "@      �?      @               @      �?                      @      @      &@       @      �?      �?      2@      .@                               @              ;@      @      5@       @      @       @       @      ,@      4@       @      @      $@      7@      1@              @      @      @      �?      &@              &@              �?                       @      @       @      �?              @      "@                                       @       @              @              �?                       @       @       @      �?              �?      @                                       @      @              @                                      �?       @       @      �?              �?      �?                                               @                              �?                      �?                                              @                                       @      @               @                                              �?                              @      @                                             �P@      A@     �W@      ,@      =@      4@      C@      9@     @S@      8@     �A@     �H@      Y@      ]@      @      7@      =@     �A@      ;@      :@      "@      @@              $@      @      @      *@      7@      @      "@      *@     �J@      ?@              @      *@      (@       @      :@      "@      =@              @      @      @      *@      7@       @      "@      (@      I@      ?@              @      *@      (@       @      $@      @      &@                       @       @      @      2@      �?      @      @      6@      "@                      @      �?      @       @       @      @                                      @      $@               @      �?      .@      "@                      @      �?               @      �?      @                       @       @      �?       @      �?      �?      @      @                              @              @      0@      @      2@              @      �?      @      @      @      �?      @       @      <@      6@              @      @      &@      @       @              (@                                       @      @               @              &@      @              �?              @      @       @      @      @              @      �?      @      @       @      �?      @       @      1@      3@              @      @      @      �?                      @              @                                      �?              �?      @                                                     �D@      9@     �O@      ,@      3@      1@      @@      (@      K@      5@      :@      B@     �G@     @U@      @      2@      0@      7@      3@      8@      @      .@      @      @      @      @       @      $@      @      @       @      2@      1@               @       @      $@      @      @              @      �?      �?              �?      �?       @      @                      @       @                               @               @              �?              �?              �?      �?       @      �?                      @      �?                                               @               @      �?                                               @                      �?      @                               @              4@      @      (@      @      @      @      @      �?       @      @      @       @      (@      "@               @       @       @      @      @       @      @              �?              @      �?      �?      @       @              �?      @                                              .@       @       @      @      @      @                      @               @       @      &@      @               @       @       @      @      1@      5@      H@      "@      ,@      ,@      ;@      $@      F@      ,@      6@      A@      =@      Q@      @      0@      ,@      *@      0@      ,@      4@      G@      @      &@      @      :@      $@     �D@      $@      4@      ;@      =@     �P@      �?      (@       @      $@      "@      $@      &@     �@@      @      @               @       @      2@      @      1@      $@      3@      ;@              (@      @       @      @      @      "@      *@       @      @      @      2@       @      7@      @      @      1@      $@     �C@      �?              @       @       @      @      �?       @       @      @      @      �?              @      @       @      @               @      @      @      @      @      @       @      �?      �?       @                                              @       @      @               @      @      @               @      @      �?              �?              @      @      �?              @      �?              �?                       @              @      �?      @      o@     �F@     �c@      2@      :@      @     �D@     �{@     �z@      :@      A@     @R@      x@     @o@       @      7@      4@      O@      $@     �i@      A@      `@      ,@      3@      @      <@     �w@     �w@      7@      =@     �O@     �s@     @f@      �?      2@      1@     �G@       @     �I@      @      @@       @      @      @      &@      L@     @]@      @      @      @     @T@     �I@              @      @      "@       @      @@              ,@      �?      �?               @      F@     @W@      �?      �?       @      D@      ;@              �?              @              3@              @              �?               @     �D@      N@      �?      �?       @      7@      (@              �?               @              ,@              @                               @      =@     �H@      �?      �?      �?      &@      "@              �?              �?              @              @              �?                      (@      &@                      �?      (@      @                              �?              *@               @      �?                      @      @     �@@                              1@      .@                              @              �?                                                              3@                              &@       @                                              (@               @      �?                      @      @      ,@                              @      @                              @              3@      @      2@      �?      @      @      @      (@      8@      @      @      @     �D@      8@              @      @      @       @      0@      @      (@      �?       @      �?      @      @      6@      @      @      @      7@      7@              @      @      @       @       @      @      @      �?       @              @      @      &@              @      @      1@      (@               @      @      �?       @      ,@       @      @                      �?              @      &@      @                      @      &@              @      �?      @              @      �?      @              @       @              @       @                      �?      2@      �?                                              @      �?                               @                                                      @                                                                      @              @                      @       @                      �?      .@      �?                                             `c@      <@     @X@      (@      (@      �?      1@     0t@     pp@      1@      6@      L@     �l@     �_@      �?      &@      *@      C@      @     �K@       @      8@               @      �?      �?     �a@     �[@      @      $@      ,@     �Q@     �F@              �?       @      @       @      9@              5@               @                     @X@      R@      @      @      &@     �K@      @@                       @      @      �?       @              �?                                      4@      @                              @                                                      7@              4@               @                     @S@     �P@      @      @      &@      J@      @@                       @      @      �?      >@       @      @                      �?      �?      G@      C@       @      @      @      .@      *@              �?                      �?      *@      @      �?                      �?      �?      E@      =@       @      @      @      *@       @                                              1@      �?       @                                      @      "@                               @      @              �?                      �?      Y@      4@     @R@      (@      $@              0@     �f@      c@      (@      (@      E@      d@     �T@      �?      $@      &@      A@      @      H@      @      8@      @      @               @     @[@     @U@       @      @      *@      P@     �A@               @      @      $@             �G@      @      3@      @      @               @     @[@     @U@      @      @      "@     �O@      ;@                      @      $@              �?              @                                                      �?              @      �?       @               @                              J@      1@     �H@      @      @               @     �Q@      Q@      @       @      =@     @X@     �G@      �?       @      @      8@      @      .@      @      @                              �?     �H@     �B@              �?      $@      B@      (@              �?      �?      @             �B@      (@      E@      @      @              @      6@      ?@      @      @      3@     �N@     �A@      �?      @      @      4@      @     �E@      &@      ;@      @      @      �?      *@      O@      H@      @      @      $@     �R@      R@      �?      @      @      .@       @      9@      @      (@      �?              �?      @     �B@      8@      �?       @      @      B@      6@              @       @      @      �?      9@              &@      �?              �?      @     �B@      6@      �?       @      @     �@@      6@                       @      @      �?       @              @      �?              �?              (@      "@                      @      5@      "@                                              @              �?                      �?              @      @                               @      @                                              �?               @      �?                              @      @                      @      *@      @                                              1@               @                              @      9@      *@      �?       @      �?      (@      *@                       @      @      �?      (@              @                                      6@      *@               @      �?      @      (@                              �?      �?      @              �?                              @      @              �?                      @      �?                       @      @                      @      �?                                               @                              @                      @               @              2@      @      .@      @      @              "@      9@      8@       @      @      @      C@      I@      �?      �?      �?       @      �?      ,@      @      &@      @       @              @      5@      ,@       @      @      @      <@      @@      �?      �?              @      �?                                                              "@                                              @                                              ,@      @      &@      @       @              @      (@      ,@       @      @      @      <@      9@      �?      �?              @      �?      (@      @      "@       @      �?              �?      @       @       @      @      @      ,@      $@      �?                       @               @      @       @      �?      �?               @      "@      @                      @      ,@      .@              �?              @      �?      @      �?      @              @              @      @      $@                              $@      2@                      �?       @                              �?                                       @      @                              �?      @                                              @      �?      @              @              @       @      @                              "@      (@                      �?       @              @      �?      �?               @              @       @      @                              "@      @                      �?       @              �?               @              @              @                                                       @                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJgo�MhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         >                   �5@N�"5u��?�	           ��@                           @� c7��?\           <�@                           �?)F�=�:�?�           ��@                           �?�+R�vg�?&           �|@                            @��v��?�            �s@                           @���Y��?s            `e@������������������������       ��P�[��?k            `c@������������������������       �      �?             0@	       
                   �4@�������?]            `b@������������������������       ��:��8{�?J            @]@������������������������       ���Q���?             >@                          �4@S��^�?V            �a@                            @�B�K/W�?H            @]@������������������������       ��2A]j�?1            @T@������������������������       ���a�2��?             B@������������������������       �$������?             9@                           �?Cy�5��?|            �@                           @fx+d\�?b            �c@                           �?��8���?=             X@������������������������       �L�.�3z�?#            �K@������������������������       �L�J��}�?            �D@                           @.����?%            �O@������������������������       ���ˠ�?             &@������������������������       ��q-�?             J@                          �4@�������?           |@                           @x����?�            v@������������������������       �����l�?�            `k@������������������������       � Qb$��?V            �`@                           �?�q��?;             X@������������������������       �YsW&�?)            �Q@������������������������       ���q���?             9@        /                    @강/���?�           ȑ@!       (                   �0@ѿ�Sr�?�           @�@"       %                     �?     `�?;             X@#       $                    @4և����?             E@������������������������       ��q�q�?             8@������������������������       ��������?             2@&       '                    @��Eac��?"             K@������������������������       �      �?             @@������������������������       ���#��Z�?             6@)       ,                    @�K�`�u�?�           @�@*       +                    @ٕ书��?           p|@������������������������       �֬�f��?	           �z@������������������������       �ݾ�z�<�?             :@-       .                     �?u�n\��?�             l@������������������������       ��ŏ1w�?@             Y@������������������������       �֑#����?J            @_@0       7                    �?�P/a���?�            �v@1       4                   �1@�{�q��?j            `f@2       3                     �?�ݒ�� �?             E@������������������������       ��e��a��?             9@������������������������       �J,�ѳ�?             1@5       6                    @|�I��?O             a@������������������������       �)C/Ap��?F            @^@������������������������       �     @�?	             0@8       ;                   �4@Ocq�21�?r            �f@9       :                    �?�Hx�5�?Y             b@������������������������       ��+\&p�?'             O@������������������������       ������?2            �T@<       =                     �?8��,�?            �C@������������������������       �^N��)x�?             ,@������������������������       ��D���J�?             9@?       Z                    �?b���/-�?9           ��@@       O                   �9@3���|�?�           8�@A       H                   �6@QL�K���?            z@B       E                    �?�b����?M            �^@C       D                     @�q�q��?              H@������������������������       �H�
R���?            �@@������������������������       ��X�%��?             .@F       G                    �?_�����?-            �R@������������������������       �^K�=��?             9@������������������������       �c�ZB>��?             I@I       L                    �?w��Qa�?�            pr@J       K                    �?�����?=            �X@������������������������       �������?             =@������������������������       �f ���?(            @Q@M       N                   �7@%�~��6�?|            �h@������������������������       �     ��?-             P@������������������������       �����?O            �`@P       W                   @@@�Xd�	�?�            Pp@Q       T                   �=@���kO��?�            �k@R       S                    @�� t���?t            �d@������������������������       �Ro�T���?I             [@������������������������       ��+�J��?+             M@U       V                     �?��e�S�?%            �L@������������������������       �������?             <@������������������������       �Ĝ�-�?             =@X       Y                    @�����?             C@������������������������       �<+	���?             .@������������������������       ��s-s��?             7@[       j                   �=@�O�]�k�?�           �@\       c                     @س��7�?&           x�@]       `                   �;@�;��K�?�            �@^       _                   �9@p�Im��?V           h�@������������������������       �P!�s���?           �x@������������������������       ��ز����?R            �_@a       b                    �?��Rw�$�?0            �T@������������������������       �Dy�5��?
             3@������������������������       �     ��?&             P@d       g                    @^ɏ���?�            �p@e       f                    @����&��?�            @l@������������������������       �j�]ث�?H            @^@������������������������       � �����?=            @Z@h       i                    @��`d�k�?            �F@������������������������       �     ��?             @@������������������������       ��1G����?             *@k       r                     @�|P�l�?a            �b@l       o                    �?1��N��?D            �Y@m       n                    �?w�J���?!            �I@������������������������       �]��N��?             3@������������������������       �      �?             @@p       q                   �@@g�M�4��?#            �I@������������������������       ��6c���?             A@������������������������       ��@�m�?             1@s       v                    �?B)�®�?            �G@t       u                   �@@�����?             ;@������������������������       ���&T���?             1@������������������������       ���Q��?             $@������������������������       �q=
ףp�?	             4@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       @{@      U@     0t@      :@     �Q@      :@      U@     ��@     `�@      R@      V@     `d@     ��@     p|@      *@     �R@     �H@     @_@     �N@     �q@      9@     `a@      @      4@      @      F@     {@     py@      4@     �A@     �R@     0x@      i@              <@      "@     �O@      :@      b@      ,@      T@      @      .@      @      =@      `@     @f@      ,@      5@     �F@      i@      \@              ,@      @      D@      3@      R@       @      =@               @       @      @     �R@     �T@       @       @      3@      Y@     �A@              @              0@      @      K@      �?      9@               @              @     �J@      F@      �?       @      *@     �P@      9@              @              "@      @      A@              (@              �?               @      A@      ;@              @      @     �A@      @              �?               @      @      8@              "@              �?               @      A@      ;@              @      @      A@      @              �?               @      @      $@              @                                                              �?              �?      �?                                              4@      �?      *@              �?              �?      3@      1@      �?      @      @      @@      2@              @              @       @      2@      �?      &@              �?              �?      2@      .@      �?      @      @      <@      $@              �?              @               @               @                                      �?       @                       @      @       @              @              @       @      2@      �?      @                       @              6@      C@      �?              @     �@@      $@                              @              1@                                       @              4@      @@      �?              @      7@      $@                              @              $@                                                      1@      5@                      @      *@      "@                              @              @                                       @              @      &@      �?              �?      $@      �?                                              �?      �?      @                                       @      @                      �?      $@                                                     @R@      (@     �I@      @      *@       @      :@      K@      X@      (@      *@      :@      Y@     @S@               @      @      8@      (@      8@      @       @                              @      (@      *@       @      @      &@      B@      1@               @      @      @       @       @      @      @                              @      $@      @              @      @      ?@      (@               @       @      �?              @       @      @                              @      @      @              @      @      (@      @              �?       @      �?              @      @       @                                      @       @                              3@      @              �?                              0@              @                              �?       @      @       @              @      @      @                      �?      @       @      @                                              �?                                       @      �?                              �?                      $@              @                                       @      @       @              @      @      @                              @       @     �H@      @     �E@      @      *@       @      4@      E@     �T@      @       @      .@      P@      N@              @      �?      1@      $@      D@      @     �C@      @      "@              @     �B@     �Q@              @      $@     �K@      G@              @              (@       @      2@      @      =@      @       @              @      <@     �A@              @       @      A@      ;@              �?              @      @      6@      �?      $@              �?                      "@      B@              �?       @      5@      3@              @              @      �?      "@      @      @              @       @      ,@      @      (@      @       @      @      "@      ,@              �?      �?      @       @      @       @       @              @       @       @       @       @      @       @      @      @      (@              �?      �?      @       @       @      �?       @                              @      @      @                              @       @                               @             `a@      &@     �M@       @      @              .@      s@     �l@      @      ,@      >@     `g@      V@              ,@      @      7@      @      T@      @      F@      �?      �?              @     �m@     `c@      @      &@      2@     �`@      N@               @       @      *@      @      &@              @              �?                      K@      0@                              @      @                               @              "@              @                                      .@       @                              @       @                               @              @                                                      &@      @                              �?                                                      @              @                                      @      �?                               @       @                               @               @                              �?                     �C@       @                               @       @                                               @                              �?                      8@       @                              �?       @                                                                                                      .@      @                              �?                                                     @Q@      @     �D@      �?                      @      g@     `a@      @      &@      2@      `@      L@               @       @      &@      @     �H@      @      @@      �?                      @      Z@     �T@      @      "@      0@     �X@     �C@               @       @      @      @      G@      @      ?@      �?                       @      X@     �T@      �?       @      0@     @V@     �C@               @       @      @      @      @              �?                               @       @               @      �?              "@                                                      4@      �?      "@                                      T@      L@      �?       @       @      ?@      1@                              @              (@               @                                      ;@      8@      �?       @              6@      $@                                               @      �?      @                                     �J@      @@                       @      "@      @                              @             �M@      @      .@      �?      @              &@     �P@     �R@       @      @      (@     �J@      <@              (@      @      $@       @      9@      �?       @              @              @     �D@      E@       @       @      @      ?@      "@               @              @               @              �?                                      3@       @                      @      @      �?                                              �?                                                      &@      @                      @      @                                                      �?              �?                                       @      @                              �?      �?                                              7@      �?      @              @              @      6@      A@       @       @      �?      8@       @               @              @              6@      �?      @              @                      4@     �@@       @       @      �?      2@       @               @               @              �?                                              @       @      �?                              @                                       @              A@      @      @      �?      �?              @      9@      @@              �?      @      6@      3@              $@      @      @       @      5@      @      @      �?      �?              @      3@      <@                      @      5@      *@              $@      @      @              1@      @      �?              �?              @      @      @                              "@      @              @       @      �?              @      @      @      �?                              *@      5@                      @      (@      @              @      �?      @              *@               @                              @      @      @              �?      �?      �?      @                                       @      @               @                              @      �?      �?                                      @                                              "@                                                      @      @              �?      �?      �?      @                                       @      c@     �M@      g@      3@     �I@      6@      D@     �Y@     �j@      J@     �J@      V@     �k@     �o@      *@      G@      D@      O@     �A@      P@      3@     @T@      @      (@      �?      ,@      I@      `@      @      2@      8@     �W@      X@              2@      2@      1@      *@      C@      @     �E@      @      @      �?      @     �B@     @W@      �?      $@      2@      N@     @Q@              @      (@      &@       @       @              *@      @      @              �?      *@      @@               @              ;@      0@                      @                      @              $@      @      �?              �?       @      @               @              ,@      �?                       @                      @              "@              �?              �?       @      @               @              "@      �?                                              �?              �?      @                                       @                              @                               @                      @              @               @                      &@      :@                              *@      .@                       @                      �?                                                      �?      &@                              @       @                                               @              @               @                      $@      .@                              "@      @                       @                      >@      @      >@                      �?      @      8@     �N@      �?       @      2@     �@@     �J@              @       @      &@       @      2@              @                              �?      @      <@              @      @      &@      (@              �?              @      �?      @              @                              �?              @              @      �?      �?       @              �?              @      �?      (@              @                                      @      7@                      @      $@      $@                                              (@      @      7@                      �?      @      1@     �@@      �?      @      *@      6@     �D@              @       @       @      �?      $@      �?      @                                       @      $@               @      @      "@      *@              �?              @      �?       @      @      4@                      �?      @      "@      7@      �?       @      $@      *@      <@               @       @      @              :@      ,@      C@      �?      "@              @      *@      B@      @       @      @      A@      ;@              ,@      @      @      &@      5@      ,@     �A@      �?      "@              @      *@      A@       @      @      @      @@      7@              @       @      @      "@      *@      *@      @@      �?      @              @      $@      :@      �?       @      @      6@      .@              @       @      @      @      @      @      :@               @               @      @      7@               @      @      @      &@              @      �?      @       @      @      @      @      �?      �?               @      @      @      �?                      0@      @              �?      �?              @       @      �?      @              @                      @       @      �?      @      �?      $@       @                               @       @       @      �?      @                                      �?      @      �?      @               @      @                               @      �?      @                              @                       @      @              �?      �?       @      �?                                      �?      @              @                              @               @      @       @      �?       @      @              @      @               @      @              �?                                                               @      �?                              @                              �?               @                              @               @      @                       @      @                      @               @      V@      D@     �Y@      ,@     �C@      5@      :@     �J@      U@      G@     �A@      P@     �_@     �c@      *@      <@      6@     �F@      6@     �T@     �A@     �U@      *@      ?@      *@      7@     �I@     �T@      <@      :@      H@     @^@     `a@      @      :@      $@      C@      2@      Q@      0@     @Q@      "@      2@       @      0@     �D@      J@      6@      1@      ;@     �W@     �T@      @      7@      "@      9@      &@      M@      *@      P@      @      2@       @      ,@     �D@     �D@      5@      *@      8@     �T@     �R@      @      4@      @      7@      @     �I@      "@     �F@      @      &@      �?      *@      <@     �B@      *@      &@      3@     �Q@      I@       @      ,@      @      ,@              @      @      3@              @      �?      �?      *@      @       @       @      @      (@      8@       @      @              "@      @      $@      @      @      @                       @              &@      �?      @      @      (@       @       @      @      @       @       @              �?                                       @               @              @              @                                              �?      $@       @      @      @                                      @      �?              @      "@       @       @      @      @       @      @      .@      3@      2@      @      *@      &@      @      $@      >@      @      "@      5@      :@     �L@      �?      @      �?      *@      @      $@      (@      2@      @       @      &@      @      "@      =@      @      "@      4@      (@      I@              @      �?      &@      @      "@      �?      @      @      @      @       @       @      7@      @      @      *@      $@      5@               @      �?      @      @      �?      &@      (@      �?      @      @      @      @      @      �?      @      @       @      =@              �?              @      @      @      @                      @              �?      �?      �?                      �?      ,@      @      �?                       @              @      @                       @                      �?      �?                      �?      &@      �?      �?                       @                                              @              �?                                              @      @                                              @      @      0@      �?       @       @      @       @       @      2@      "@      0@      @      4@      @       @      (@      @      @      @      @      ,@      �?       @      @      @              �?      "@      @      (@      @      .@               @      $@      @                       @      @      �?      @      @       @                      @      @      @               @               @       @      @                       @       @              @               @                              @       @                              �?       @                                      @      �?      �?      @                              @      �?      @               @              �?      @      @              @      �?      "@               @      �?      �?              �?      @              @      @      *@                       @      @                              @               @                              �?      @              @      @      "@                       @      �?              @      �?       @                      �?      �?                                       @              @                              @               @       @       @                      @               @      �?      "@      @      @              @      @               @              @      �?       @      �?                       @                      �?       @      @                       @      @               @              @      �?       @      �?                       @                      �?       @      @                       @                                       @                                                                                      �?                              @               @               @      �?              �?                      �?               @              @              @              @      �?                                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��|hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKqhnh4h7K ��h9��R�(KKq��hu�B�         8                   �2@�D�Xx��?�	           ��@                           @0y[ܨ��?�           ��@                           �?����[�?�           p�@                            @�k�{�?�            �s@                           �?�娈/H�?n            �f@                            �?�q�q�?,             R@������������������������       ���5�TB�?&             O@������������������������       �p=
ףp�?             $@	       
                    @��P��?B             [@������������������������       �U�6|���?              J@������������������������       �:/����?"             L@                          �1@HE$d�?K            �`@                           @8��,�?,            �S@������������������������       ���/5�?            �C@������������������������       ����З�?            �C@                           �?�Cc}h�?             L@������������������������       �     ��?	             0@������������������������       �q=
ףp�?             D@                           @��.b���?�            @u@                           @��;�L��?�            �l@                            @������?�            �i@������������������������       �1/�o���?N            @^@������������������������       �⎸#��?9            �U@������������������������       �'�%����?             7@                          �0@b)g���?@            �[@������������������������       �p�u=q��?             7@                           �?��ܞ��?5            �U@������������������������       �.��D�|�?            �A@������������������������       �O��N���?              J@       )                   �0@�7��ƻ�?            z@       $                    �?�X�C�??            �X@        !                    @2u�+���?$             M@������������������������       ��n���?             "@"       #                    @�|����?            �H@������������������������       �b+��c�?            �B@������������������������       ���8��8�?             (@%       &                    �?��Q���?             D@������������������������       ��q�q�?             (@'       (                     �? �Cc}�?             <@������������������������       ���X��?             ,@������������������������       �������?             ,@*       1                    @33333��?�             t@+       .                   �1@8�$�#��?�            �l@,       -                    �?2�tk~X�?E             [@������������������������       ����eP*�?             F@������������������������       �     (�?)             P@/       0                    @&}|�xI�?L            �^@������������������������       �R���Q�?             D@������������������������       ��^�X�=�?6            �T@2       5                    @l�����?;            @V@3       4                     �?<+	���?             >@������������������������       ��X�%��?	             .@������������������������       ��r����?             .@6       7                    @D[�F��?+            �M@������������������������       ���4��g�?            �A@������������������������       �UUUUUU�?             8@9       T                    �?��v���?	           2�@:       G                    �?��5��C�?U           �@;       @                     �?��!7r�?�            0x@<       ?                   �;@�A`��"�?:             Y@=       >                    �?2I�v���?3            �V@������������������������       �Few���?            �D@������������������������       �-�?���?            �H@������������������������       �333333�?             $@A       D                    �?P��`��?�            �q@B       C                     �?�;Z��?C            @Z@������������������������       ������j�?             H@������������������������       �z�J��?&            �L@E       F                    �?�\Z�Ny�?w            �f@������������������������       ��%`)���?<            �Z@������������������������       ���S����?;             S@H       M                    �?G�x�?a           ȍ@I       L                   �?@Й.���?�            �t@J       K                     �?�$���?�            �s@������������������������       �6y��D�?E            �Z@������������������������       ��C���?�             j@������������������������       ��θ�?             *@N       Q                   �>@�y,	�o�?�           ��@O       P                    �?
�i�?c           @�@������������������������       �Zy5� �?�            �i@������������������������       ��Ҕ!��?�            �u@R       S                    @�_|sܣ�?0            @R@������������������������       �     ��?             @@������������������������       ��O�`�I�?            �D@U       d                     @'4�Mp�?�           t�@V       ]                     �?	&��;�?�           ؒ@W       Z                    @�Na!�?           ��@X       Y                   �9@e�^����?<           �~@������������������������       �ဃ�][�?�            x@������������������������       ��є�!�?C            @Z@[       \                   �5@����k+�?�            pv@������������������������       �䙢�c�?n             g@������������������������       ��j U��?o            �e@^       a                    �? *4>HR�?�            Pv@_       `                    @�t����?`            `a@������������������������       �]����?E            @Y@������������������������       ��h�*$��?             C@b       c                   �5@���ފ��?�            @k@������������������������       ��A�e�?:            @W@������������������������       ��K�b��?K            @_@e       j                    �?���a��?�            pr@f       i                    @������?U            �_@g       h                    @Ç2�j��?N             ]@������������������������       ��ѳ�wY�?             A@������������������������       �h�T�B�?7            �T@������������������������       �ffffff�?             $@k       n                    �?��tG�?a             e@l       m                    @�q��/��?            �H@������������������������       ��ˠT�?	             6@������������������������       ���F�� �?             ;@o       p                   �5@贁N��?I             ^@������������������������       �$Vn\1��?             G@������������������������       �:��i~�?+            �R@�t�bh�h4h7K ��h9��R�(KKqKK��h��BC       �|@      U@     @u@      @@     �Q@      :@     �R@     H�@     ��@     �M@      \@      c@     ��@     �z@      3@     �O@     �J@     @`@      L@      _@      (@     �T@              @              "@     @q@     �k@      @      1@      8@     �g@     �O@              (@      @      ;@      @      V@      @     �K@              @              @     �\@     `a@      @      1@      3@      _@      G@              @      @      5@      @     �D@      @      0@                               @     @S@     @R@       @      @      @     �L@      4@              @               @              5@      @      @                                     �I@     �K@              @      @      8@      @                               @               @      �?      @                                      <@      .@              @              &@       @                                               @               @                                      <@       @              @              &@       @                                                      �?       @                                              @                                                                                      *@      @      @                                      7@      D@              �?      @      *@      @                               @              �?      @      @                                       @      7@                      �?      "@      @                                              (@                                                      .@      1@              �?      @      @      �?                               @              4@              "@                               @      :@      2@       @               @     �@@      *@              @              @              ,@              @                                      ,@      "@       @               @      7@      @                                              @                                                      $@       @      �?               @      1@       @                                              "@              @                                      @      @      �?                      @      @                                              @               @                               @      (@      "@                              $@      @              @              @              @                                                                                              �?      @              @              @              �?               @                               @      (@      "@                              "@       @                              @             �G@      @     �C@              @               @      C@     �P@       @      *@      (@     �P@      :@               @      @      *@      @      A@      @      7@              @              �?      @@      A@      �?       @      $@      H@      2@               @      @      "@      �?      >@      @      7@              @              �?      @@      @@      �?       @      $@     �B@      1@               @              @      �?      0@              &@              �?              �?      :@      *@      �?       @      "@      9@      @               @              @      �?      ,@      @      (@               @                      @      3@              @      �?      (@      $@                              �?              @                                                               @                              &@      �?                      @       @              *@              0@              �?              �?      @      @@      �?      @       @      3@       @                              @       @       @                              �?                              2@                               @                                                      &@              0@                              �?      @      ,@      �?      @       @      1@       @                              @       @       @              @                                               @      �?               @       @      @                              @              @              "@                              �?      @      @              @              .@      @                                       @      B@      @      ;@                              @      d@      U@                      @     @P@      1@              @              @              @              @                                     �M@      (@                      �?      &@      @                              �?              @              @                                     �A@       @                              @                                                       @                                                      @                                      @                                                      @              @                                      ?@       @                              @                                                                      @                                      :@      @                              @                                                      @                                                      @      @                              �?                                                       @              �?                                      8@      @                      �?      @      @                              �?                                                                       @      @                              �?                                                       @              �?                                      0@      �?                      �?      @      @                              �?               @                                                       @                              �?       @                                      �?                              �?                                       @      �?                              �?      @                                              =@      @      7@                              @     �Y@      R@                      @      K@      ,@              @              @              6@      @      1@                              @     @P@      L@                             �F@      &@              @               @              (@      �?      @                               @      ;@     �B@                              7@       @                              �?               @              �?                               @      0@      $@                              @                                                      @      �?       @                                      &@      ;@                              0@       @                              �?              $@      @      ,@                              @      C@      3@                              6@      "@              @              �?              @              *@                                       @      �?                              &@       @                                              @      @      �?                              @      >@      2@                              &@      @              @              �?              @              @                                     �B@      0@                      @      "@      @              @              @                              @                                      .@      @                      �?      �?                      @                                              @                                       @      @                      �?      �?                       @                                                                                      *@                                                               @                              @              �?                                      6@      (@                      @       @      @                              @              @              �?                                      0@      @                       @      @      @                                              @                                                      @      @                      �?      @                                      @             0u@      R@      p@      @@     �P@      :@     �P@     �n@     0w@     �K@     �W@      `@     |@     �v@      3@     �I@      I@     �Y@     �J@     �c@      B@     ``@      1@     �G@      4@     �A@     @P@      `@     �@@     �P@     �K@     `i@      e@      "@     �@@     �B@     �N@     �C@     �O@      "@     �A@      @      &@      @      @      2@     �L@      @      4@      *@      Q@     �G@       @      @      @       @      @      2@               @               @              @      @      2@       @      @      @      :@      @                       @      �?              (@              @               @              @      @      1@       @      @      @      :@      @                       @      �?              @               @                              @      �?      @              @       @      1@      �?                      �?                      @              @               @                       @      &@       @              @      "@      @                      �?      �?              @              �?                                              �?              �?                      �?                                             �F@      "@      ;@      @      "@      @      @      .@     �C@      @      0@      @      E@     �D@       @      @      @      @      @      "@       @      @               @                      "@      4@       @      *@      @      ,@      3@               @       @               @      �?       @      �?                                      @      &@              @      �?       @      (@                                      �?       @              @               @                      @      "@       @      @       @      @      @               @       @              �?      B@      @      5@      @      @      @      @      @      3@      �?      @      @      <@      6@       @       @       @      @      @      5@      @      .@               @                      @      ,@              @      �?      2@      0@       @       @              @      �?      .@      @      @      @      @      @      @      @      @      �?               @      $@      @                       @       @      @     �W@      ;@      X@      ,@      B@      ,@      =@     �G@     �Q@      <@      G@      E@     �`@     @^@      @      =@      ?@     �J@     �@@      F@      @      1@              1@      @       @      :@      :@      ,@      &@      ,@     �P@      :@              (@      @      2@      ,@      F@      @      1@              &@      @       @      :@      :@      ,@      "@      (@     �P@      :@              $@      @      1@      ,@      $@       @       @              @       @      @      @      @               @      @      <@      "@              @      @      @      $@      A@      @      "@               @      �?      @      7@      6@      ,@      @      @      C@      1@              @      @      $@      @                                      @                                               @       @                               @              �?              I@      6@     �S@      ,@      3@      &@      5@      5@     �F@      ,@     �A@      <@     @Q@     �W@      @      1@      8@     �A@      3@      H@      5@     �R@      "@      *@      @      2@      5@     �D@      &@      <@      :@     @Q@      W@      @      .@      1@      ?@      $@      5@      @      7@      @       @      �?       @      ,@      7@               @      $@      ?@      <@              @      *@      @       @      ;@      0@      J@      @      &@      @      $@      @      2@      &@      4@      0@      C@      P@      @      $@      @      <@       @       @      �?      @      @      @      @      @              @      @      @       @              @      @       @      @      @      "@       @      �?      @      �?                                       @      @      @                      @      �?       @              @      @                      �?      @      @      @      @               @              �?       @                      @              @      �?      @     �f@      B@     �_@      .@      4@      @      ?@     �f@     `n@      6@      =@     �R@     �n@      h@      $@      2@      *@      E@      ,@     @c@      6@     �Z@      @      ,@      @      1@     �b@     �j@      5@      9@     �J@     `i@      b@      @      .@      (@      A@      "@     �Z@       @     �R@      @       @       @      (@     �V@     �c@      0@      6@      C@      b@     �\@              $@      &@      7@      @      O@      @     �A@              @       @      "@      @@     �Z@      &@      &@      <@     �T@      S@              @      @      .@      �?     �E@       @      <@              �?      �?       @      :@      Y@      @      &@      8@     �N@      N@              @       @       @      �?      3@      @      @               @      �?      �?      @      @      @              @      5@      0@                      @      @             �F@      @      D@      @      @              @      M@      J@      @      &@      $@      O@      C@              @      @       @      @      >@              5@       @      @               @     �C@      <@       @      @      @      C@       @              �?                       @      .@      @      3@       @       @              �?      3@      8@      @      @      @      8@      >@              @      @       @      @     �G@      ,@      @@       @      @       @      @      M@      K@      @      @      .@     �M@      ?@      @      @      �?      &@      @      8@      @      &@       @      �?       @      @      =@      7@       @      �?      @      @      (@              @      �?      @      @      &@      @      "@      �?      �?       @      @      9@      4@              �?      @      @      "@              @      �?                      *@      �?       @      �?                              @      @       @                      �?      @               @              @      @      7@      @      5@              @               @      =@      ?@      @       @      (@      J@      3@      @                       @              1@       @       @               @                      3@      2@       @                      6@      @                              @              @      @      3@              @               @      $@      *@      �?       @      (@      >@      ,@      @                      @              <@      ,@      4@      "@      @       @      ,@      @@      >@      �?      @      5@     �E@      H@      @      @      �?       @      @      &@      �?      @               @      �?      @      9@      &@      �?      @      @      6@      8@               @      �?      @       @      $@      �?      @               @      �?              9@      &@      �?      @      @      6@      5@               @      �?      @       @      @              @                      �?              @      @                      @      @       @              �?                              @      �?       @               @                      3@       @      �?      @      �?      2@      *@              �?      �?      @       @      �?               @                              @                                                      @                                              1@      *@      *@      "@      @      �?      $@      @      3@                      0@      5@      8@      @      �?              @      @      $@       @              @                       @       @      $@                      @      @      @              �?              �?              "@      @               @                                      @                      �?               @                              �?              �?      @              �?                       @       @      @                      @      @      �?              �?                              @      @      *@      @      @      �?       @      @      "@                      $@      2@      5@      @                      @      @      @              "@      @       @              @       @      @                      @      "@      @                              �?              @      @      @      @       @      �?      @      @      @                      @      "@      2@      @                      @      @�t�bub��%     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ:��RhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKyhnh4h7K ��h9��R�(KKy��hu�Bx         >                    @�dU��?�	           ��@       !                   �4@_�Q.|��?�           ¡@                          �3@�紼�?$           x�@                           @ک'N��?�           p�@                           �?l{�%9`�?3           @@                            @S=��M�?�            @o@������������������������       �D� ʿ�?\            `c@������������������������       �<�-2W~�?0            �W@	       
                     @��U���?�            @o@������������������������       ��a�}��?]             b@������������������������       �Z������?J            @Z@                           @#(���?{            @g@                           �?uS�[�8�?W             `@������������������������       ���Coul�?            �B@������������������������       �����7��??             W@                          �1@Z��f��?$            �L@������������������������       �����K�?             2@������������������������       ��A�A�?            �C@                            �?���[�q�?v             h@                           �?P\>w��??            �[@                            �?zJ���?            �C@������������������������       �g\�5�?             :@������������������������       ��T�6|��?             *@                            �?�)O�?,             R@������������������������       �y�N����?            �@@������������������������       ���RT��?            �C@                           �?��� �?7            �T@                           @7��d��?             A@������������������������       ��q�q�?             8@������������������������       ���Q��?             $@                            @�����j�?             H@������������������������       �������?             2@������������������������       ��d��0�?             >@"       /                    �?1���=�?]           ȕ@#       *                     @������?�            x@$       '                   �;@}R�̈́�?�             o@%       &                   �8@�V�D.(�?�            `i@������������������������       ��^L���?`            �b@������������������������       �-����4�?&            �J@(       )                     �?��x�(�?!             G@������������������������       ��C��2(�?             &@������������������������       �p�_�Q�?            �A@+       .                   �=@�F����?S             a@,       -                    �?�q4;���?K            �]@������������������������       ��w�����?            �@@������������������������       �;"Z��?8            �U@������������������������       �4%���?             1@0       7                    �?��m~�?�?c           ��@1       4                    @������?�            pv@2       3                   �=@T9�vW��?m            �e@������������������������       ����:6�?]            �b@������������������������       ���c����?             :@5       6                    @Tmh����?s             g@������������������������       �u��,��?(            @P@������������������������       �v���� �?K             ^@8       ;                    @Z����l�?�           P�@9       :                   �=@���بD�?`            �e@������������������������       ��k���?R             b@������������������������       �/�����?             <@<       =                     @��|�<�?#           �}@������������������������       �.K�Bb�?�            �r@������������������������       �����o��?n            @f@?       \                   �2@�e�����?(           ��@@       O                    @} �==�?`           x�@A       H                    @���R�?           �z@B       E                     @��(�r�?�            �n@C       D                    �?�3e��k�?t            �d@������������������������       �@���4�?B            �V@������������������������       �^�(!�?2            @S@F       G                    @�p=
ף�?3             T@������������������������       �B���?             �H@������������������������       �w���<�?             ?@I       L                    @8@dO�%�?n            �f@J       K                    �?6 ��P��?            �A@������������������������       ��S����?	             3@������������������������       �      �?
             0@M       N                     @� �q��?[             b@������������������������       �!�nS�2�?U            �`@������������������������       �}��7�?             &@P       U                    @o�ŏ1�?K             Y@Q       T                     �?�J]�'G�?#            �G@R       S                   �0@     @�?             @@������������������������       ���Q��?             $@������������������������       ��!pc��?             6@������������������������       �0��b�/�?
             .@V       Y                    �?�M�84�?(            �J@W       X                   �1@+7����?             7@������������������������       �*L�9��?             &@������������������������       ��q�q�?             (@Z       [                   �1@�`�`�?             >@������������������������       �     ��?
             0@������������������������       �^N��)x�?             ,@]       l                   �8@~��g�?�           d�@^       e                     @%�$d��?'           Ȋ@_       b                    @я���?�           x�@`       a                    @s�I�Ж�?�           8�@������������������������       ��v�;�H�?           P|@������������������������       ��DaI7�?�            @h@c       d                    @����[�?)             R@������������������������       ��-؂-��?!             N@������������������������       ��������?             (@f       i                    @(�[�5�?Z            @a@g       h                    @�MJ��%�?4             U@������������������������       ��If%�9�?            �B@������������������������       � Q�"T��?            �G@j       k                   �4@}�����?&             K@������������������������       ��r
^N��?             <@������������������������       ����t���?             :@m       r                     �?    �+�?�             p@n       q                   �>@4ܪ'z�?,            �O@o       p                    @����X�?"            �H@������������������������       �333333�?             4@������������������������       ��کB���?             =@������������������������       �����X�?
             ,@s       v                     @�\^^�.�?u             h@t       u                    @LM�]�?[             c@������������������������       �L4S�u�?*            �P@������������������������       �
��r�c�?1            @U@w       x                    @�rcí�?            �D@������������������������       ����>4��?             ,@������������������������       ��L-���?             ;@�t�bh�h4h7K ��h9��R�(KKyKK��h��B�G       �{@     @V@     Pu@      =@     @T@      6@      W@     ��@     ��@     �R@     �U@     `c@     P�@     @}@      (@      P@     �F@     �]@      Q@     pp@      I@      m@      4@     �O@      6@     @P@     �g@     �r@      J@     �K@      [@     u@     `r@      @     �G@     �A@      T@     �J@     �`@      "@     �O@      �?       @              "@     �a@     `c@       @      (@     �@@     `d@     �U@              *@      @      5@      0@     �[@       @      J@      �?      @              @     �_@     @^@       @      (@      7@      ^@     �J@              $@      @      0@      $@     �U@       @      @@      �?      @              @     @[@      T@       @       @      0@     @U@      D@              @      �?      @       @     �G@       @      &@                              @     @R@     �E@       @      @      @     �A@      1@                              @       @      @@       @      $@                                     �H@      =@              @      @      *@      &@                              �?              .@              �?                              @      8@      ,@       @              @      6@      @                              @       @     �C@      @      5@      �?      @               @      B@     �B@              @      "@      I@      7@              @      �?      @      @      7@      �?      @      �?       @               @      8@      <@               @      @      8@      ,@              @               @      @      0@      @      ,@              @                      (@      "@               @      @      :@      "@               @      �?      �?              9@              4@              �?                      1@     �D@      @      @      @     �A@      *@              @       @      "@       @      &@              .@                                      ,@      A@      @              @      8@      "@                       @      "@       @       @              @                                              @      @              @      @      @                       @      @       @      "@              (@                                      ,@      =@                      �?      3@      @                              @              ,@              @              �?                      @      @       @      @       @      &@      @              @                              �?              @                                      @      �?      �?              �?      @                                                      *@              �?              �?                              @      �?      @      �?      @      @              @                              8@      �?      &@              �?              @      0@      A@                      $@     �E@      A@              @      �?      @      @      2@              @                               @      @      ;@                      @      5@      2@              @               @      @      �?                                              �?              &@                      @      0@      �?                                      @                                                      �?               @                              .@                                               @      �?                                                              @                      @      �?      �?                                      @      1@              @                              �?      @      0@                       @      @      1@              @               @              (@              @                                       @      �?                       @      @      @              �?               @              @                                              �?      @      .@                              �?      &@               @                              @      �?       @              �?               @      $@      @                      @      6@      0@                      �?      @               @              @              �?                      @      @                              @       @                               @               @                              �?                      @      @                              @      @                                                              @                                                                              �?       @                               @              @      �?      @                               @      @      @                      @      0@       @                      �?      �?              @      �?                                       @      @       @                       @              @                      �?      �?              �?              @                                               @                      @      0@      @                                              `@     �D@     @e@      3@     �K@      6@      L@      G@     �b@      F@     �E@     �R@     �e@     �i@      @      A@      ?@     �M@     �B@      E@      .@      D@      @       @      @      "@      *@     @R@      *@      ,@      6@      H@      G@      �?      @      @      (@      @      =@       @      7@      @      @      @      "@      @      K@      "@      $@      (@     �A@      8@      �?       @      @      "@      @      ;@      @      4@       @      @      @       @      @      F@      @      @      &@      A@      4@      �?       @      @      @      @      .@      @      0@               @       @       @      @      C@      @      @      "@      =@      (@               @      �?       @      @      (@      �?      @       @       @      �?                      @       @               @      @       @      �?               @      @               @      @      @      �?      �?              @      �?      $@      @      @      �?      �?      @                               @              �?              �?                                              @              �?      �?              �?                                              �?      @       @      �?      �?              @      �?      @      @      @              �?      @                               @              *@      @      1@       @      @      �?               @      3@      @      @      $@      *@      6@              @      @      @       @      (@      @      ,@       @      @      �?               @      3@      @              $@      "@      6@               @      �?      @       @      �?      �?       @                                      @       @      @              @              @              �?                              &@      @      (@       @      @      �?              @      &@                      @      "@      .@              �?      �?      @       @      �?              @                                                              @              @                      @       @                     �U@      :@     @`@      ,@     �G@      2@     �G@     �@@     �R@      ?@      =@     �J@     �_@      d@      @      ;@      9@     �G@      >@      C@      @     �B@      @      $@       @       @      0@     �@@      @      $@      *@     �P@     �P@              @      $@      $@      2@      2@      @      6@              @              @      (@      &@      @      @      @      4@     �C@              @       @      @      @      (@       @      6@              @              @      &@      &@      �?      @      @      3@      B@              @       @      @       @      @      �?                                              �?               @       @      �?      �?      @               @              @      @      4@      @      .@      @      @       @      @      @      6@              @      @      G@      <@              �?       @      @      (@      @       @      @      @      @              @      �?      $@              @       @      &@      @                                      @      .@      �?       @      @      �?       @      �?      @      (@               @      @     �A@      5@              �?       @      @      @      H@      4@     @W@       @     �B@      0@     �C@      1@      E@      <@      3@      D@      N@     �W@      @      5@      .@     �B@      (@      @      @      .@              "@      @      "@      @      3@      .@              @      5@      7@      �?      @      @      3@      �?      @      @      .@              "@      �?      "@      @      2@      @              @      4@      2@              @      @      3@      �?                                              @                      �?      &@               @      �?      @      �?      @                              F@      *@     �S@       @      <@      &@      >@      $@      7@      *@      3@     �@@     �C@     �Q@      @      .@      $@      2@      &@      =@      @      G@      @      6@      @      1@      "@      ,@      &@      *@      8@      >@     �@@              (@      @      (@      @      .@      @      @@       @      @      @      *@      �?      "@       @      @      "@      "@      C@      @      @      @      @       @     �f@     �C@      [@      "@      2@              ;@      v@     Pr@      7@      ?@     �G@      o@     �e@      @      1@      $@      C@      .@      G@      @      A@              �?              @     �g@      [@      @      �?       @     �S@     �B@              @              @              >@      @      @@              �?              @     �e@     �U@       @      �?      @      N@      9@                                              5@      @      <@              �?              @      V@     �D@       @      �?      @      D@      ,@                                              &@      @      @                              @      Q@      9@       @      �?       @      @@      &@                                              @      �?      �?                              @     �C@      4@                       @      0@      @                                              @      @      @                              �?      =@      @       @      �?              0@       @                                              $@              5@              �?                      4@      0@                      �?       @      @                                              @              4@                                      @      "@                      �?      @      �?                                              @              �?              �?                      .@      @                              �?       @                                              "@              @                              �?     @U@      G@                      @      4@      &@                                              @                                                      8@       @                              @                                                                                                              0@                                      @                                                      @                                                       @       @                               @                                                      @              @                              �?     �N@      F@                      @      .@      &@                                              @              @                                      N@     �C@                      �?      .@      &@                                              �?                                              �?      �?      @                      @                                                              0@       @       @                              �?      1@      5@       @              �?      2@      (@              @              @               @      �?                                      �?      $@       @                               @      $@                              �?              @      �?                                      �?      @      @                              @      @                              �?               @                                                      @       @                              �?                                                      @      �?                                      �?       @      @                              @      @                              �?              �?                                                      @      �?                              @      @                                               @      �?       @                                      @      *@       @              �?      $@       @              @              @              @      �?      �?                                      @       @       @                      @      �?                                              @                                                       @      @                              @                                                              �?      �?                                      �?      @       @                      �?      �?                                              @              �?                                      @      @                      �?      @      �?              @              @              @              �?                                               @                              @                      �?              �?                                                                      @      @                      �?              �?               @              @             �`@     �@@     �R@      "@      1@              5@     �d@      g@      3@      >@     �C@     `e@      a@      @      ,@      $@     �@@      .@      \@      0@     �H@      "@      @              .@      c@     �d@      "@      5@      7@     �`@     �X@      @      $@      @      7@      @      X@      ,@     �E@      @      @              &@     �`@     `b@       @      ,@      3@     �[@     �Q@      �?      $@      @      3@      @     @V@      ,@      A@      @      @              $@      ^@     `a@      @      "@      1@     �W@     �Q@      �?      $@      @      1@      @     �Q@      @      ;@       @      �?              @     �V@     �W@      @      @      &@      Q@      J@              @              @      @      3@      @      @       @      @              @      >@     �F@       @      @      @      :@      2@      �?      @      @      &@      �?      @              "@      �?                      �?      .@       @       @      @       @      1@      �?                       @       @              @               @                              �?      (@       @              @       @      .@                                       @                              �?      �?                              @               @                       @      �?                       @                      0@       @      @      @                      @      2@      1@      �?      @      @      6@      ;@      @                      @       @      &@       @       @       @                       @      (@      .@      �?      �?      �?      ,@      3@                                       @      @              �?       @                               @      @                              @      $@                                       @      @       @      �?                               @      @      (@      �?      �?      �?      @      "@                                              @              @       @                       @      @       @              @      @       @       @      @                      @              @              @       @                              �?      �?              @      @      �?      @                              @               @              �?                               @      @      �?                              @      @      @                      �?              7@      1@      9@              (@              @      &@      5@      $@      "@      0@      C@     �C@       @      @      @      $@       @      "@      �?      @              �?               @      @      @      �?              @      @      2@                      @      @              @      �?      @                              �?      @      @      �?              �?      @      2@                      @      @              �?      �?       @                                      @      @                                      @                       @      @              @              �?                              �?      �?              �?              �?      @      ,@                      �?                      @              @              �?              �?              �?                       @                                               @              ,@      0@      2@              &@              @      @      1@      "@      "@      *@      A@      5@       @      @       @      @       @      $@       @      0@              &@              �?      @      0@      "@      "@      (@      8@      2@       @      �?               @      @      @               @              &@                      @      "@      @       @      @       @      $@       @      �?              �?              @       @      ,@                              �?       @      @      @      @       @      0@       @                              �?      @      @       @       @                              @              �?                      �?      $@      @              @       @      @      �?      @      @                                                                                      @                      �?                      �?              @       @                              @              �?                      �?      @      @               @       @      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�a2hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         <                    �?u`��?�	           ��@       !                    @��?� ��?t            �@                          �2@.?�跙�?V           ��@                          �1@���%q��?�            �l@                            �?��d�&4�?O            ``@                           �?<��KM��?.             S@������������������������       ��ˠT�?             6@������������������������       �Һ��Ea�?              K@	       
                   �0@,��Y��?!            �K@������������������������       ����>4��?             ,@������������������������       ��E��{�?            �D@                           @��7���?B            @X@                           �?�9��%��?+            �O@������������������������       �~X�<��?             ;@������������������������       �������?             B@                            @%����?             A@������������������������       ����,�?             3@������������������������       ��������?	             .@                           �?Y�4=��?�           h�@                           @�X�wN�?}            @h@                          �3@U����1�?N             ]@������������������������       ��ˠT�?             &@������������������������       �'Cta���?F            @Z@                          �9@�.y0���?/            �S@������������������������       �2�PZi�?!            �J@������������������������       ���~j�t�?             9@                          �5@��&1��?H           X�@                            �?������?s            @f@������������������������       ����w��?:            @V@������������������������       �
�g����?9            @V@                           �9@g.I�/�?�            �u@������������������������       ��D��?|            �h@������������������������       �K?�'|��?Y            �b@"       1                    @򝿉�n�?           ��@#       *                   �2@ʁ쯷��?s           0�@$       '                    @�qv�F��?�            p@%       &                   �0@@�bY�p�?Z            �b@������������������������       ��������?             4@������������������������       �     !�?L             `@(       )                    �?ĘT���??            @[@������������������������       �l�L���?              M@������������������������       �� =[y�?            �I@+       .                    @���J7�?�            Pt@,       -                    @~�5τ��?~            �g@������������������������       �g�6���?G            @[@������������������������       �.��#VL�?7            �S@/       0                   �8@������?\             a@������������������������       �B���%%�?N            �\@������������������������       ��T�x?r�?             6@2       7                     @�6�����?�            q@3       6                    @5yy8,�?�             k@4       5                   �5@\��"e��?{            �h@������������������������       �>���L�?N            �`@������������������������       �����r�?-            @P@������������������������       �P7�Z�?             3@8       ;                   �8@�m۶m��?#             L@9       :                   �3@�J�կ�?            �E@������������������������       ����^B{�?             2@������������������������       ��
F%u�?             9@������������������������       ��q-��?             *@=       Z                     @�'�n�?9           ��@>       K                    �?5�s��?�           0�@?       F                   �>@q_�[9�?O           ��@@       C                    �?:m����?5            ~@A       B                   �9@�jA��?T            �`@������������������������       ����C&�?A            �X@������������������������       �%����?             A@D       E                    @,
l���?�            �u@������������������������       �"mdk���?�             u@������������������������       �}��7�?             &@G       H                    @     ��?             H@������������������������       �333333�?             4@I       J                     �?���S�r�?             <@������������������������       �����W�?             *@������������������������       ��A��S�?             .@L       S                   �5@0�� �w�?S           ��@M       P                    @^�?8�~�?R           H�@N       O                     �?�S�����?K            �^@������������������������       �a��"A�??             Z@������������������������       �R�n��?             2@Q       R                    �?���c�e�?           �z@������������������������       ���/����?Z            �a@������������������������       �O��e�?�             r@T       W                    @�[O�)�?           0y@U       V                    @�E�)��?�            0r@������������������������       ��2WW���?�            `n@������������������������       �UUUUUU�?             H@X       Y                    @�)x9o�?C             \@������������������������       �nqwZ���?<            @X@������������������������       ���A���?             .@[       j                    @R�ԛ@�?�           ��@\       c                    @�
�1�?�            �w@]       `                    @_fȪ G�?�            0t@^       _                    @H�V�:V�?�            @r@������������������������       ��镲q�?�             i@������������������������       �C%��N��?<             W@a       b                   �1@������?             ?@������������������������       ��h$���?
             .@������������������������       �     ��?             0@d       g                   �2@�X�C�?%             L@e       f                    �?�ˠT��?             6@������������������������       �      �?             (@������������������������       ��������?             $@h       i                   �5@%����?             A@������������������������       �0��b�/�?	             .@������������������������       �P7�Z�?             3@k       r                   �4@"�Q*�	�?�            @o@l       o                   �2@7mD<+�?J            �_@m       n                    @����^D�?'            �O@������������������������       �A�@���?            �E@������������������������       ��������?             4@p       q                    @      �?#             P@������������������������       �� =[y�?
             1@������������������������       �ހ���?            �G@s       v                   �=@3�a���?Q            �^@t       u                    @�$I�$��?J             \@������������������������       ���	A��?6            �R@������������������������       ��,�El�?            �B@������������������������       ��T�x?r�?             &@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       Pz@     @S@     Pu@     �A@      Q@     �@@     @V@     x�@     ��@     @Q@     �U@     @f@     @�@     `x@      1@     @Q@      M@     @^@     �N@     @h@      F@     @b@       @      1@      @      <@     �u@      u@      6@      <@     �I@     `s@      c@       @      =@      2@     �B@      7@     �[@      9@     @X@       @      ,@      @      5@     �\@     @c@      &@      3@     �B@      c@     �V@       @      8@      1@      6@      5@      9@       @      "@                                     �P@     �O@      @      �?      @      @@      ,@               @              @              &@              @                                      G@     �C@      @      �?      �?      3@       @                               @               @              �?                                      B@      6@              �?      �?      "@       @                               @                              �?                                      @      @                      �?      @       @                                               @                                                      >@      .@              �?              @                                       @              "@              @                                      $@      1@      @                      $@                                                      �?              @                                      @       @                               @                                                       @              �?                                      @      .@      @                       @                                                      ,@       @      @                                      4@      8@                      @      *@      (@               @              @              @       @       @                                      (@      5@                               @      "@              �?               @              @      �?                                              @      @                              @      @              �?               @              �?      �?       @                                      @      .@                              @      @                                               @              �?                                       @      @                      @      @      @              �?               @              @              �?                                      @       @                      @       @      �?                                              �?                                                      @      �?                              @       @              �?               @             �U@      7@      V@       @      ,@      @      5@     �H@     �V@      @      2@     �@@      ^@      S@       @      6@      1@      0@      5@      4@      @      1@               @       @      @      0@      >@      @      @      "@      F@      0@              @              @      @      "@       @      1@                              @      @      6@      @      @      @      6@      $@              @              @      @                       @                                       @      �?                       @              @                                              "@       @      .@                              @      @      5@      @      @      @      6@      @              @              @      @      &@      �?                       @       @       @      "@       @      @      @      @      6@      @              @               @              $@      �?                      �?       @              @       @      @      @      @      @      @              @              �?              �?                              �?               @      @                                      .@       @                              �?             �P@      4@     �Q@       @      (@      @      0@     �@@     �N@              (@      8@      S@      N@       @      .@      1@      &@      0@      <@              1@              @       @       @      5@      >@              @      @     �@@      7@               @              @      @      0@               @              �?               @      *@      0@               @      @      1@      @               @              @              (@              "@               @       @               @      ,@              �?      @      0@      2@                              �?      @      C@      4@      K@       @      "@      �?      ,@      (@      ?@              "@      1@     �E@     �B@       @      *@      1@      @      *@      5@      @      A@      @      @      �?      &@      &@      5@              @      *@      2@      9@      �?       @       @       @              1@      *@      4@      @      @              @      �?      $@               @      @      9@      (@      �?      @      "@      @      *@     �T@      3@     �H@              @              @     @m@     �f@      &@      "@      ,@     �c@     �O@              @      �?      .@       @      J@      "@     �B@              @              @      g@     �\@       @      @      @     �Z@     �A@              @      �?      "@      �?      5@      @      (@                              @     @]@      N@                              ?@      $@                                              .@      @      &@                              @      L@     �B@                              0@      @                                              �?                                                      *@      @                               @                                                      ,@      @      &@                              @     �E@     �@@                              ,@      @                                              @              �?                                     �N@      7@                              .@      @                                              �?              �?                                      F@      @                              @                                                      @                                                      1@      1@                              "@      @                                              ?@      @      9@              @               @     �P@     �K@       @      @      @      S@      9@              @      �?      "@      �?      .@      @      1@               @               @      ;@      =@       @      @      @      G@      .@              �?      �?      "@              *@      @      @                               @      *@      6@      @       @      �?      9@      "@                               @               @       @      (@               @                      ,@      @       @      @      @      5@      @              �?      �?      �?              0@      �?       @              �?                      D@      :@              �?      �?      >@      $@               @                      �?      &@               @                                      C@      8@              �?      �?      8@      @                                      �?      @      �?                      �?                       @       @                              @      @               @                              ?@      $@      (@                               @      I@     �P@      @       @       @     �I@      <@               @              @      �?      <@      @      &@                                      E@     �O@      �?       @      @      C@      5@              �?                      �?      9@      @      &@                                     �C@      O@      �?       @      @      ?@      4@                                              2@      �?      "@                                      @@      F@      �?              �?      4@      @                                              @       @       @                                      @      2@               @      @      &@      *@                                              @                                                      @      �?                       @      @      �?              �?                      �?      @      @      �?                               @       @      @       @               @      *@      @              �?              @              �?              �?                               @      @      @       @               @      *@      @              �?              @                                                               @      @       @                       @      @      �?              �?                              �?              �?                                      @      �?       @                      @      @                              @               @      @                                              �?      �?                                                                       @             `l@     �@@     `h@      ;@     �I@      <@     �N@     @j@      r@     �G@     �M@     �_@      s@     �m@      .@      D@      D@      U@      C@     �c@      ,@     `a@      .@      ;@      0@     �A@      g@      j@     �@@     �E@     @U@      m@     @b@      @      ;@     �@@     @P@      4@      G@       @     �O@      @      ,@      $@      4@      C@      I@       @      ;@     �C@     @T@      M@      �?      (@      .@      9@      ,@      G@       @     �M@      @      &@      @      3@      C@      H@      @      8@      7@     @T@      M@      �?      &@      "@      8@      (@      7@              "@               @              @      &@      3@              @      @      .@      2@      �?      �?      @      &@       @      4@              @                               @      &@      1@              @      @      (@      &@              �?      @       @       @      @               @               @              @               @                              @      @      �?                      "@              7@       @      I@      @      "@      @      (@      ;@      =@      @      3@      1@     �P@      D@              $@      @      *@      $@      5@       @      I@      @      "@      @      (@      ;@      =@      @      1@      1@     �P@     �A@              $@      @      *@       @       @                                                                               @                      @                                       @                      @       @      @      @      �?               @      �?      @      0@                              �?      @      �?       @                      @      �?      �?                                      �?      @      "@                              �?                                                      �?       @      @      �?               @                      @                                      @      �?       @                                              @      �?                                      @                                              �?       @                              �?       @                               @                      @                                      @                     �[@      (@      S@      $@      *@      @      .@     @b@     �c@      9@      0@      G@     �b@      V@      @      .@      2@      D@      @     �S@      @     �A@      @       @      �?      @     @]@     �Y@      @       @      7@     �W@     �C@              @      @      1@      @      0@               @      �?      �?      �?      @      .@      F@      @       @              *@      &@              �?               @      �?      .@              @      �?              �?       @      *@     �D@      @       @              $@       @              �?               @      �?      �?              @              �?              �?       @      @                              @      @                                              O@      @      ;@       @      @              @     �Y@     �M@       @      @      7@     @T@      <@               @      @      .@       @      .@              (@              �?              �?     �D@      ;@      �?      @      @      2@      ,@              �?              @      �?     �G@      @      .@       @      @              @     �N@      @@      �?      @      3@     �O@      ,@              �?      @      &@      �?      @@      "@     �D@      @      @      @       @      =@      L@      4@       @      7@     �L@     �H@      @      (@      (@      7@      @      8@      "@      0@      @      @      @      @      7@     �I@      .@       @      ,@      I@      @@      @      @      @      ,@      �?      5@      @      0@      @      @      @       @      0@     �B@      .@      @      &@      F@      ?@       @      @      @      (@      �?      @      @                                      @      @      ,@              @      @      @      �?       @      �?               @               @              9@       @                      @      @      @      @              "@      @      1@              @      "@      "@       @       @              1@       @                       @      @      @      @              "@      @      (@              @      "@       @       @                       @                              �?                                                      @                              �?             �Q@      3@      L@      (@      8@      (@      :@      :@     �S@      ,@      0@      E@     �R@     �V@      $@      *@      @      3@      2@     �G@      &@      B@       @      1@      $@      $@      5@     �L@      @       @      6@     �I@      D@      @      $@       @       @      "@      C@      $@      =@      @      1@      "@       @      3@     �G@      @       @      5@     �B@      B@      @      @      �?       @      "@      @@       @      <@      @      1@      "@       @      ,@      E@      @       @      4@      B@      <@      @      @      �?       @       @      1@      @      1@      @      .@      "@      @      "@      @@       @      @      *@      4@      3@      @      @      �?       @      @      .@      @      &@      �?       @               @      @      $@      @      @      @      0@      "@              �?                       @      @       @      �?      �?                              @      @                      �?      �?       @                                      �?      �?                                                      @      @                      �?              @                                              @       @      �?      �?                                      �?                              �?      @                                      �?      "@      �?      @      �?              �?       @       @      $@                      �?      ,@      @              @      �?                       @              @                              �?       @       @                              @      �?                                                              @                              �?      �?                                      @                                                       @              @                                      �?       @                              �?      �?                                              @      �?              �?              �?      �?               @                      �?      @      @              @      �?                      @                      �?                                      @                              �?                      @                                      �?                              �?      �?              @                      �?      @      @                      �?                      8@       @      4@      @      @       @      0@      @      6@       @       @      4@      7@     �I@      @      @      @      &@      "@      ,@              "@               @                      @      1@      @      @      "@      2@      <@               @       @      "@      @      @              @               @                      @      &@              @       @      @      *@               @      �?      @      @      @              @                                       @      @              @              �?      *@               @      �?      @      �?                                       @                      �?      @                       @      @                                      �?      @      $@              @                                              @      @              @      (@      .@                      �?       @              �?              @                                              �?                      �?      @      @                                              "@              �?                                              @      @              @      @      &@                      �?       @              $@       @      &@      @      @       @      0@       @      @      �?      @      &@      @      7@      @      �?      @       @      @      "@       @      &@       @      @       @      0@       @      @      �?      @      "@      @      7@      @      �?      @      �?       @      @      @      @              @       @      @      �?      @      �?      @      @      @      3@      �?      �?      @      �?       @      @       @      @       @      �?              &@      �?                      �?      @              @       @                                      �?                       @      �?                                                       @                      �?                      �?      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJdP*hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         6                    �? ��~���?�	           ��@                           �?[�^u��?           ��@                            �?G\2��?y           ��@                          �1@�E]t�?n             f@������������������������       ��Ҍ���?             7@       	                    �?�W�g��?a             c@                          �5@��ͽ1��?.            �R@������������������������       ��E��ӭ�?             B@������������������������       �cT!)��?             C@
                           @��~�\��?3            �S@������������������������       ��RN�ڷ�?'            �M@������������������������       ���(\���?             4@                           �?q���?           `z@                          �1@�N�'��?r            �e@                            @]ON���?             ;@������������������������       �>;n,��?             &@������������������������       �      �?	             0@                            �?������?b            �b@������������������������       ��L�y��?(            �N@������������������������       �R����?:            �U@                           @����?�            �n@                           @�X��'�?�             l@������������������������       ���P�	��?_            �b@������������������������       �4lF��=�?,            @S@                            @�ˠT�?             6@������������������������       ���E���?             "@������������������������       ��1G����?             *@       +                   �=@�S+ю.�?�           T�@       $                    �?�p����?Y           x�@       !                    �?��U�#o�?�            r@                           �2@���(\��?L             ^@������������������������       ��d�����?             3@������������������������       �u6��$�??            @Y@"       #                   �5@�8\3��?j             e@������������������������       ��q�Q�?:             X@������������������������       �>��^[��?0            @R@%       (                    �?|��h���?�           p�@&       '                    �?��2���?�            �o@������������������������       ����(\��?             $@������������������������       �?^!���?�            �n@)       *                     @�|?5^��?            y@������������������������       ��U�(���?�            �i@������������������������       ���g��?            �h@,       1                     �?��7i��?E            �Y@-       0                   @@@P1��w�?            �C@.       /                    @�|�j��?             >@������������������������       �n�����?             .@������������������������       �0��b�/�?             .@������������������������       ������H�?             "@2       3                     �?�MՕm�?/            �O@������������������������       �     ��?
             0@4       5                    @��;�?%            �G@������������������������       �G���t��?            �A@������������������������       ��q�q�?	             (@7       T                    �?VzĢ��?�           ��@8       E                   �2@h�(��?�           �@9       @                    @f	�/!��?�            �w@:       =                     @�z���?8            �V@;       <                     �?     t�?(             P@������������������������       �A�<;���?!            �J@������������������������       �t�E]t�?             &@>       ?                   �1@g�WH��?             ;@������������������������       �pƵHP�?             *@������������������������       ��X�C�?             ,@A       D                    @w�@����?�            �q@B       C                    @sW����?�            �p@������������������������       �,�ѳ��?Y             a@������������������������       �     �?J             `@������������������������       ���|���?             6@F       M                    @Ra�����?�            �@G       J                    @�u��:��?�            �s@H       I                   �=@��m{�?�            `m@������������������������       �H	��{�?�            �k@������������������������       �����>�?             ,@K       L                    @r����?-            @S@������������������������       �)\���(�?!             I@������������������������       �#����?             ;@N       Q                    @@$,�o��?           �x@O       P                    @�L�^	C�?�            pv@������������������������       ��Yqs��?�             h@������������������������       ���mjP��?q            �d@R       S                    @vK�B#��?            �@@������������������������       �}��7�?             &@������������������������       ��X����?             6@U       d                   �5@.Ĵ�x�?�           ��@V       ]                    @����_�?�           P�@W       Z                   �1@�3_<�?E           �@X       Y                   �0@�'���?f            �d@������������������������       �g\�5�?!             J@������������������������       �v�w�<0�?E            @\@[       \                   �2@�D�ς��?�            0u@������������������������       �fY�eY��?:             U@������������������������       �� ��P��?�            �o@^       a                   �3@�M��?h            @f@_       `                    @���~�?H             _@������������������������       �"n���?$            �Q@������������������������       ��i�+$��?$             K@b       c                     �?I��D�?              K@������������������������       �     ��?             @@������������������������       ��9����?             6@e       l                    @o���?B           �@f       i                     @���`��?�            �v@g       h                    @^�u6�?�            �r@������������������������       �z�-U_��?�             p@������������������������       �:(!�;\�?            �C@j       k                   �9@�>��DM�?+            @Q@������������������������       �F��ӭ��?             B@������������������������       �,j�J��?            �@@m       p                    �?b��7��?^            �a@n       o                   �:@      �?             @@������������������������       ���6�80�?             3@������������������������       �ƵHPS!�?             *@q       r                   �;@��5*q�?K            @[@������������������������       ��������?7             T@������������������������       �K�]l���?             =@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       P{@     �Q@     v@      E@     @Q@      A@     �R@     8�@      �@     �P@     �W@     �b@     Ȃ@     �{@      $@     �O@     �K@      ^@     @Q@     �f@     �B@     �e@      9@     �E@      9@      B@     �\@     `g@     �B@      L@     @R@     �o@     �i@       @      D@     �A@     �K@     �K@     @U@       @     �F@      �?      0@       @      (@     �O@      Q@      3@      6@      ?@     @Z@      P@              ,@      "@      (@      6@      8@      @      *@      �?      @       @      @      1@      &@      �?      @      "@      G@      1@              @      @      @      @      @                                                      $@       @                      @      �?      �?                                              2@      @      *@      �?      @       @      @      @      "@      �?      @      @     �F@      0@              @      @      @      @      *@      �?      @                                      �?       @      �?       @       @      :@      $@              �?       @      @      �?       @                                                      �?      @                       @      2@      @                                              @      �?      @                                              @      �?       @               @      @              �?       @      @      �?      @      @      $@      �?      @       @      @      @      �?              �?      @      3@      @              @       @      �?      @      @      @      @      �?      @       @      @      @                      �?      @      *@       @              �?       @      �?      @       @              @                              �?              �?                              @      @               @                             �N@       @      @@              &@               @      G@     �L@      2@      3@      6@     �M@     �G@              $@      @       @      1@      9@              *@              �?               @      @@      A@      @      @      @      >@      (@              @      �?      �?      @       @                                                      ,@      @      @                      �?                                                      �?                                                      @      @                                                                                      �?                                                      "@       @      @                      �?                                                      7@              *@              �?               @      2@      ;@      @      @      @      =@      (@              @      �?      �?      @      ,@              @              �?                      (@      (@      �?      @              @       @                                      @      "@              @                               @      @      .@      @      @      @      6@      $@              @      �?      �?      �?      B@       @      3@              $@              @      ,@      7@      &@      (@      3@      =@     �A@              @      @      @      *@      >@       @      ,@              $@              @      *@      7@      "@      (@      3@      6@     �A@              @      @      @      *@      4@       @      $@              @              @      &@      3@      @      @      "@      2@      ;@              @      �?       @      @      $@              @              @              @       @      @      @      @      $@      @       @                      @      @       @      @              @                                      �?               @                      @                                      �?              �?                                                                       @                      @                                      �?              @              @                                      �?                                       @                                                     @X@      =@      `@      8@      ;@      7@      8@      J@     �]@      2@      A@      E@     �b@     �a@       @      :@      :@     �E@     �@@     �V@      =@     �]@      4@      6@      .@      5@      J@     �]@      *@      6@     �C@     �b@     @a@      @      4@      1@      ?@      :@      C@       @      9@      @      (@      @      @      *@     �B@      @       @      &@      L@     �E@       @      �?      �?      .@      "@      1@      �?      "@      @       @              �?      @      0@               @      �?      >@      1@       @      �?              &@      �?      @                                                      @                                       @      @                              @              *@      �?      "@      @       @              �?              0@               @      �?      <@      *@       @      �?               @      �?      5@      @      0@      @      $@      @       @      @      5@      @              $@      :@      :@                      �?      @       @      ,@      @       @              @      �?      �?      @      4@      �?              @      (@      $@                      �?      @       @      @      @       @      @      @       @      �?              �?      @              @      ,@      0@                                      @      J@      5@     �W@      ,@      $@      (@      2@     �C@     @T@      "@      4@      <@      W@     �W@      �?      3@      0@      0@      1@      :@      @     �@@      @      @      @      @      ;@      A@              @      @      F@      >@              @       @      @      @                       @                                      @      �?                                      �?                                              :@      @      ?@      @      @      @      @      5@     �@@              @      @      F@      =@              @       @      @      @      :@      1@     �N@      $@      @       @      *@      (@     �G@      "@      ,@      5@      H@     @P@      �?      *@       @      $@      &@      ,@      @      ?@      @      @              @      &@      6@       @      &@      @      <@      >@               @      @      @      @      (@      ,@      >@      @               @       @      �?      9@      �?      @      ,@      4@     �A@      �?      @       @      @      @      @              "@      @      @       @      @              �?      @      (@      @       @      @      @      @      "@      (@      @      @                      �?              @                      �?              &@       @               @                      @      "@      �?      @                      �?              @                      �?               @                       @                       @       @              @                      �?                                      �?               @                                                       @                                                      @                                      @                       @                       @                      �?                                                                              @       @                                      �?      �?      �?      @              "@      @      @      @      @                      @      �?      �?       @       @      @      @      @      @      @                      @      �?                      �?                      @              �?                               @      �?      @              @              @       @      @      @       @                       @      �?               @       @      @      @      @              @      @              @      �?       @      @       @                       @      �?                       @      �?      @      @              @                              �?      @                                                               @              @               @                     �o@      A@     �f@      1@      :@      "@      C@     @{@     �z@      =@     �C@      S@     �u@     �m@       @      7@      4@     @P@      ,@      _@      &@     �S@      �?      @      �?      &@     �p@     �k@      &@      2@      :@     �d@     @X@              @      @      =@      @      E@      �?      3@                               @      a@     �W@      @      �?      @     �F@      9@                              �?              0@              @                                      1@      =@      �?      �?      �?      *@       @                              �?              @              @                                      1@      ;@              �?      �?      @      @                              �?              @              @                                      0@      4@              �?      �?       @      @                              �?                              �?                                      �?      @                               @                                                      (@                                                               @      �?                      "@      @                                              @                                                              �?      �?                      @                                                       @                                                              �?                               @      @                                              :@      �?      .@                               @     �]@     �P@      @              @      @@      1@                                              4@      �?      .@                               @     �Z@     �P@      @              @      >@      1@                                               @              "@                                     �J@      C@                      @      5@      @                                              (@      �?      @                               @     �J@      <@      @              �?      "@      *@                                              @                                                      *@                              �?       @                                                     �T@      $@      N@      �?      @      �?      "@     �`@     �_@      @      1@      4@     �^@      R@              @      @      <@      @     �H@      @      1@              @      �?      @     �H@      L@      @      @      *@     �J@      A@                       @      .@      �?      E@      @      (@              @      �?      @      B@      I@      �?      @      &@      C@      4@                               @      �?     �D@      @      (@               @      �?      @     �A@      H@      �?       @      &@      >@      4@                               @      �?      �?                              �?                      �?       @              �?               @                                                      @       @      @                              �?      *@      @      @               @      .@      ,@                       @      @              @       @      @                                       @      @      �?               @      @       @                       @      @              �?               @                              �?      @       @       @                       @      @                                             �@@      @     �E@      �?      �?               @     �T@     �Q@      @      ,@      @     @Q@      C@              @      �?      *@      @      =@      @      C@      �?                              T@     �P@      @      ,@      @     �P@      A@              @              $@      �?      .@      @      4@                                     �J@      ?@       @      @       @      D@      .@              �?              @      �?      ,@      �?      2@      �?                              ;@      B@      �?       @      @      :@      3@              @              @              @      �?      @              �?               @      @      @                              @      @              �?      �?      @       @                      @              �?                      @      �?                                                              �?                      @      �?                                       @               @                              @      @              �?              @       @     ``@      7@     @Y@      0@      6@       @      ;@      e@     �i@      2@      5@      I@     `f@     `a@       @      1@      1@      B@      $@     @W@      @     �E@      @       @      �?      (@     `a@     @b@      �?      "@      8@     @Z@     �O@              @      @      &@      @     �S@      @      >@      @       @      �?       @     �\@     �V@      �?      @      2@     @U@      E@              @      @      @      @      5@              @                              �?      F@      E@              @       @      :@      $@                               @      �?      @              �?                                      1@      $@                      �?      &@      @                               @              ,@              @                              �?      ;@      @@              @      @      .@      @                                      �?     �L@      @      7@      @       @      �?      @     �Q@     �H@      �?      @      $@     �M@      @@              @      @      @      @      *@      �?      @                               @      9@      �?      �?                      7@      @              �?       @      �?       @      F@      @      2@      @       @      �?      @     �F@      H@              @      $@      B@      9@               @      @      @      �?      .@      @      *@       @      @              @      9@     �K@              @      @      4@      5@                              @               @               @      �?      @              �?      .@     �G@                      @      (@      3@                              @              @              @      �?      @              �?       @     �B@                      �?      @       @                              �?              @              @                                      *@      $@                      @      @      &@                              @              @      @      @      �?      �?              @      $@       @              @       @       @       @                              �?               @              @      �?      �?                      @       @              @               @       @                              �?              @      @                                      @      @                               @      @                                                      C@      0@      M@      "@      ,@      @      .@      =@      M@      1@      (@      :@     �R@      S@       @      ,@      &@      9@      @      8@      $@     �@@      @      $@      @      &@      8@      I@      (@      (@      6@     �L@      L@       @      "@      @      .@       @      4@      @     �@@      @      "@      @      @      2@      B@      &@      (@      1@      J@     �B@      �?      @      @      *@              1@      @      =@       @      @      @      @      1@     �A@      &@      $@      1@      H@      ?@      �?      @      @      @              @              @      @      @              �?      �?      �?               @              @      @              �?              @              @      @                      �?              @      @      ,@      �?              @      @      3@      �?       @               @       @       @                                               @      @      (@                       @      @      @                               @      �?       @      @                      �?               @      �?       @      �?              @       @      (@      �?       @                      �?      ,@      @      9@      @      @              @      @       @      @              @      1@      4@              @      @      $@      @              @      @              �?                      �?      @      �?              �?      @      @              @       @       @      @               @      @              �?                      �?      �?      �?                      @       @              @       @                               @                                                      @                      �?               @                               @      @      ,@       @      6@      @      @              @      @      @      @              @      ,@      0@               @      @       @      �?      $@       @      2@              @               @      @      @       @               @       @      0@               @      @      @              @              @      @                       @                       @              �?      @                               @      @      �?�t�bub�R     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJC(chG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKkhnh4h7K ��h9��R�(KKk��hu�Bh         4                   �2@=G�?R��?�	           ��@                           �?�i���?�           ��@                           �?�����?�            �t@                           @��H����?]            `a@                            �?ȶ���?W            �_@                           �?]"?ӧ
�?/             O@������������������������       �����?             C@������������������������       �r�q��?             8@	       
                    �?;2C+6��?(            @P@������������������������       ���QN�?             ?@������������������������       �~2�P�?             A@������������������������       �9��8���?             (@                           �?����?s             h@                          �1@4և����?&             L@                            @V>�� =�?             ?@������������������������       ���]�`��?
             *@������������������������       �O��E�?
             2@                            �?�A`��"�?             9@������������������������       �}��7�?             &@������������������������       �s
^N���?
             ,@                          �0@��y�b��?M             a@������������������������       �R���Q�?             4@                            @K�~�y��?B            @]@������������������������       �Դ��K.�?#            @Q@������������������������       ���8���?             H@       )                    @����"o�?�            �@       "                    @,��h��?e           8�@                           @M�ة���?i            @d@                           �?�z����?L            �^@������������������������       ����.��?/            �S@������������������������       �U�x?r��?             F@        !                   �0@ffffff�?             D@������������������������       ������?             3@������������������������       ��E�_���?             5@#       &                     @|B]�?�            Px@$       %                    @g������?�            �s@������������������������       �]pOx�:�?�            �j@������������������������       ������?=            �X@'       (                   �1@��Դ��?2             S@������������������������       ��D[�� �?            �H@������������������������       � ��?Z�?             ;@*       1                     @z7e�?Q            @_@+       .                     �?�-�2�7�?A            �Y@,       -                    @�������?!            �I@������������������������       �Dc}h��?             <@������������������������       ��C4T2�?             7@/       0                    �?*Mp���?             �I@������������������������       �"�����?             5@������������������������       � d��0u�?             >@2       3                    �?J��LQ�?             7@������������������������       ���"e���?             "@������������������������       ��m۶m��?
             ,@5       R                   �8@��c���?M           ��@6       C                    �?��0_���?�           ̞@7       >                   �7@J������?@           (�@8       ;                     �?d�50K��?�           ��@9       :                    �?���x��?           �y@������������������������       �����KF�?`            �b@������������������������       ��m��1�?�            @p@<       =                    @�����?�            �u@������������������������       �ǽq���?�            �m@������������������������       ��o5���?J            @[@?       B                    @����~�?H             \@@       A                    @�m�|,�?A            �Y@������������������������       �����[��?+             R@������������������������       �c�/��b�?             >@������������������������       �R���Q�?             $@D       K                    �?NB6�j��?�           8�@E       H                    @�]�?�?�             w@F       G                   �7@?�ܵ�|�?�             i@������������������������       �2�����?o            `e@������������������������       �f"΃�?             =@I       J                    @��8Yz�?k            @e@������������������������       ��Q�	"�?<            �X@������������������������       �����S��?/            �Q@L       O                    @(4	���?�           ��@M       N                     @���Aq��?�           �@������������������������       �r7-���?)           @~@������������������������       �趶����?�            �k@P       Q                   �4@�������?             9@������������������������       ���E���?             "@������������������������       �     @�?             0@S       \                    �?T��n%��?]           0�@T       [                    @�F/((�?�            �j@U       X                   �;@�ob����?}             h@V       W                    �?ڭ)x��?F            �Z@������������������������       �f|�We��?!            �J@������������������������       ��?����?%             K@Y       Z                    �?Uj ��k�?7            �U@������������������������       �\��[���?            �C@������������������������       �*�6(���?            �G@������������������������       ��V���?             6@]       d                    �?[Q�f6��?�           x�@^       a                    @�FqS1�?�            `o@_       `                     �?�[ A�c�?"             I@������������������������       �R�n��?             2@������������������������       �     ��?             @@b       c                     �?6�>����?�             i@������������������������       ���C~���?M            @[@������������������������       �$e?��Z�??             W@e       h                   @@@�ҧ���?           @}@f       g                    @�u���d�?�            @y@������������������������       �-V�T<�?�            r@������������������������       ��Ty���?P            �\@i       j                     �?     <�?#             P@������������������������       �     ��?             @@������������������������       �     0�?             @@�t�bh�h4h7K ��h9��R�(KKkKK��h��B�?       P|@     �V@     Pv@      =@      T@      =@      V@     ؀@      �@     �P@      V@     �d@     8�@     z@      *@      R@     �B@     �`@      N@     �`@      @     �M@              @              $@     `q@     �i@      @      @      7@     @d@      S@              (@       @      8@      @     �J@              >@               @              @      O@      D@      @      �?      .@     �M@      C@              @      �?      3@       @      :@              "@                               @      B@      3@                       @      5@       @              @              @              6@              @                               @      B@      3@                       @      3@       @              �?              @              1@              �?                                      6@      (@                      @      @       @                                              "@              �?                                      .@      @                      @       @      �?                                               @                                                      @      @                              @      �?                                              @              @                               @      ,@      @                      @      ,@      @              �?              @              @              @                                      @      @                      @      @      �?              �?              �?              �?              �?                               @      $@      �?                       @       @      @                              @              @               @                                                                               @                       @               @              ;@              5@               @               @      :@      5@      @      �?      @      C@      >@                      �?      (@       @      @               @                               @      @      @      �?              @      (@      @                              @              @              @                                      @      �?      �?              @      @      @                               @              @                                                       @      �?      �?              @      @                                                       @              @                                      @                                      @      @                               @               @              @                               @      �?      @                              @      @                               @                              @                                               @                               @                                       @               @                                               @      �?       @                              @      @                                              4@              *@               @                      3@      0@       @      �?      @      :@      7@                      �?       @       @      $@              �?                                      @                                              @                                              $@              (@               @                      *@      0@       @      �?      @      :@      4@                      �?       @       @      @              @              �?                      (@      "@       @              @      3@      @                              @       @      @              @              �?                      �?      @              �?      �?      @      ,@                      �?      @             �T@      @      =@              �?              @      k@     �d@      @       @       @     �Y@      C@              "@      �?      @      �?      L@       @      ;@              �?              @      h@     �`@      @       @      @     �T@      @@              �?      �?      @      �?      3@              @                               @     �C@     �J@      @               @      5@      $@              �?      �?      @              .@              @                               @      C@      =@       @               @      2@      @              �?      �?      @              (@              �?                                      >@      4@                              $@       @                              @              @              @                               @       @      "@       @               @       @      @              �?      �?                      @              �?                                      �?      8@      �?                      @      @                              �?                                                                      �?      ,@                               @       @                                              @              �?                                              $@      �?                      �?      @                              �?             �B@       @      4@              �?              @      c@     @T@               @      @      O@      6@                                      �?      5@       @      &@                              @     �`@     �P@                      @      J@      5@                                               @       @      @                              �?      Y@     �I@                      �?      B@      &@                                              *@              @                               @      @@      .@                      @      0@      $@                                              0@              "@              �?                      5@      .@               @              $@      �?                                      �?       @                              �?                      4@      ,@               @              @      �?                                               @              "@                                      �?      �?                              @                                              �?      :@      @       @                              �?      8@      ?@      �?              �?      4@      @               @              �?              :@      @      �?                              �?      2@      9@      �?              �?      *@      @              @              �?              &@      @                                      �?      *@      (@                      �?       @                                      �?              @       @                                      �?      @       @                              @                                                      @       @                                              "@      @                      �?      �?                                      �?              .@              �?                                      @      *@      �?                      @      @              @                              @                                                      @      @      �?                       @       @                                              "@              �?                                       @      @                              @       @              @                                              �?                                      @      @                              @       @              �?                                              �?                                      @      �?                               @      �?                                                                                                       @      @                              @      �?              �?                             �s@     @U@     �r@      =@     @S@      =@     �S@     Pp@     py@      N@     @U@     �a@     Pz@     Pu@      *@      N@     �A@     @[@     �L@     �m@      H@     @i@      3@      >@      &@     �C@     �k@     �t@      =@     �H@     �U@     �r@      m@      @      6@      1@     �P@      ?@     @[@      $@     �Q@      �?      "@      �?      $@     @]@     �d@      &@      3@      >@     `d@     @W@              "@      "@      ?@      &@     �Y@      @      M@              "@      �?      @     �Y@     �a@       @      1@      :@     �c@     �S@              @      @      ;@      @     �N@      @     �@@              @              @     �F@      U@      @      *@      "@     @U@     �D@              @       @      ,@       @      :@      �?      *@              @              �?      "@      0@      �?      @       @     �D@      4@              @              @       @     �A@       @      4@                              @      B@      Q@      @      @      @      F@      5@                       @      "@              E@      @      9@              @      �?             �L@     �L@       @      @      1@     �Q@      C@               @      @      *@      @     �C@      @      .@               @      �?              E@      D@       @      @      "@      B@      >@               @       @      @      @      @              $@              @                      .@      1@              �?       @     �A@       @                       @      @              @      @      *@      �?                      @      .@      8@      @       @      @      @      ,@              @      @      @      @      @      @      *@      �?                      @      (@      8@      @       @      @      @      ,@               @       @      �?      @      @      @      &@      �?                      @      @      3@               @      @      @      @               @       @              @      �?               @                              �?      "@      @      @                               @                              �?                                                                      @                                       @                      �?      �?      @             �_@      C@     ``@      2@      5@      $@      =@      Z@     �d@      2@      >@     �L@     �`@     �a@      @      *@       @     �A@      4@      F@      @      :@      �?      @      @      @      G@     @R@      @      @      ,@     �F@      M@               @      @       @      @      6@      @      0@              @      @      @      ,@     �E@      @      @      &@      9@      9@              @      �?      @      �?      5@      @      (@              @      @      @      ,@      D@      @      @      "@      2@      *@              @      �?      @      �?      �?              @                                              @                       @      @      (@                                              6@       @      $@      �?                       @      @@      >@                      @      4@     �@@              @       @       @      @      "@      �?       @      �?                              :@      2@                      @      $@      8@                                      @      *@      �?       @                               @      @      (@                              $@      "@              @       @       @      �?     �T@      @@     @Z@      1@      .@      @      7@      M@      W@      (@      8@     �E@     @V@     �T@      @      @      @      ;@      *@      T@      @@     �Y@      (@      .@      @      1@      M@      W@      (@      7@     �E@      V@     �R@      @      @      @      ;@      *@     �K@      3@     �Q@      @      $@              &@     �I@      O@      @      ,@      ?@      Q@     �D@      �?      @      @      3@      (@      9@      *@     �@@      @      @      @      @      @      >@      @      "@      (@      4@      A@      @               @       @      �?      @               @      @                      @                              �?              �?      @                                              �?               @                                                                              �?      @                                               @                      @                      @                              �?                       @                                             �T@     �B@      X@      $@     �G@      2@     �C@      D@     @S@      ?@      B@     �K@      _@      [@      "@      C@      2@     �E@      :@      <@      "@      &@      @      @      @      "@       @      :@      @      (@      $@      ?@      =@       @      "@      �?       @      @      <@      "@      &@      @      @      @      @       @      7@      @      (@      "@      >@      9@       @       @      �?       @       @      5@      @      @      �?      @      �?      �?      �?      *@              �?      @      4@      1@       @      @              @      �?      $@      @      �?                                              *@              �?      @      $@      @               @               @              &@       @      @      �?      @      �?      �?      �?                              �?      $@      &@       @      @               @      �?      @      @      @       @      �?      @      @      �?      $@      @      &@      @      $@       @              @      �?      @      �?      @      �?      @                              �?      �?      @              @      �?      @      @              @                              @       @      @       @      �?      @      @              @      @      @      @      @       @                      �?      @      �?                                      �?               @      @      @       @              �?      �?      @              �?                      �?      K@      <@     @U@      @      E@      *@      >@      @@     �I@      9@      8@     �F@     @W@     �S@      @      =@      1@     �A@      7@      9@      *@      5@      �?       @              *@      4@      ;@       @      $@      @      D@      =@              "@      @      &@      &@       @      �?      &@               @              @      @      �?       @      �?      �?      @      @              @      �?      @              @      �?      �?                              @      �?              �?      �?                                       @              @              @              $@               @                       @      �?      �?              �?      @      @               @      �?                      1@      (@      $@      �?      @              "@      1@      :@              "@      @     �B@      8@              @      @       @      &@      "@      @      @              �?               @      &@      0@              @      @      ,@      3@              @       @      @      "@       @       @      @      �?      @              @      @      $@              @              7@      @               @      @       @       @      =@      .@      P@      @      A@      *@      1@      (@      8@      7@      ,@      D@     �J@      I@      @      4@      &@      8@      (@      :@      *@      M@      @      A@      "@      0@      (@      7@      7@       @      8@     �I@     �H@       @      2@      @      0@      "@      *@      &@      F@      @      8@       @      @      (@      5@      7@      @      2@     �C@      @@      �?      &@      @      *@      @      *@       @      ,@       @      $@      �?      (@               @              @      @      (@      1@      �?      @      @      @      @      @       @      @                      @      �?              �?              @      0@       @      �?      @       @      @       @      @       @                                              �?              �?              @      &@       @                      �?       @      @      �?      �?       @      @                      @                                      �?      @              �?      @      �?       @       @       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�"hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKuhnh4h7K ��h9��R�(KKu��hu�B�         >                   �2@�6�Ț��?�	           ��@                           �?<Y�/��?�           x�@                           @4ٹ<S�?J           ��@                           �?��g\���?�            `l@                           �?-�%�xE�?5            �U@                          �1@9��8���?             8@������������������������       �؂-؂-�?	             .@������������������������       �0�����?             "@	       
                     �?�+Z���?%            �O@������������������������       �     ��?             @@������������������������       ���b�=�?             ?@                            �?x9/���?T            �a@                            �?���Z��?)            @P@������������������������       �g�W���?             A@������������������������       �R�5�`��?             ?@                           �?��ݓ���?+            �R@������������������������       �ZZZZZZ�?             �I@������������������������       ��q�q�?             8@                           @�!T_��?�            �s@                          �1@̄���?�            �n@                            �?��(\���?a             d@������������������������       �2��=��?            �B@������������������������       �t�W��w�?L            �^@                            �?3,Ң�?5            �U@������������������������       �贁N��?             >@������������������������       ��>4և��?#             L@                            @�ە%��?+            @Q@                          �0@�lÎ��?$             M@������������������������       �b���i��?             &@������������������������       �����<�?            �G@������������������������       �}��7�?             &@        /                    @    `��?7            �@!       (                    @6��ԭ�?�            �r@"       %                     @�/�eo��?�            �k@#       $                    �?�~��?F             [@������������������������       �'�Tk��?            �F@������������������������       ��#Y�'�?*            �O@&       '                   �1@�#�d��??            @\@������������������������       ��~���B�?&            �N@������������������������       �^�`���?             J@)       ,                     �?�\�>$��?9            �T@*       +                    �?~e�.y0�?$             J@������������������������       ��ƖJ��?             ?@������������������������       ��T�	��?             5@-       .                    @�z�G��?             >@������������������������       ��������?             2@������������������������       �UUUUUU�?             (@0       7                    @�h�*$��?y             j@1       4                   �0@#��U��?N            @`@2       3                    @E�ϣ1��?             C@������������������������       ��T�	��?             5@������������������������       ��W��H��?             1@5       6                    @UP��g��?;             W@������������������������       ��y})�?            �G@������������������������       �>M�k%�?            �F@8       ;                    @�s�Z���?+            �S@9       :                     �?{���CA�?             O@������������������������       ����З�?            �C@������������������������       �\")�i��?             7@<       =                     �?�@�m�?             1@������������������������       ��(\����?             $@������������������������       �������?             @?       V                    �?gb�q��?           V�@@       I                    �?�s��=\�?           X�@A       H                   �?@��*���?           0}@B       E                    �?�zQ7���?           P|@C       D                    �?�	U��6�?Q             a@������������������������       ��H6��%�?.            @R@������������������������       �&7)��?#            �O@F       G                    �?�n:o��?�            �s@������������������������       �N�zv�?C            �[@������������������������       �9�\@��?z            �i@������������������������       ���>4և�?             ,@J       Q                   �@@����p�?           �@K       N                    �?T�pN�?�           �@L       M                    �?=c��#��?�            �s@������������������������       �>α�
��?H            �Z@������������������������       �Ȩ�I��?�            �j@O       P                   �>@��(K|�?           �y@������������������������       �Ƿdp�a�?           �x@������������������������       ���a_j�?             3@R       S                   @A@�].��?             C@������������������������       ���8��8�?             (@T       U                     @θ	�?             :@������������������������       ���(\���?             $@������������������������       �     ��?
             0@W       f                     @�៻d_�?�           T�@X       _                    �?#�M�E�?E           �@Y       \                   �7@gC�t���?}           0�@Z       [                    @�������?           �y@������������������������       ��!!pϯ�?�            �w@������������������������       ��Cc}�?             <@]       ^                    �?_�E�x�?x            �i@������������������������       ��S@ذ�?'            �P@������������������������       �)��ח�?Q            `a@`       c                     �?j�]ث�?�           ��@a       b                    @���\��?�            �p@������������������������       �.�-�c�?3            �V@������������������������       �x<���?j            @f@d       e                   �:@�M�7H�?+           �|@������������������������       ���Զ|��?�            x@������������������������       ���[��"�?.             R@g       n                    @���l�?�            �q@h       k                   �5@p���r�?\            �a@i       j                    @ÇՊ~��?,            �L@������������������������       ��Sy'��?#             E@������������������������       ��������?	             .@l       m                   �;@      �?0             U@������������������������       �     ��?%             P@������������������������       �\���(\�?             4@o       r                   �3@8��!n��?[            �a@p       q                    �?�A`��"�?             9@������������������������       �ƵHPS!�?             *@������������������������       �r�q��?	             (@s       t                    @���/�#�?G            �\@������������������������       ���ӭ�a�?             B@������������������������       ��)���?4            �S@�t�bh�h4h7K ��h9��R�(KKuKK��h��BxE        {@      U@     �u@      B@     �S@      :@     @Q@     P�@     �@     �R@      X@     �c@     ��@     @y@      3@     �M@     �G@      `@     �L@     @^@      $@     �R@      @      @              *@     �q@     `k@      @      "@      7@     `e@     �R@              "@      @      8@      @     �M@      @      9@                              @     �f@      `@              @      "@     �R@      B@              @              &@             �@@              &@                                      L@      H@              @      @     �D@      .@              @              &@              2@               @                                      9@      @               @       @      0@      @               @              @              @               @                                       @       @                       @               @               @              �?              @               @                                      @      �?                       @              �?                                               @                                                       @      �?                                      �?               @              �?              *@                                                      1@      @               @              0@      @                              @              @                                                      .@       @               @              @       @                                              @                                                       @       @                              (@      @                              @              .@              "@                                      ?@      E@               @      �?      9@       @              @              @              "@              �?                                      (@      <@               @              "@       @                               @              @              �?                                       @      $@                              "@                                       @              @                                                      @      2@               @                       @                                              @               @                                      3@      ,@                      �?      0@      @              @               @               @              @                                      0@      @                      �?       @      @              @               @              @               @                                      @      @                               @                                                      :@      @      ,@                              @     �_@     @T@                      @     �@@      5@                                              1@      @      "@                              @      [@      P@                      �?      :@      ,@                                              &@      @      @                              @     �S@     �D@                              0@      @                                              @                                               @      5@      &@                                                                                       @      @      @                               @     �L@      >@                              0@      @                                              @              @                                      >@      7@                      �?      $@      $@                                              �?                                                      @      0@                      �?      @      @                                              @              @                                      ;@      @                              @      @                                              "@              @                                      3@      1@                      @      @      @                                               @               @                                      ,@      0@                      @      @      @                                              @                                                      @      @                              �?                                                      @               @                                      &@      *@                      @      @      @                                              �?              @                                      @      �?                              �?                                                      O@      @      I@      @      @              "@     @Y@     �V@      @      @      ,@     @X@     �C@              @      @      *@      @     �C@      @      B@      @      @              @      E@      H@      @      @       @      Q@      :@              �?      @      @       @      @@      @      :@      @      @              @      ?@      :@       @      @      @      K@      0@              �?      @      @               @      �?      &@              �?              @      3@      .@       @      �?      @      ?@      @                      @       @              @               @                                      .@      (@              �?      �?       @      �?                               @              @      �?      "@              �?              @      @      @       @              @      7@      @                      @                      8@      @      .@      @      @                      (@      &@              @              7@      (@              �?      �?       @              ,@              @              @                      &@      @               @              "@       @              �?      �?                      $@      @       @      @                              �?      @              �?              ,@      @                               @              @              $@              �?                      &@      6@      �?      �?       @      ,@      $@                              �?       @                      @                                      $@      4@      �?               @      &@      @                                                               @                                      $@       @      �?               @      @       @                                                              @                                              (@                              @      �?                                              @              @              �?                      �?       @              �?              @      @                              �?       @      @              @              �?                               @                              �?      @                              �?       @       @               @                                      �?                      �?               @      @                                              7@      @      ,@                              @     �M@      E@                      @      =@      *@              @       @       @      �?      &@              $@                               @      H@      =@                      @      *@      $@                              �?      �?                                                              9@      @                              �?      @                              �?                                                                      &@      @                                      @                                                                                                      ,@                                      �?      �?                              �?              &@              $@                               @      7@      6@                      @      (@      @                                      �?      @              "@                                      (@      @                      �?      $@      @                                              @              �?                               @      &@      2@                      @       @      �?                                      �?      (@      @      @                              @      &@      *@                      �?      0@      @              @       @      @              &@      @      @                              @      $@      &@                              *@      @                              @              &@      @                                      @      @      @                              @      �?                              @                              @                                      @      @                              "@       @                                              �?                                                      �?       @                      �?      @                      @       @      @                                                                               @                      �?                               @       @      @              �?                                                      �?                                      @                      �?              �?             �s@     �R@     0q@     �@@     @R@      :@      L@     �p@     `x@     �Q@     �U@     �`@     �|@     �t@      3@      I@      D@      Z@      K@     ``@      ?@     �a@      (@     �J@      6@      >@     @P@     @_@      =@     �O@      Q@     `d@      c@      *@     �@@      9@      H@     �A@      L@      &@     �C@       @      6@      @      $@      @@     �J@      "@      3@      5@      V@     �H@              "@      ,@      (@      1@      K@      &@     �C@       @      0@      @      $@      @@      J@      "@      .@      4@      V@     �H@              "@      ,@      (@      1@      0@      @       @              @              @      "@      @@              @       @      3@      .@              @      @      �?      @      @      @      @                                      @      =@              @       @      *@      @                                       @      &@              @              @              @      @      @              �?              @      &@              @      @      �?      @      C@      @      ?@       @      &@      @      @      7@      4@      "@      "@      2@     @Q@      A@              @      "@      &@      &@      *@       @      @               @      @       @      &@      *@       @      @      @      =@      "@              @       @      @       @      9@      @      9@       @      "@              @      (@      @      @      @      .@      D@      9@              �?      @      @      "@       @                              @                              �?              @      �?                                                             �R@      4@     @Y@      $@      ?@      2@      4@     �@@      R@      4@      F@     �G@     �R@     �Y@      *@      8@      &@      B@      2@     �R@      4@     �X@      "@      9@      2@      4@     �@@     �Q@      2@     �E@     �C@     �R@     �Y@      @      8@      &@     �A@      (@     �F@      @      G@      �?      $@      @      @      2@     �C@              4@      0@      E@      C@      �?      @      @      &@      @      9@       @      $@              @              �?      �?      &@               @      @      4@      *@      �?       @              @      �?      4@      @      B@      �?      @      @      @      1@      <@              (@      (@      6@      9@               @      @      @      @      =@      ,@     �J@       @      .@      .@      *@      .@      @@      2@      7@      7@     �@@     @P@      @      4@      @      8@      @      =@      ,@     �J@      @      ,@      "@      *@      .@      @@      .@      6@      7@     �@@     �O@      @      2@      @      8@      @                               @      �?      @                              @      �?                       @               @                       @      �?               @      �?      @                              �?       @      �?       @                      "@                      �?      @      �?              �?              @                                                       @                      �?                      �?      @                      �?      �?      @                              �?       @      �?      @                       @                              @                      �?      �?                                      �?       @              @                                                                                              @                                              �?      �?                       @                              @     �f@     �E@     �`@      5@      4@      @      :@     �i@     �p@      E@      8@     �P@     �r@      f@      @      1@      .@      L@      3@     �c@     �A@     @]@      1@      1@       @      4@     �f@     �l@      C@      3@      J@     �n@     @_@       @      0@      (@      D@      *@     @S@      *@     �D@      @      @              @     @Z@      `@      ,@      &@      3@     �\@     �I@              @       @      ,@      @      I@      @      6@               @              �?     �P@      Z@       @      @      ,@     �U@      <@                       @      $@      @      H@      @      5@               @              �?     �N@     �Y@      @      @      ,@      S@      <@                      �?       @      @       @              �?                                      @      �?      @                      &@                              �?       @              ;@       @      3@      @      @              @      C@      8@      @      @      @      <@      7@              @              @      �?      0@       @      @                                      $@      ,@      �?       @       @       @      @              �?                              &@      @      .@      @      @              @      <@      $@      @      @      @      4@      0@              @              @      �?     @T@      6@      S@      ,@      $@       @      0@      S@     �Y@      8@       @     �@@     @`@     �R@       @      $@      $@      :@      "@      4@      @     �A@      "@      @       @      *@      :@      8@      *@      @       @      I@      9@              @      @      .@       @       @              1@      @       @       @       @      @       @      �?      @      @      2@      @                       @      @              (@      @      2@      @      @              @      3@      0@      (@      @      @      @@      6@              @      @      &@       @     �N@      1@     �D@      @      @              @      I@     �S@      &@      �?      9@      T@     �H@       @      @      @      &@      @     �H@      $@      :@      @      @              @      I@     �R@      @      �?      3@     �Q@      F@       @      @      @      @      @      (@      @      .@       @                                      @      @              @      "@      @                       @      @      �?      8@       @      2@      @      @       @      @      8@      A@      @      @      ,@     �J@      J@      @      �?      @      0@      @      ,@      @      "@      @       @      �?       @      @      9@      �?              "@      7@      6@      �?              @      "@      @      @       @      @              �?      �?      �?      @      $@                      @      *@      @                      @       @              @       @      @              �?      �?              @       @                       @       @      @                              �?              �?                                              �?               @                       @      @                              @      �?              @       @       @      @      �?              �?      @      .@      �?              @      $@      3@      �?                      @      @      @               @      @      �?              �?      @      $@                      @       @      1@                              @      @      @       @                                                      @      �?              �?       @       @      �?                      @              $@      @      "@      �?      �?      �?      @      1@      "@      @      @      @      >@      >@      @      �?              @              @               @                               @              @              @      @      �?      @                                              �?                                              �?              @              @      �?      �?      @                                               @               @                              �?              @                      @              �?                                              @      @      @      �?      �?      �?       @      1@      @      @       @      �?      =@      :@      @      �?              @               @              @      �?                              (@      �?               @              "@      @                              �?              @      @      @              �?      �?       @      @       @      @              �?      4@      6@      @      �?              @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��zhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKohnh4h7K ��h9��R�(KKo��hu�BH         >                     @P{�d��?�	           ��@                           �?�Tn�f�?�           ��@                           @Ė�k}��?2           ē@                           �?��\��-�?�           ��@                           @��vD=x�?�            �x@                           �?�3��2s�?�            @s@������������������������       ��"�F�?h            �d@������������������������       ��e�	��?^            �a@	       
                     �?���5S��?1            �U@������������������������       ��~VC�1�?             E@������������������������       ����i�V�?             F@                            �?��堭^�?�            Pu@                          �4@��@�?�             q@������������������������       �     z�?R             `@������������������������       ��b���?Z            @b@                          �;@��HIc�?.            �P@������������������������       �\;U���?'             M@������������������������       ���"e���?             "@                           @�G�P�r�?a           ��@                          �0@_6��Z�?C           �~@                           @ֱ߹���?%            �L@������������������������       ��>$�*��?            �D@������������������������       �     @�?             0@                            �?����.��?            {@������������������������       ��3�`���?�            �r@������������������������       ��8"C��?_             a@                          �2@�7���?            �C@������������������������       �     ��?             0@                            �?��/��@�?             7@������������������������       �ffffff�?             $@������������������������       ��T�6|��?             *@        /                   �4@Q�5���?�           p�@!       (                    �?Ph���?�           �@"       %                     �?�F��41�?y            �g@#       $                    @�mdG�+�?9            @W@������������������������       ������?             �J@������������������������       ��������?             D@&       '                    �?3�l��N�?@            �X@������������������������       �#8̺�8�?             G@������������������������       �PS!����?"             J@)       ,                    @�~70���?           @|@*       +                    �?"Q5��?�            `u@������������������������       �}<��Z�?C            @Z@������������������������       ��@Wx|��?�            �m@-       .                    �?L��a���?F            �[@������������������������       �m��1G�?!             J@������������������������       �^s]ev�?%             M@0       7                   �;@_�J��H�?)           Ȋ@1       4                    �?r@_N_��?�           ��@2       3                    @-w�Ǒ�?�            �q@������������������������       ��Dn���?k            @e@������������������������       ���z����?E            @\@5       6                     �?
}���?�            pw@������������������������       ���VBwI�?R            @_@������������������������       ���$?�W�?�            @o@8       ;                   @A@�gE��?�            �h@9       :                   @@@2���|�?l            �d@������������������������       ���'#��?c            �b@������������������������       �����H�?	             2@<       =                    �?,j�J��?            �@@������������������������       �J�w�"w�?             3@������������������������       �4և����?             ,@?       V                    �?D�a���?�           �@@       M                    �?���O2�?�           ��@A       F                    �?.C�*��?�            �q@B       E                   �7@�G�z��?7             T@C       D                   �6@�	4-���?'            �J@������������������������       ��	j*D�?            �C@������������������������       �d}h���?             ,@������������������������       �'��}��?             ;@G       J                   �4@vq���?�             i@H       I                    @}����i�?6            �V@������������������������       �ҽe�J�?             E@������������������������       ��q�q�?             H@K       L                    �?�
����?L            �[@������������������������       �`����x�?             =@������������������������       �����!s�?8            �T@N       O                   �0@H�D�>�?           Pz@������������������������       ���8��8�?             (@P       S                    �?f~�ϐ>�?           �y@Q       R                   �7@/�����?P            �`@������������������������       ��zv��?7             V@������������������������       �-�D���?            �F@T       U                    @p<�54�?�            @q@������������������������       �Z0Rb�?I             ]@������������������������       ���Q�5�?l             d@W       d                   �5@B�����?           �{@X       ]                   �3@;)�%�w�?�            pq@Y       \                    @�"D�O[�?z            @g@Z       [                    �?�Мk#�?t            �e@������������������������       �|>�+78�?0            �Q@������������������������       �� �f���?D            �Y@������������������������       ��]�`��?             *@^       a                    �?^��o2��?8            @W@_       `                   �4@�e����?            �B@������������������������       �~VC�1��?             5@������������������������       �     ��?	             0@b       c                    @Y�Cc�?"             L@������������������������       �,�Œ_,�?             >@������������������������       ���1G���?             :@e       j                    @iQjG�?h            �d@f       i                    @�&%�ݒ�?C            @Z@g       h                    @��8��x�?=             X@������������������������       ��.y0���?              J@������������������������       � 9�����?             F@������������������������       ���E���?             "@k       l                    �?�SF�\c�?%             O@������������������������       ��E��ӭ�?
             2@m       n                    @�#��Z=�?             F@������������������������       ���.sxQ�?             ;@������������������������       ��ѳ�w�?	             1@�t�bh�h4h7K ��h9��R�(KKoKK��h��B�A       0~@      T@     �u@     �@@     @T@      =@     �T@     ؀@     ��@     @P@     �R@     `e@     h�@     �y@      (@      J@      P@     `a@     �I@     �u@     �I@     �l@      3@     �J@      @     �K@     �{@     �|@     �I@      K@      _@     �y@     @o@      @      B@     �B@     �W@     �@@      f@      5@     @X@      @      0@              2@     �n@      p@      ,@      6@     �E@     @g@      Z@              $@      @      C@      "@      ]@      *@     �I@       @      *@              1@     �X@     @b@      "@      1@      @@      Y@     @P@              $@      @     �@@       @     @P@      @      A@               @              &@      G@     �K@       @      .@      *@     �P@      @@              "@      @      1@       @     �K@      @      >@              @              &@      =@     �D@      �?      $@      $@     �I@      =@              "@      @      &@      @      A@       @      .@              @               @      2@      :@      �?      @      @      7@      0@                              "@      @      5@      @      .@               @              @      &@      .@              @      @      <@      *@              "@      @       @       @      $@       @      @               @                      1@      ,@      �?      @      @      0@      @                              @      @      @       @      @                                       @      @              �?              ,@      �?                              @       @      @              �?               @                      "@      &@      �?      @      @       @       @                               @      �?     �I@      @      1@       @      @              @      J@     �V@      @       @      3@     �@@     �@@              �?              0@              D@      @      .@       @       @              @     �C@     �T@      @       @      .@      5@      7@              �?              .@              .@               @       @                       @      ?@      I@               @      @      @      @                              @              9@      @      *@               @              @       @      @@      @              "@      ,@      0@              �?              &@              &@      �?       @              @                      *@      "@      �?              @      (@      $@                              �?              &@      �?       @                                      *@      "@                      @      $@      @                              �?                                              @                                      �?                       @      @                                             �N@       @      G@       @      @              �?     `b@     �[@      @      @      &@     �U@     �C@                              @      �?      H@       @     �D@       @      @              �?      a@      [@      @      @      &@      T@      C@                              @              @                                                      A@      &@                              @                                                       @                                                      <@      @                              @                                                      @                                                      @      @                              �?                                                     �D@       @     �D@       @      @              �?     �Y@     @X@      @      @      &@     �R@      C@                              @              >@       @      ?@       @       @              �?     �K@     �Q@      @       @      $@     �K@      ?@                               @              &@      @      $@              �?                      H@      :@       @      @      �?      4@      @                               @              *@              @                                      $@       @                              @      �?                              �?      �?      "@                                                      @      �?                              �?                                                      @              @                                      @      �?                              @      �?                              �?      �?       @              @                                                                              @      �?                                               @              �?                                      @      �?                               @                                      �?      �?     �e@      >@     �`@      .@     �B@      @     �B@     �h@     `i@     �B@      @@     @T@     �l@     @b@      @      :@      @@     �L@      8@      V@      @     �F@      @      @               @     �a@      ^@      @       @      =@     �W@      I@              (@       @      2@       @      3@      �?      3@      �?       @              @      6@      ?@               @      3@     �B@      2@              @              @      @      @      �?      .@      �?                       @      $@      .@               @      @      9@      @                              @      �?      @      �?      �?                               @      @      (@               @      @      2@      @                              �?              @              ,@      �?                              @      @                              @      @                               @      �?      *@              @               @              �?      (@      0@                      ,@      (@      &@              @              @      @       @                                              �?      �?       @                      $@      @      @              @                      @      @              @               @                      &@       @                      @      @      @                              @       @     @Q@      @      :@       @      @              @     �]@     @V@      @      @      $@      M@      @@               @       @      &@       @     �E@              5@       @      �?              @     �Y@      S@      @      @      @      H@      3@               @      �?      @       @      "@               @                                      A@     �A@              @      @      $@      @                                      �?      A@              3@       @      �?              @     @Q@     �D@      @       @      @      C@      *@               @      �?      @      �?      :@      @      @              @              �?      0@      *@                      @      $@      *@              @      �?       @              3@      �?      @              �?                      (@      @                              @      @              @      �?      �?              @      @       @              @              �?      @      "@                      @      @      $@              @              @             �U@      9@     @V@      (@      >@      @      =@      L@     �T@     �@@      8@      J@     �`@      X@      @      ,@      >@     �C@      0@     @Q@      4@     @Q@      @      .@      @      2@      L@     �Q@      5@      2@      A@     �]@      S@       @      $@       @     �@@       @     �C@      &@      ;@      �?      "@               @      *@      2@      $@      *@      .@     �E@      E@       @      @      @      1@      @      =@      $@      1@      �?      @              @      (@      (@      @      @      "@      8@      9@       @      �?      @      @      @      $@      �?      $@              @              @      �?      @      @      "@      @      3@      1@              @              &@      @      >@      "@      E@      @      @      @      $@     �E@     �J@      &@      @      3@      S@      A@              @      @      0@      �?      $@              5@      @              @      @      *@      "@      �?       @      "@      :@      &@               @              "@              4@      "@      5@      @      @      �?      @      >@      F@      $@      @      $@      I@      7@              @      @      @      �?      1@      @      4@      @      .@       @      &@              (@      (@      @      2@      .@      4@      �?      @      6@      @       @      1@      @      *@      @      .@       @      &@              &@       @      @       @      .@      3@      �?      @      4@      @      @      .@      @      (@      @      *@       @      &@              $@       @      @      @      *@      2@      �?      @      (@      @      @       @              �?               @                              �?                      �?       @      �?                       @                               @      @      �?                                      �?      @              $@              �?              �?       @      �?      @                       @      �?                                      �?      �?               @                              �?       @              @               @      @                                                      @               @              �?                              �?             �`@      =@     @]@      ,@      <@      7@      <@     @X@     �b@      ,@      5@     �G@     �e@     @d@      "@      0@      ;@      F@      2@     �Q@      3@     �T@      "@      7@      4@      (@      F@     �S@      *@      3@      B@     �V@      Y@      @      (@      :@      ;@      ,@      ;@      @      7@      @       @      @      @      A@      F@      �?      @      &@      E@     �C@      �?      @      *@      "@      @      3@      @      @              @                      @      &@      �?                      $@      ,@      �?       @              @      �?      *@              �?              @                      @      @      �?                      @      *@      �?      �?              @      �?      @                              @                      @      @      �?                      @      $@              �?              @      �?      @              �?                                                                               @      @      �?                                      @      @      @                                              @                              @      �?              �?                               @       @      1@      @      @      @      @      <@     �@@              @      &@      @@      9@              @      *@      @      @       @              "@                              �?      8@      1@               @      @      4@      @              �?              @      �?                       @                              �?      1@      @                      �?      (@       @                                      �?       @              @                                      @      &@               @      @       @       @              �?              @              @       @       @      @      @      @      @      @      0@              �?      @      (@      5@              @      *@       @       @                      @                      �?      �?              @                       @      @      @              �?      �?       @      �?      @       @       @      @      @       @      @      @      $@              �?      @      @      2@               @      (@              �?     �E@      ,@      N@      @      .@      1@      @      $@     �A@      (@      0@      9@      H@     �N@      @      @      *@      2@      $@      @                                                       @                                      @                                                      B@      ,@      N@      @      .@      1@      @       @     �A@      (@      0@      9@     �F@     �N@      @      @      *@      2@      $@      7@       @      1@              @              �?      @      (@      @      @      @      0@      3@              @      @      @      @      .@       @      (@              @              �?      @      (@      @      @      @      "@      @              �?      @       @      @       @              @               @                      @              �?              �?      @      *@               @      �?       @              *@      (@     �E@      @      $@      1@      @       @      7@      @      (@      4@      =@      E@      @      @      @      ,@      @      @      @      "@      @      "@      *@              �?      1@      @      @       @      (@      "@      @      �?       @      "@       @       @      @      A@      @      �?      @      @      �?      @      @       @      (@      1@     �@@      �?       @      @      @      @      O@      $@      A@      @      @      @      0@     �J@     @Q@      �?       @      &@      U@      O@      @      @      �?      1@      @      G@      @      5@       @      �?       @      @     �C@      G@      �?      �?      @     �O@      8@               @              *@      �?     �A@       @      0@       @      �?              @      >@      B@      �?      �?      @     �@@      *@               @              @             �A@       @      0@       @      �?              �?      >@      ?@              �?      @      @@      &@               @              @              .@              (@                              �?       @      $@              �?      @      (@      @              �?                              4@       @      @       @      �?                      6@      5@                       @      4@      @              �?              @                                                              @              @      �?                      �?       @                                              &@       @      @                       @       @      "@      $@                              >@      &@                              $@      �?      @       @                               @              @      @                              @      @                              @      �?       @                                       @              @       @                              @      @                                      �?      �?       @                                                      @                              @       @                              @               @              @                               @      @      @                              8@      @                              @              @              @                                       @      @                              &@      �?                              @              @                                               @      �?                                      *@      @                               @              0@      @      *@      @      @      �?      "@      ,@      7@              �?      @      5@      C@      @       @      �?      @      @      0@      �?      "@      @      �?               @      (@      1@              �?      @      @      :@               @              @      @      &@      �?      @      @      �?               @      (@      1@              �?      @      @      9@              �?              @      @      &@              @      @      �?                      @      "@              �?      �?      @      &@              �?              @       @              �?      @                               @      "@       @                       @       @      ,@                              �?      �?      @               @                                                                                      �?              �?                                      @      @              @      �?      @       @      @                       @      0@      (@      @              �?                              @      �?                                       @      @                              @      @                                                       @      @              @      �?      @              @                       @      (@      @      @              �?                              �?                      �?      �?      @              @                       @      (@       @      �?              �?                              �?      @               @              @                                                      @       @                                �t�bub��#     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�)*hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmK{hnh4h7K ��h9��R�(KK{��hu�B�         >                   �3@�ˣ͂��?�	           ��@       !                     @��y�2��?�           8�@                          �1@��6ndC�?r           ��@                           �?;�J�i�?            {@                          �0@�8��8��??             X@                           �?w��o	�?             =@������������������������       �3�R�f�?             3@������������������������       �R���Q�?             $@	       
                    �?�d� ��?0            �P@������������������������       ��9+�Q�?             =@������������������������       �窷uJ��?             C@                           @R@x���?�             u@                           @�)H�?�            Pq@������������������������       �������?�            @l@������������������������       �AZs����?$            �I@                          �0@��D�E��?+            �N@������������������������       ���[��"�?             2@������������������������       ���{�<�?            �E@                           @9�!/9��?V           h�@                            �? �sR���?�            p@                           �?d}o4O�?I            �]@������������������������       �=���D�?            �@@������������������������       ���M��?6            @U@                          �2@�&Z̉`�?W            `a@������������������������       ��Z��%,�?-            @R@������������������������       ���-��?*            �P@                           @t#�m�G�?�            �r@                            �?�N�"���?x            `g@������������������������       ��Y���?L            @]@������������������������       �`�j��?,            �Q@                             �?,�]U��?>            @\@������������������������       �AW/���?            �H@������������������������       �     |�?%             P@"       1                    @d5��\��?           �z@#       *                    @\��"e��?�             r@$       '                   �1@v�XԖ�?�            �j@%       &                   �0@��`so��?1            �R@������������������������       �VUUUUU�?             8@������������������������       �|a2U0�?#             I@(       )                    �?��i�<]�?S            @a@������������������������       ��["5��?"            �J@������������������������       �ÛtM&��?1            @U@+       .                    �?����a�?2             S@,       -                   �1@d����?             =@������������������������       �������?
             ,@������������������������       ���2Tv�?
             .@/       0                    �? ����?            �G@������������������������       �     @�?             0@������������������������       ��w�u��?             ?@2       9                    @�n?�6d�?Z            �a@3       6                    �?g	J�R��?8            �U@4       5                    @M�h���?              J@������������������������       ��$I�$I�?             <@������������������������       �r�q��?             8@7       8                   �2@:!��d�?            �A@������������������������       ��e��a��?             9@������������������������       ����Q��?             $@:       ;                    @������?"             L@������������������������       �������?	             ,@<       =                   �2@���S�r�?             E@������������������������       ����Mb�?             9@������������������������       �	6c����?             1@?       ^                    �?���o
�??           v�@@       O                   �=@F�e&d�?�           ��@A       H                    @�T-_�?�           ��@B       E                    �?��؟���?B           x�@C       D                    �?����X/�?�             l@������������������������       �x�)�J�?1            @U@������������������������       �*���o��?Z            `a@F       G                     @p�����?�            �r@������������������������       ��X��?h             f@������������������������       ��M�N��?O            �_@I       L                    @�kݴ��?_           ��@J       K                   �4@��)S��?k            `d@������������������������       �RM�ı��?             =@������������������������       �Weׇ�n�?\            �`@M       N                    �?����>�?�            @w@������������������������       �������?c            `b@������������������������       ���)k8+�?�             l@P       W                    �?���7��?[            @b@Q       T                    @/�����?             E@R       S                      @q=
ףp�?             4@������������������������       ��ˠT�?             &@������������������������       ��<ݚ�?             "@U       V                   @@@��.���?             6@������������������������       �r�q��?             (@������������������������       ��������?	             $@X       [                    @�ջ����?=             Z@Y       Z                     @�`�`�?             >@������������������������       �����H�?             2@������������������������       �UUUUUU�?             (@\       ]                   �?@@�|���?+            �R@������������������������       ��&%�ݒ�?             5@������������������������       �Bռ(���?            �J@_       n                    �?m�T�σ�?C           �@`       g                     @����-��?           �x@a       d                   �7@~�z݆�?�            `t@b       c                    �?
uI��~�?�            �k@������������������������       ���D=��?P             _@������������������������       �     0�?C             X@e       f                    �?�9O|�?A            �Z@������������������������       ��p�r�m�?            �H@������������������������       �������?&            �L@h       k                    @�6*����?.            �Q@i       j                    �?~�O�+�?             ?@������������������������       ��������?             1@������������������������       �4և����?             ,@l       m                   �7@ƵHPS!�?            �C@������������������������       �������?             7@������������������������       �     ��?             0@o       v                   �:@����ı�?A           ��@p       s                    @ݲ�6�>�?�           �@q       r                   �7@,�uK�B�?Q            �`@������������������������       ��x��ݳ�?6            �U@������������������������       �Ũ�oS��?            �F@t       u                   �8@��$�O�?z           ��@������������������������       ��P��;�?5           �}@������������������������       ��L!��?E            @Y@w       x                    �?��	;���?v            �f@������������������������       �      �?
             4@y       z                   �<@H�z�g�?l             d@������������������������       �YsW&�?/            �Q@������������������������       �d��c��?=            @V@�t�bh�h4h7K ��h9��R�(KK{KK��h��BI       �}@      U@     �u@     �A@      U@      7@     �R@     ��@     `�@     @P@     �S@     �c@     P�@     �z@      (@     �L@      J@     �^@     @Q@     �h@      ,@     �Y@      @      @              "@     �u@     �q@      $@      4@      F@     �l@     �Y@              @      @      =@      (@      a@      $@      K@      �?                       @     �q@      k@       @      *@      @@     @b@     �L@                      @      &@       @      I@      @      4@                              @     �a@     �X@      @      @      "@      S@      "@                              @      @      .@              @                                      4@      1@      @      �?      @      7@      �?                              �?      @      @              @                                      @      "@                              @                                                      @               @                                       @       @                              @                                                      @               @                                      @      �?                              �?                                                      "@               @                                      .@       @      @      �?      @      2@      �?                              �?      @      @               @                                      @      @              �?      @      @      �?                                      @      @                                                       @      @      @              �?      ,@                                      �?       @     �A@      @      ,@                              @     �^@     @T@              @      @     �J@       @                              @              4@      @      *@                              @     @[@      Q@              @      @     �D@      @                                              1@      @      (@                              @     �W@      H@              @       @      B@      �?                                              @              �?                                      ,@      4@                       @      @      @                                              .@       @      �?                                      *@      *@                      �?      (@      �?                              @              "@                                                      @      @                               @                                                      @       @      �?                                      "@      $@                      �?      $@      �?                              @             �U@      @      A@      �?                       @      b@     �]@      @      @      7@     �Q@      H@                      @      @      @      G@      @      0@      �?                      �?     �I@      P@              @      .@      =@      4@                              @      @      8@      @      @      �?                              6@      8@               @      @      4@      @                              �?       @      @      @      @                                      @      @                      �?      @      @                              �?              1@      �?      @      �?                              1@      5@               @      @      *@      @                                       @      6@              $@                              �?      =@      D@              �?      "@      "@      ,@                              @      �?      0@              @                              �?      .@      8@              �?       @      @      @                                              @              @                                      ,@      0@                      @      @      @                              @      �?      D@      �?      2@                              �?     @W@      K@      @      @       @     �D@      <@                      @      @              6@              ,@                              �?      S@      8@      @      @      @      :@      ,@                              �?              0@              @                              �?     �B@      .@       @      @      @      5@      *@                                              @               @                                     �C@      "@      �?                      @      �?                              �?              2@      �?      @                                      1@      >@       @              @      .@      ,@                      @       @              $@      �?       @                                      @      (@                      @      "@       @                      @      �?               @               @                                      &@      2@       @               @      @      (@                       @      �?             �N@      @      H@      @      @              �?      M@     �Q@       @      @      (@     @U@      G@              @       @      2@      @     �E@      @      ;@              �?                      ;@      F@       @      @      @      P@      D@              @       @      1@      @     �B@      @      4@              �?                      7@      >@              @      @     �L@      2@              @              $@       @      9@      �?       @              �?                      .@      @                      @      &@      @                                              $@      �?       @                                       @                                       @      �?                                              .@              @              �?                      @      @                      @      "@       @                                              (@      @      (@                                       @      7@              @      �?      G@      .@              @              $@       @      &@      �?       @                                      @       @               @              "@      @              @              @              �?       @      @                                      @      .@              �?      �?     �B@      &@                              @       @      @              @                                      @      ,@       @              @      @      6@              �?       @      @      �?      �?                                                       @      (@      �?              �?      @      @              �?               @              �?                                                      �?      @      �?                       @      @                                                                                                      �?      @                      �?      @      �?              �?               @              @              @                                       @       @      �?               @       @      2@                       @      @      �?      @               @                                                      �?                              @                       @       @      �?      �?              @                                       @       @                       @       @      ,@                              @              2@              5@      @       @              �?      ?@      :@              @      @      5@      @              @              �?      �?      "@              5@      @       @                      3@      (@              @      @      (@      @                                              @              2@       @                              @      @               @      �?      &@      @                                              @              @       @                               @      �?               @      �?       @       @                                              �?              &@                                      @      @                              @      �?                                              @              @      �?       @                      (@       @              �?       @      �?                                                      @               @               @                      (@      �?                       @      �?                                                                      �?      �?                                      @              �?                                                                      "@                                              �?      (@      ,@              �?       @      "@      @              @              �?      �?      @                                              �?      @      @                                                                              �?      @                                                       @      &@              �?       @      "@      @              @              �?              �?                                                       @      @                               @      @                              �?              @                                                              @              �?       @      �?                      @                             pq@     �Q@     `n@      ?@     @T@      7@     �P@     �h@     �t@     �K@      M@     @\@     0v@     pt@      (@      I@     �F@     �W@     �L@     �^@     �@@     ``@      ,@     �I@      .@      F@      N@     @^@      =@     �G@      P@     @c@     �c@      @      >@      @@     �H@      G@     �]@      ?@      ^@      @      C@      &@     �B@      N@     �\@      2@      @@     �H@      c@     �b@       @      9@      4@      E@     �B@     �G@      3@     �J@      @      0@       @      2@     �A@     @S@      "@      "@      =@     �V@     �O@       @      $@      $@      7@      &@      >@      @      8@               @               @      2@      B@       @      @      $@     �G@      3@      �?      @      �?      @      @      @      @      ,@                              @      @      5@       @      @      �?      0@                       @                      @      8@              $@               @              @      &@      .@              �?      "@      ?@      3@      �?      @      �?      @      �?      1@      (@      =@      @      ,@       @      $@      1@     �D@      @      @      3@      F@      F@      �?      @      "@      2@      @      ,@       @      6@      @      @              @      *@      4@      @      @      @      B@      8@      �?      �?       @      @      �?      @      @      @              $@       @      @      @      5@      @      �?      (@       @      4@              @      @      (@      @     �Q@      (@     �P@      @      6@      "@      3@      9@      C@      "@      7@      4@     �N@     @U@              .@      $@      3@      :@      ?@       @      .@      @      $@       @       @      $@      *@      @      @      @      &@     �C@              @      @       @      @      @                                                      �?       @               @      �?       @      (@               @                              8@       @      .@      @      $@       @       @      "@      &@      @       @      @      "@      ;@              �?      @       @      @      D@      $@      J@      �?      (@      @      1@      .@      9@      @      3@      0@      I@      G@              (@      @      1@      5@      5@      @      (@      �?      @      @      @      "@      (@               @      @      >@      1@               @      @      @      @      3@      @      D@              "@      @      (@      @      *@      @      &@      $@      4@      =@              $@       @      ,@      0@      @       @      &@      @      *@      @      @              @      &@      .@      .@       @      &@      @      @      (@      @      "@      @              @              @              �?              @              @      �?       @      @      �?      �?       @      �?      @      @                                                              �?              @      �?              @              �?                      @      �?                                                              �?              @      �?              �?                                      @       @                                                                               @                      @              �?                              �?              @              @              �?              @                               @       @      �?               @      �?                              @              �?                              @                               @       @                              �?              �?               @              @              �?                                                              �?               @                               @      @      @      "@      @      @               @      &@      "@      ,@              @      @      @      $@      @      @                       @       @      @                                      @              �?              @      @      @      �?              �?                       @              @                                      @              �?              �?              @                                                       @                                               @                               @      @              �?              �?               @      @      @       @      @      @               @      @      "@      *@              �?              �?      "@      @      @               @      �?       @              �?      @              �?       @      �?                      �?                       @       @                              @      @       @      @                      �?      @       @      *@                              �?      @      @      @     �c@     �B@      \@      1@      >@       @      6@     @a@     �j@      :@      &@     �H@      i@      e@      @      4@      *@     �F@      &@      H@      1@      8@      �?       @      @      @     �I@     @V@       @       @      *@     �M@      J@              @              $@      @      E@      $@      6@      �?               @      @     �G@     @T@       @       @      (@     �G@     �A@              @              @       @      5@      @      *@                      �?      �?     �@@     �P@       @              $@     �B@      9@               @              @              (@      @       @                                      0@      F@       @              @      7@      $@                                              "@      �?      @                      �?      �?      1@      7@                      @      ,@      .@               @              @              5@      @      "@      �?              �?      @      ,@      ,@      @       @       @      $@      $@              @                       @      1@              @                                       @      $@      �?               @      @      @              �?                              @      @       @      �?              �?      @      (@      @      @       @              @      @               @                       @      @      @       @               @      @              @       @                      �?      (@      1@                              @      �?       @      @       @                      @               @      @                      �?      @      @                              @                      �?       @                      @               @       @                              @      @                                               @       @                                                      @                      �?              �?                              @              @      @                       @                       @      @                              "@      (@                               @      �?       @                                                       @      @                               @      (@                              �?      �?       @      @                       @                                                              @                                      �?             @[@      4@      V@      0@      <@      @      .@     �U@      _@      2@      "@      B@     �a@      ]@      @      .@      *@     �A@       @     �W@      ,@     �Q@      ,@      0@              "@     �S@     @[@      @      @      7@     �_@     �V@      @      &@       @      ;@      @      .@      �?      1@      "@                              5@      0@       @              �?      A@      $@              �?              @              ,@      �?      @      @                              1@       @      �?                      8@       @              �?              @              �?              &@      @                              @       @      �?              �?      $@       @                              �?              T@      *@      K@      @      0@              "@     �L@     @W@      @      @      6@     @W@     @T@      @      $@       @      6@      @      Q@       @      H@      @      &@              @      K@     �T@      @      @      *@      Q@     @P@      @      @       @      2@      @      (@      @      @              @               @      @      $@              �?      "@      9@      0@              @              @              ,@      @      1@       @      (@      @      @      "@      .@      (@       @      *@      .@      9@      �?      @      &@       @      @              �?       @      �?                              @              @                                                      @                      ,@      @      .@      �?      (@      @      @      @      .@      @       @      *@      .@      9@      �?      @      @       @      @      @      @       @      �?      �?      �?      @      @      $@      @       @       @      @      (@                      @      @      @      "@       @      *@              &@       @       @      �?      @      �?              &@       @      *@      �?      @              @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�&:hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         >                   �2@��绖�?�	           ��@       !                     @��y�h�?�           H�@                           �?�o�>Ɩ�?�           ��@                            �?_�g���?s             f@                           @�~	c���??            @X@                          �1@��2(&�?             F@������������������������       ��b�=y�?             9@������������������������       ��	"P7��?             3@	       
                    �?����m�?#            �J@������������������������       �     @�?	             0@������������������������       �A-�_ .�?            �B@                           �?n)��b�?4            �S@                           �?j]���~�?            �A@������������������������       �36�v[�?             7@������������������������       �9��8���?             (@                           �?���!pc�?             F@������������������������       �� =[y�?             1@������������������������       ��s��g�?             ;@                            �?
����?[            �@                           @�z0�?�            �i@                           @� ���?M             _@������������������������       �e������?-             R@������������������������       �3�E��?              J@                           @�`غ��?3            �T@������������������������       ����Dl�?            �I@������������������������       �     ��?             @@                          �0@�7L�?�            Pu@                           �?�y�}�)�?3            �Q@������������������������       �4���C�?            �@@������������������������       �x�"w���?             C@                            �?�Gm=��?�            �p@������������������������       �Bf����?e            @e@������������������������       ���v���?C             Y@"       1                   �1@�e!}�?�            �s@#       *                    �?/V"H��?m            �e@$       '                    @,R�n��?0             R@%       &                    �?N��)x9�?             <@������������������������       ��zv��?             &@������������������������       �$�ɜoB�?
             1@(       )                    �?}��7�?             F@������������������������       ��z�G��?             4@������������������������       �UUUUUU�?             8@+       .                    @�g��s��?=             Y@,       -                    @���:��?            �A@������������������������       �     @�?	             0@������������������������       �0\�Uo��?
             3@/       0                    �?R;�Uz��?*            @P@������������������������       ���IF�E�?            �@@������������������������       �     ��?             @@2       9                    @��G;��?\            @b@3       6                    @�W'�]��?A            �X@4       5                    �?r�q��?              H@������������������������       �����X�?             5@������������������������       �A��?�?             ;@7       8                    @��Q���?!             I@������������������������       ��\�l8b�?            �A@������������������������       �N贁N�?             .@:       ;                    �?��8��8�?             H@������������������������       ��)x9/�?             ,@<       =                    �?2�^��"�?             A@������������������������       �$����%�?
             3@������������������������       �؂-؂-�?             .@?       X                    �?"��@��?           n�@@       O                   �?@�Y��&J�?G           ��@A       H                    �?�����?           t�@B       E                   �7@�衖���?C           0�@C       D                     �?#JS��%�?�            @s@������������������������       �6���y��?j            `d@������������������������       �t�4���?W             b@F       G                     �?������?�            @j@������������������������       �D�>��?A            �Y@������������������������       ���1�/8�?A             [@I       L                    @H V�?�           ��@J       K                    �?/���?%           �{@������������������������       �[�n�[�?q             e@������������������������       ����oH�?�            `q@M       N                    �?Ǐ�J�x�?�            �q@������������������������       ��+&�B�?>            �X@������������������������       �%�\quQ�?o            �f@P       W                    @�K9iI�?2            @S@Q       T                   �@@     (�?*             P@R       S                    �?G���t��?            �A@������������������������       �������?             ,@������������������������       �W�7�L�?             5@U       V                     @8^s]e�?             =@������������������������       ��X�%��?             .@������������������������       �I�$I�$�?	             ,@������������������������       �؉�؉��?             *@Y       h                   �9@`3^�i�?�           4�@Z       a                   �7@(�Zߦ��?           t�@[       ^                     �?IfT���?�           $�@\       ]                    @ζ����?}           0�@������������������������       �K�V��w�?           p{@������������������������       �֝~�0�?p            �e@_       `                    @��u���?           0z@������������������������       ��ŪU{~�?�            �s@������������������������       �k+��ݓ�?B             Y@b       e                    @7V>��;�?�            �j@c       d                     �?�;m��?_            �c@������������������������       �\F���?            �D@������������������������       �h��'��?E            �\@f       g                    �?n۶m۶�?$             L@������������������������       �L$e?���?             7@������������������������       �3(&ޏ�?            �@@i       p                    �?��h�*$�?�             s@j       m                     �?�G���?N            �\@k       l                    @-�܃QN�?             ?@������������������������       �h���eP�?             6@������������������������       ���"e���?             "@n       o                   �=@�w��&��?9            �T@������������������������       ��A����?(            �L@������������������������       ���?��?             :@q       t                    �?v!�?}            �g@r       s                    @)^���?*            @P@������������������������       ��9(!�;�?            �C@������������������������       �.�T�6�?             :@u       v                    @o���?S            @_@������������������������       ��):���?B             Y@������������������������       �9��v���?             9@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F        }@     �V@     �s@      E@     �R@      <@     @U@     H�@     H�@     �Q@     �V@      b@     ��@      {@      $@     �J@      J@     �`@     �K@     �b@      @     @R@      �?      @              &@     0r@      k@       @      @      .@     `c@     �Q@              @              9@      @     �U@       @      A@              �?               @     �l@     �d@      @       @      (@     �[@      H@               @              *@      �?      <@      �?      0@              �?              �?      B@     �A@      �?      �?      $@      @@      "@                              @      �?      .@      �?      "@                                      6@      (@              �?      @      5@       @                              @              @              @                                      .@      @              �?      �?      @      @                              @               @              @                                      $@      @              �?              @      �?                                              @                                                      @                              �?      @      @                              @              $@      �?      @                                      @       @                      @      .@      @                                                              @                                              �?                       @      "@                                                      $@      �?      �?                                      @      @                       @      @      @                                              *@              @              �?              �?      ,@      7@      �?              @      &@      �?                              �?      �?      $@                                              �?      @       @      �?              @      @                                                      @                                                      @      @                      @      �?                                                      @                                              �?              @      �?              �?       @                                                      @              @              �?                      @      .@                               @      �?                              �?      �?                                                              @      @                              @      �?                                      �?      @              @              �?                       @      $@                              @                                      �?             �M@      �?      2@                              @     `h@     �`@      @      �?       @     �S@     �C@               @              "@              :@      �?       @                               @      L@      P@       @              �?      A@      ,@                              @              3@      �?       @                              �?      E@      <@                              9@      @                              �?              &@               @                                      1@      3@                              4@      @                                               @      �?                                      �?      9@      "@                              @       @                              �?              @                                              �?      ,@      B@       @              �?      "@      "@                              @              �?                                              �?      @      =@       @              �?      @       @                               @              @                                                      $@      @                              @      �?                               @             �@@              0@                              @     `a@      Q@       @      �?      �?     �F@      9@               @              @              @               @                                      C@      $@                              $@      �?                              @              @               @                                      7@       @                               @                                                      @                                                      .@       @                               @      �?                              @              :@              ,@                              @     @Y@      M@       @      �?      �?     �A@      8@               @              �?              (@              @                               @     @S@      D@                              5@      &@                                              ,@              @                              @      8@      2@       @      �?      �?      ,@      *@               @              �?             �O@      @     �C@      �?       @              @      N@      I@      @      @      @      F@      6@              @              (@       @     �C@              *@               @                     �B@     �A@      @      @       @      4@      ,@               @               @              5@              @              �?                      ,@      @      @       @       @      @       @              �?              �?              &@                              �?                       @      �?      @       @      �?      @      @                                               @                                                       @              @              �?      @                                                      "@                              �?                              �?               @              �?      @                                              $@              @                                      (@      @                      �?       @      @              �?              �?              @               @                                       @      @                                      �?                                              @              @                                      @       @                      �?       @      @              �?              �?              2@              @              �?                      7@      =@              �?              ,@      @              �?              �?               @              �?                                      @      (@                              @       @                              �?              @              �?                                      @       @                              @                                                      @                                                              $@                               @       @                              �?              $@              @              �?                      3@      1@              �?              @      @              �?                              @              @                                      (@      @                              @                                                      @               @              �?                      @      &@              �?               @      @              �?                              8@      @      :@      �?                      @      7@      .@               @      �?      8@       @               @              $@       @      3@      @      $@      �?                      �?      &@      ,@               @      �?      1@      @               @              "@              (@      @      "@                              �?       @      @              �?              $@       @                              @              @      �?      @                              �?      �?                                      @      �?                              @              @      @      @                                      �?      @              �?              @      �?                                              @      �?      �?      �?                              "@      &@              �?      �?      @      @               @              @              @      �?              �?                              @      "@                      �?      @      @                              �?              �?              �?                                       @       @              �?              �?      �?               @              @              @              0@                               @      (@      �?                              @       @                              �?       @      @              @                                      @                                               @                                               @              &@                               @       @      �?                              @                                      �?       @                      &@                               @       @                                      @                                                       @                                                      @      �?                              @                                      �?       @     �s@      U@     @n@     �D@      R@      <@     �R@     `p@      y@      O@     �T@     @`@     �{@     �v@      $@     �G@      J@     �[@      J@      a@      H@     �`@      8@      G@      5@      A@     �J@     �`@      =@      M@      O@     �h@      f@      @      ?@     �A@      P@     �C@     �`@      H@     @_@      2@     �A@      0@     �@@     �J@     �`@      9@      J@      J@     �h@     �e@      �?      =@      =@      N@      A@     �L@      &@      K@      @      *@      @      *@      <@     @S@      @      5@      0@     �X@     �P@      �?      $@       @      2@      (@      B@      �?     �C@      @      $@      @      @      8@      C@      @      &@      &@     �Q@      A@      �?      @      �?      $@      @      9@      �?      .@              @              @      ,@      1@      �?      @      @      I@      0@               @              @              &@              8@      @      @      @              $@      5@      @      @      @      4@      2@      �?      �?      �?      @      @      5@      $@      .@      @      @              $@      @     �C@              $@      @      <@      @@              @      @       @      @      @      @      @      �?                      @      @      7@               @       @      @      5@                      @      @      @      ,@      @       @      @      @              @              0@               @      @      8@      &@              @      @      �?      �?      S@     �B@     �Q@      &@      6@      (@      4@      9@     �K@      5@      ?@      B@     �X@      [@              3@      5@      E@      6@      K@      5@     �E@      @      1@      "@       @      2@     �E@      (@      &@      1@     �Q@      P@              &@      *@      4@      $@      :@      @      3@       @      &@      �?      @      @      *@      �?      �?       @      A@      8@              @      @      @      @      <@      0@      8@      @      @       @       @      (@      >@      &@      $@      .@     �B@      D@              @       @      .@      @      6@      0@      <@      @      @      @      (@      @      (@      "@      4@      3@      ;@      F@               @       @      6@      (@      $@       @      "@               @              @               @      @      @       @      &@      (@                      @      "@       @      (@      ,@      3@      @      @      @      @      @      @      @      .@      &@      0@      @@               @      @      *@      @      @              @      @      &@      @      �?                      @      @      $@               @      @       @      @      @      @      @              @      @      @      �?                              @      @      $@               @      @       @      @      @      @       @              �?      @      @      �?                              @      @      @               @              �?      @      @      �?      �?                              @                                      �?       @      @                                              �?              �?              �?      @              �?                              @       @                       @              �?      @       @      �?      �?              @      �?      �?                                               @      @                      @      �?       @      �?      @      �?              @      �?                                                      �?      @                              �?      �?      �?                               @              �?                                              �?      �?                      @              �?              @                      �?       @      @      @      �?                                                                                              �?     �f@      B@     �[@      1@      :@      @      D@      j@     �p@     �@@      9@      Q@     �n@     �g@      @      0@      1@      G@      *@      d@      6@     �U@      ,@      0@      @      A@      h@     �m@      0@      5@     �H@     �i@     �`@      @       @      "@      8@      @     @a@      ,@      R@       @      ,@      @      7@      f@     �g@      *@      (@      E@     `f@     �Z@              @      "@      5@      @     �R@      @      G@      @      @       @      0@     �W@     �`@      *@      $@      9@     �W@     @P@              @      @       @      @     �J@      @      6@      @      �?       @      ,@      Q@      [@      *@       @      0@      R@      E@              �?      @      @      @      6@      �?      8@       @      @               @      ;@      ;@               @      "@      7@      7@               @       @       @      �?     �O@      $@      :@      @      @      �?      @     @T@     �K@               @      1@      U@     �D@              @      @      *@       @      G@      "@      2@      @      @      �?      @      R@      C@               @      .@      P@      :@                      @      $@      �?      1@      �?       @              @              �?      "@      1@                       @      4@      .@              @              @      �?      7@       @      .@      @       @              &@      1@     �H@      @      "@      @      :@      <@      @       @              @              0@      @      &@      @                      "@      $@      E@      �?       @      @      5@      2@              �?                              �?       @      @                              @              @      �?      @              $@      $@                                              .@      @      @      @                      @      $@     �B@              @      @      &@       @              �?                              @      �?      @               @               @      @      @       @      �?      �?      @      $@      @      �?              @               @              �?                                      @      @       @      �?      �?              @              �?              �?              @      �?      @               @               @       @      @                              @      @      @                       @              3@      ,@      7@      @      $@      @      @      0@      =@      1@      @      3@     �D@      K@      �?       @       @      6@      @      (@      @      @      �?      @                      &@      2@      �?       @      @      7@      3@              @               @       @      @      �?       @                                      �?      @                       @       @      $@              �?               @              @      �?       @                                      �?      @                      �?              @              �?               @              @                                                                                      �?       @      @                                              @      @       @      �?      @                      $@      ,@      �?       @      �?      5@      "@              @                       @      @      @      �?      �?      @                      $@      (@              �?      �?      $@      @               @                      �?       @              �?               @                               @      �?      �?              &@      @               @                      �?      @       @      3@       @      @      @      @      @      &@      0@       @      0@      2@     �A@      �?      @       @      4@      @      �?      @      @       @       @      �?              �?      @      &@       @      @      "@       @               @      @      @      �?      �?      @       @      �?       @      �?                      @      @       @       @      "@      @                      �?      �?                      �?       @      �?                              �?      �?      @              �?              @               @      @      @      �?      @      @      .@              @      @      @      @      @      @              *@      "@      ;@      �?      �?      @      0@      @      @      @       @                      @      @      @      @       @              *@       @      6@      �?      �?      @      *@      @      �?              @              @                      �?      �?      @                      �?      @                              @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJa�ahG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKohnh4h7K ��h9��R�(KKo��hu�BH         4                    �?a��ni��?�	           ��@                          �4@^�'L9�?�           ܘ@                            @Q�GD,9�?�           X�@                           @d�~���?�            pv@                          �1@Y�ӗ�?�            �u@                           @6�:�e��?:            @X@������������������������       ��p=
ף�?&             N@������������������������       ���I!��?            �B@	       
                    @l&����?�            `o@������������������������       ��D��u�?N            �`@������������������������       �ϩ�=!�?G            �]@������������������������       ���ˠ�?             &@                          �0@$'z ��?�            @p@                           �? )O��?             2@������������������������       �      �?              @������������������������       �
ףp=
�?             $@                           �?���%��?�            @n@                           @���q�?8            �S@������������������������       ��q�%��?#            �I@������������������������       ��)x9/�?             <@                           �?�f�:���?e            `d@������������������������       �?�ܵ��?             I@������������������������       �J����V�?F            @\@       '                    �?�~�m�?u           `�@                             @�1��?�            �u@                          �5@#AM�h��?             j@                           �?     `�?             @@������������������������       �l�l��?	             .@������������������������       �U��6���?
             1@                            �?�zv��?l             f@������������������������       ��cQ�pf�?\            �b@������������������������       ���<,��?             9@!       $                    �?|�k\+�?U             a@"       #                    �?������?             B@������������������������       �/�s��?             3@������������������������       ��ѳ�w�?
             1@%       &                    �?�3��*�?>            @Y@������������������������       ����,d!�?             G@������������������������       �nh�)r��?#            �K@(       /                   �=@D�k#{�?�           ��@)       ,                   �8@�2*�?`           ��@*       +                     �?��y_�?�            Pt@������������������������       �M@�/��?i            @d@������������������������       ���]���?l            `d@-       .                     �?�J�x��?�            �i@������������������������       ���P�k�?4            �T@������������������������       ���.|��?W            �^@0       1                    @���T��?A            �X@������������������������       ���a_j�?             3@2       3                     �?���}B��?6            �S@������������������������       ���N��N�?             :@������������������������       ��q�MU�?&            �J@5       R                   �3@=�NUp��?�           $�@6       E                     @^��z�?X           H�@7       >                   �0@��6����?�           x�@8       ;                    �?�Y�}��?S            ``@9       :                     �?:�RHm�?1            @S@������������������������       �$߼�x�?$             N@������������������������       �V��6���?             1@<       =                     �?j"�=��?"             K@������������������������       ��iQT�?            �E@������������������������       ����k���?             &@?       B                     �?
�j^q�?�           `�@@       A                    @�_�����?           �|@������������������������       �:|z3��?�             u@������������������������       ���gE#�?C             ^@C       D                    @s����b�?t            �h@������������������������       ���Q�%�?a             d@������������������������       �h/�����?             B@F       M                   �2@�0�=��?y            @g@G       J                    �?�~�#��?X            �`@H       I                    @�Ĝ��?'             M@������������������������       ������?             ?@������������������������       ��dIG���?             ;@K       L                    �?�T�x?r�?1            @S@������������������������       ��H���?             ?@������������������������       �vLB�?�?             G@N       O                    @�W�g��?!            �I@������������������������       �b���i��?             &@P       Q                    @��Q��?             D@������������������������       ��q-�?             *@������������������������       ���k���?             ;@S       b                    �?Yz)�"��?W           $�@T       [                     �?������?           {@U       X                   �5@'���6�?�            `m@V       W                    �?��n2���?9            �X@������������������������       �M=ֱ߹�?             �L@������������������������       �R����d�?            �D@Y       Z                    �?�'+dP��?X             a@������������������������       �fffff��?3             T@������������������������       �|�%~oI�?%            �L@\       _                    �?+���H �?}            �h@]       ^                     @�K����?>            �Y@������������������������       ��X�C�?#             L@������������������������       �~K$e?��?             G@`       a                   �:@�8��8��??             X@������������������������       �����H�?1             R@������������������������       ��������?             8@c       h                   �8@����ܾ�?I           ��@d       g                    @wi���2�?}           �@e       f                    �?��T��?r           ��@������������������������       � �s-��?�            �o@������������������������       ��o�5��?�            @u@������������������������       ����S�r�?             ,@i       l                    �?u�)>�.�?�            ps@j       k                   �;@�z�G��?             >@������������������������       ����Q��?             $@������������������������       ���Q���?	             4@m       n                    @��4b��?�            �q@������������������������       ���#�a �?�            @l@������������������������       �}Vb��N�?#            �K@�t�bh�h4h7K ��h9��R�(KKoKK��h��B�A        {@     @V@     �u@      9@     �W@      <@     �T@     @�@     p�@     @R@      W@     �d@     P�@     z@      *@     �P@      G@     @`@      J@     �c@      D@     �d@      $@     �M@      4@      B@      _@      g@     �A@      K@      X@      k@     �i@      @      F@     �@@     �P@      C@     �Q@      @      M@      �?      @               @     �V@     �Z@       @      1@      B@     �Z@      L@              *@      @     �@@      @     �D@       @     �@@      �?      �?               @      M@     @R@      @       @      :@     @P@      6@              @              $@      @      D@       @     �@@      �?                       @     �L@     @R@      @       @      :@     @P@      0@              @              $@      @      $@              @                                      <@      4@      @              @      4@       @                                              @              @                                      4@      "@                      @      1@      �?                                              @              �?                                       @      &@      @              @      @      �?                                              >@       @      ;@      �?                       @      =@     �J@               @      3@     �F@      ,@              @              $@      @      (@       @      &@                              �?      *@      A@               @      @      >@      *@               @              @       @      2@              0@      �?                      �?      0@      3@              @      *@      .@      �?              @              @       @      �?                              �?                      �?                                              @                                       @      =@      @      9@              @                      @@     �@@      @      "@      $@      E@      A@              @      @      7@      �?      @               @                                      @                                      �?       @                                               @              �?                                      @                                              �?                                              @              �?                                      @                                      �?      �?                                              7@      @      7@              @                      9@     �@@      @      "@      $@     �D@      @@              @      @      7@      �?      @              @                                      .@      *@               @       @      ,@      (@              �?              "@              @                                                      (@      @              �?       @      &@      $@                              @               @              @                                      @      @              �?              @       @              �?              @              0@      @      3@              @                      $@      4@      @      @       @      ;@      4@              @      @      ,@      �?      @       @       @              @                      @      @              @              @      @               @               @              &@      �?      &@                                      @      *@      @      �?       @      6@      1@              @      @      (@      �?      V@     �A@     �Z@      "@      K@      4@      A@      A@     �S@      ;@     �B@      N@     �[@     �b@      @      ?@      <@     �@@      ?@      I@      $@      @@       @      .@       @       @      "@     �A@      0@      ,@      *@      E@      K@       @      *@      @      "@      "@      C@      @      6@      �?      @               @      @      7@       @      (@      $@      >@      =@              @      @      "@      �?      *@               @                              �?              @               @       @       @                                      @              @              �?                              �?              @                               @                                      �?              @              �?                                              @               @       @                                               @              9@      @      4@      �?      @              @      @      0@       @      $@       @      <@      =@              @      @      @      �?      2@      @      2@      �?      @              @      @      (@      @      "@      @      ;@      <@               @      @      @      �?      @               @                                              @       @      �?      @      �?      �?              @                              (@      @      $@      �?      (@       @              @      (@       @       @      @      (@      9@       @       @      �?               @      @      �?                       @                       @      @      @       @      �?       @      "@               @                       @      @      �?                                              �?      @      @       @      �?       @      @                                                                               @                      �?      �?      @                              @               @                       @      "@      @      $@      �?      $@       @              @       @       @               @      $@      0@       @      @      �?              @      @       @      @                                      @      @                              @      *@              @                      @       @      @      @      �?      $@       @                      @       @               @      @      @       @       @      �?              @      C@      9@     �R@      @     �C@      (@      :@      9@      F@      &@      7@     �G@      Q@     �W@      @      2@      8@      8@      6@     �@@      4@      P@      @      ?@       @      5@      7@      C@      $@      1@     �B@     �P@      W@              .@      .@      4@      ,@      ;@       @     �E@      @      &@      @      &@      5@      :@      @      .@      5@      A@     �L@              @      @      2@      "@      ,@      @      1@               @              @      3@      $@      �?       @      @      :@      >@               @       @      "@      @      *@      @      :@      @      @      @       @       @      0@      @      @      0@       @      ;@              @      @      "@      @      @      (@      5@      �?      4@      @      $@       @      (@      @       @      0@     �@@     �A@              $@       @       @      @      �?      "@      @      �?      $@      �?      @      �?      @      �?       @       @      .@      *@              $@       @              �?      @      @      0@              $@       @      @      �?      @      @              ,@      2@      6@                      @       @      @      @      @      &@      @       @      @      @       @      @      �?      @      $@      �?       @      @      @      "@      @       @      @      �?      @              �?                              @              �?                      �?      �?      �?                              �?      @      @      @      @      @      @       @      �?      �?      @      $@      �?      �?      @       @      "@      @       @              @                              @      @              �?              @      @              �?                       @       @      @      �?      �?      @      @      @      �?       @       @              �?      �?      @      �?              @       @      @       @      @     @q@     �H@     `f@      .@     �A@       @      G@     �z@     P{@      C@      C@     �Q@     w@     �j@      @      7@      *@      P@      ,@     @[@      &@      Q@      @      @              &@     �p@     @j@      @      $@      6@     `c@      M@              @      @      *@      @     @U@      &@     �D@       @       @               @     @m@     @g@      @      @      1@     �]@      I@               @      @      "@       @      0@                                                     �J@     �D@               @      �?      0@      �?                              �?              @                                                      B@      7@               @              "@                                                      @                                                      7@      5@               @              @                                                                                                              *@       @                               @                                                      "@                                                      1@      2@                      �?      @      �?                              �?              @                                                      $@      2@                      �?      @      �?                              �?               @                                                      @                                       @                                                     @Q@      &@     �D@       @       @               @     �f@      b@      @       @      0@     �Y@     �H@               @      @       @       @     �L@      "@      8@       @                      @     �]@     �W@       @       @      .@     �R@     �@@               @      @       @       @      F@      �?      *@       @                      @     @Z@      Q@      �?       @      &@      L@      5@              �?      @       @       @      *@       @      &@                               @      ,@      :@      �?              @      3@      (@              �?      @      @              (@       @      1@               @               @      O@     �I@      @              �?      <@      0@                                              $@       @      *@               @               @      M@      A@      @              �?      7@      (@                                               @              @                                      @      1@                              @      @                                              8@              ;@      @      @              @      B@      8@              @      @      B@       @              @              @      �?      3@              6@              @              �?      @@      (@              @      @      :@      @               @              @      �?      @              5@                              �?       @      @               @      �?      *@      �?                                              @              @                                      @      @               @      �?      @      �?                                                              .@                              �?      @       @                              @                                                      *@              �?              @                      8@      @              �?      @      *@      @               @              @      �?       @                                                      .@      �?                              @      �?                                              @              �?              @                      "@      @              �?      @      @      @               @              @      �?      @              @      @       @               @      @      (@              @      �?      $@       @               @                              �?                               @                       @                              �?      @                                                      @              @      @                       @       @      (@              @              @       @               @                                                      @                              �?      @                               @                                                      @              @                               @      �?      @              @              @       @               @                             �d@      C@     �[@      $@      <@       @     �A@     �c@     `l@     �@@      <@     �H@     �j@     `c@      @      1@      @     �I@      &@      J@      3@      8@       @      @      @      @      K@     @X@      @      (@      0@     �P@     �M@               @              @       @      6@              1@              �?              @     �B@     �L@      @      @      &@     �A@      C@               @              �?               @               @              �?              �?      8@      0@               @       @      .@      5@                                              @               @                                      1@       @              �?      @      ,@      @                                              @                              �?              �?      @       @              �?      @      �?      ,@                                              ,@              .@                               @      *@     �D@      @      @      @      4@      1@               @              �?              "@              "@                                      @     �A@      �?       @      �?      *@      @                                              @              @                               @      $@      @      @      @       @      @      $@               @              �?              >@      3@      @       @      @      @              1@      D@      �?      @      @      ?@      5@              @              @       @      2@      @       @               @      �?               @      :@               @      @      2@      ,@              �?              �?              *@      @       @                                      @      0@               @       @      "@      @              �?                              @      @                       @      �?              @      $@                      �?      "@      &@                              �?              (@      *@      @       @      @       @              "@      ,@      �?      @       @      *@      @              @              @       @      $@      @      @      �?      @      �?              "@      *@      �?                      *@      @              @              �?               @       @              �?              �?                      �?              @       @               @                               @       @     �\@      3@     �U@       @      6@      @      @@      Z@     @`@      <@      0@     �@@     �b@      X@      @      "@      @      G@      "@     �V@      $@      I@      @      &@              7@     �T@      [@      &@      (@      0@     @Y@      K@      @      @      @      5@      @     �V@      $@      H@       @      $@              6@     �T@      [@       @      (@      0@     �X@     �J@      @      @      @      5@      @      ;@      �?      1@                              @     �L@      O@               @      @     �F@      :@              �?               @      �?     �O@      "@      ?@       @      $@              2@      :@      G@       @      $@      (@     �J@      ;@      @       @      @      *@       @                       @      @      �?              �?                      @                      @      �?                                              9@      "@     �B@      @      &@      @      "@      5@      6@      1@      @      1@     �G@      E@      �?      @      @      9@      @              @      "@               @                       @       @      @                      @      �?                      @                                      @                                      �?      �?                              �?                                                              @       @               @                      �?      �?      @                       @      �?                      @                      9@      @      <@      @      "@      @      "@      3@      4@      *@      @      1@      F@     �D@      �?      @      �?      9@      @      2@      @      5@      @      @      @      @      0@      3@      "@      @      1@     �C@      =@      �?      @      �?      7@      @      @      �?      @              @              @      @      �?      @                      @      (@              �?               @      @�t�bub�R"     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJtP�vhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         8                    �?R辳]��?�	           ��@                           �?_N��R,�?           �@                          �4@g$zX���?�           ��@       	                   �1@N�Q����?�            �n@                            �?�V����?(            @P@������������������������       �ףp=
��?             4@                            @�ks����?            �F@������������������������       ��l� {�?             1@������������������������       �c}h���?             <@
                            �?�6탵�?n            �f@                           �?������?             B@������������������������       ����k���?             6@������������������������       ����X�?             ,@                          �3@n&,���?U             b@������������������������       ��T��n�?8            @X@������������������������       �r�q�?             H@                          �>@*�)����?           �x@                          �7@��{`��?�            0v@                           @���1�A�?s            �d@������������������������       �$�_�0�?m            �c@������������������������       �      �?              @                          �9@�d�����?z            �g@������������������������       ��g5n�?8            �U@������������������������       ����a��?B            @Y@                          @@@�Rͦ$�?            �B@                           �?�����?             6@������������������������       ��G�z��?             $@������������������������       �r�q��?	             (@������������������������       �t�@�t�?             .@       -                   �=@�p*�W�?u           ��@       &                   �6@T.#��?9           ��@        #                   �4@�r����?E           P@!       "                     �?\mg�wo�?�             u@������������������������       ���钹H�?Z            �a@������������������������       �"���;�?�            �h@$       %                     @#Ĝ�5�?f            `d@������������������������       �����c��?7             U@������������������������       ��ϗkaY�?/            �S@'       *                   �7@�x� v�?�            pz@(       )                    @,Z�}2�?+            @Q@������������������������       ���6�80�?             C@������������������������       ��߸�ǒ�?             ?@+       ,                    @h�+���?�             v@������������������������       �����1��?�            �s@������������������������       �2���h��?             C@.       3                   �?@r�qW�?<             X@/       0                    �?)\���(�?            �A@������������������������       �*L�9��?             &@1       2                     �?�8��8��?             8@������������������������       ������H�?             "@������������������������       ��.�?�P�?
             .@4       5                     �?}R��ɞ�?$            �N@������������������������       �ƵHPS!�?             *@6       7                     �?UUUUU��?             H@������������������������       ��.�?�P�?	             .@������������������������       ����#���?            �@@9       X                   �4@���2��?�           ��@:       I                     @@��#_�?�           |�@;       B                   �0@�AZ����?L           ��@<       ?                    �?0��>���?U             a@=       >                     �?8tM���?"            �L@������������������������       �$G�h��?             7@������������������������       ��������?             A@@       A                    @�������?3            �S@������������������������       ��ۑ��?            �B@������������������������       �>��t�?             E@C       F                    @r+?�h�?�           p�@D       E                   �2@���N�?�?�           ��@������������������������       �Xf�E�?�            �y@������������������������       ��mq�v/�?�            �u@G       H                     �?�,騷}�?"             K@������������������������       �/��.���?            �B@������������������������       �*�8�G��?             1@J       Q                    @����?�             m@K       N                    @��P�B�?P            �^@L       M                    �?����?;            @V@������������������������       �3�E��?4            �S@������������������������       �2(&ޏ�?             &@O       P                   �3@X��H��?             A@������������������������       �+7����?             7@������������������������       ��C��2(�?             &@R       U                    @[nh�)r�?K            �[@S       T                    �?�z�G��?$             I@������������������������       ��^|�!�?             7@������������������������       �#����?             ;@V       W                   �2@�:m���?'             N@������������������������       ��b-�I�?             C@������������������������       �h���eP�?             6@Y       h                    �?My�r���?�           ��@Z       a                    �?�bq�Z��?�            Ps@[       ^                     @	W����?f            �d@\       ]                    @��o�	'�?V            @a@������������������������       ��y��/�?3            �S@������������������������       ��3����?#            �M@_       `                    @m��
I��?             ;@������������������������       ������H�?             "@������������������������       ��q�q�?
             2@b       e                   �8@����HY�?b             b@c       d                    @-��rҐ�?;            �U@������������������������       �&5DSb�?,             Q@������������������������       ��������?             2@f       g                   �=@io8�?'             M@������������������������       �/�����?             E@������������������������       �     ��?	             0@i       p                    @P�b����?�           ؇@j       m                   �;@�$ĺ���?�           h�@k       l                    @<KQ�^�?[           �@������������������������       ��V�W )�?�            �v@������������������������       ��ڎ&�U�?m            �f@n       o                    @�z�dC
�?H            �Z@������������������������       ��ƺ�W�?/            @R@������������������������       ��IєX�?             A@q       t                     @G^�X7��?B            �[@r       s                     �?9ǽ��2�?.            �Q@������������������������       ��uϪ~�?!            �H@������������������������       ��zv��?             6@u       v                   �7@!�����?            �C@������������������������       �K�]l���?             =@������������������������       ���Q��?             $@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       �y@      N@     Pt@     �@@     @U@      A@     �W@     �@     @�@     �L@     �Z@     �c@     X�@     �{@      &@     �L@     �O@     �a@     �N@     �g@      @@     �d@      2@      J@      ;@     �J@     @Y@      h@      ;@     �P@     �T@     `l@     �k@      @     �@@      E@     @R@     �F@     @U@      &@      K@      @      .@       @      3@     �O@     �W@      @      7@      4@      [@     �R@      @      (@      (@      6@      *@      <@      @      .@              @                     �D@     �I@      @      "@       @      G@      9@              @              &@       @      &@              @                                      4@      &@       @                      $@      @                                               @              @                                      @      �?                               @      �?                                              @              @                                      0@      $@       @                       @      @                                              �?                                                       @       @                              @      �?                                               @              @                                       @       @       @                      @       @                                              1@      @       @              @                      5@      D@       @      "@       @      B@      5@              @              &@       @      @      �?      �?                                      @      @               @      �?      0@                                              �?      @                                                              @                              ,@                                                      @      �?      �?                                      @                       @      �?       @                                              �?      $@      @      @              @                      2@      B@       @      @      �?      4@      5@              @              &@      �?      @      @      @                                      "@      7@       @      @              2@      ,@              @              &@              @               @              @                      "@      *@              @      �?       @      @              �?                      �?     �L@      @     �C@      @      &@       @      3@      6@     �E@              ,@      2@      O@      I@      @       @      (@      &@      &@      J@      @     �B@      @       @       @      *@      6@     �D@              &@      2@     �N@      E@      �?       @      $@      $@      "@     �@@      �?      3@       @      @      �?       @      *@      .@              @      @      @@      ,@      �?      @      @      @      �?      @@      �?      2@       @      @      �?       @      &@      ,@              @      @      @@      &@      �?      @      @      @      �?      �?              �?                                       @      �?                                      @                                              3@      @      2@      �?       @      �?      @      "@      :@              @      *@      =@      <@              @      @      @       @      @               @                      �?      @      @      1@                      @      &@      6@               @      @       @      �?      .@      @      $@      �?       @              �?      @      "@              @      @      2@      @               @      @      @      @      @               @              @              @               @              @              �?       @       @               @      �?       @      �?              �?              �?              @               @               @              �?       @                              �?       @                                                       @               @                              �?      @                              �?              �?              �?              �?              �?                               @                      @                                       @      @              �?               @              @                              �?                               @               @                     �Z@      5@     @\@      .@     �B@      9@      A@      C@     �X@      7@      F@      O@     �]@     �b@       @      5@      >@     �I@      @@     @Z@      4@      Z@      $@      A@      3@      @@      C@      W@      .@     �A@     �H@     �]@     `b@              0@      2@     �F@      :@     �Q@      $@     �J@      @      0@      @      ,@      ?@      Q@       @      .@      =@     �Q@     �O@               @      @      =@      @     �F@      @     �C@      @      @              @      =@     �H@      �?      "@      4@      K@     �F@              @       @      4@      @      &@              .@      @      �?              @      .@      9@               @      $@      8@      ,@                              *@      @      A@      @      8@              @                      ,@      8@      �?      @      $@      >@      ?@              @       @      @      @      9@      @      ,@              &@      @      $@       @      3@      @      @      "@      0@      2@              @      @      "@              4@      �?      @                              @       @      (@       @      @      @      "@      $@               @               @              @      @      @              &@      @      @              @      @       @      @      @       @               @      @      �?             �A@      $@     �I@      @      2@      0@      2@      @      8@      @      4@      4@     �H@      U@               @      *@      0@      4@       @      �?       @      �?      @      @      �?      �?      @       @       @      �?      @      @                      @       @      "@       @      �?      @      �?       @      @              �?      @      �?              �?      @      �?                       @      �?                               @               @              �?                      �?       @                      @                      �?      �?      "@      ;@      "@     �E@      @      ,@      &@      1@      @      4@      @      (@      3@     �F@     @S@               @      $@      ,@      &@      6@       @      >@      @      ,@      &@      0@      @      1@      @      (@      1@      E@     �R@              @      $@      &@      &@      @      �?      *@                              �?      @      @                       @      @      @              �?              @              �?      �?      "@      @      @      @       @              @       @      "@      *@              �?       @      @      (@      @      @      �?      �?      @                       @       @              @      @       @                      �?               @      @      @                      �?      @                               @                                                      �?                      @                      �?               @                       @                      @      @       @                                       @      @      @              �?                                      �?                      �?               @                                              @      �?                               @                      �?                      @      @                                               @               @                              @      @      @      @                      �?      @      @      *@                       @      @      @      @      @                       @                      @                                      �?      �?                               @               @      �?                       @      @      @                              �?      @      @      (@                       @      �?      @      �?      @                              @       @                              �?      @              @                                      �?                                       @      �?      �?                                      �?      @      "@                       @      �?      @      �?      @     @k@      <@     �c@      .@     �@@      @     �D@     �{@     pz@      >@      D@      S@     �x@     `k@      @      8@      5@      Q@      0@     @W@       @     �M@      @      "@      �?      &@     0t@     0p@      @      1@      >@      l@     @Y@              @      @      :@      @     @R@       @     �E@      @      @              "@     �q@     �k@      @      "@      7@     @d@      S@              @      @      4@      @      "@              @                                      N@      F@              �?       @      *@       @                               @              @              @                                      C@      $@              �?              �?                                                      �?                                                      &@      "@              �?              �?                                                      @              @                                      ;@      �?                                                                                      @                                                      6@      A@                       @      (@       @                               @                                                                      @      7@                              @      �?                                              @                                                      .@      &@                       @      @      �?                               @              P@       @      D@      @      @              "@     �k@     `f@      @       @      5@     �b@     �R@              @      @      2@      @     �L@       @     �B@      @      @              @      k@     @e@      @       @      1@     �`@     �R@              @      @      .@      @      6@      �?      .@                              @     �`@     �X@       @       @      @     @S@     �F@              �?      �?      @       @     �A@      �?      6@      @      @              �?     �T@      R@      @      @      *@     �K@      =@              @      @      "@      �?      @              @               @              @      @      "@                      @      1@                                      @               @              @                              @      @      @                      @      $@                                      @              @                               @                      �?       @                              @                                                      4@              0@      @      @      �?       @     �D@      B@               @      @      O@      9@               @              @      �?      *@              &@       @       @      �?       @      0@      2@               @      �?      D@      .@                                              (@              &@       @       @      �?              "@      &@              �?      �?      @@      @                                              (@              $@       @       @      �?               @      $@              �?      �?      8@      @                                                              �?                                      �?      �?                               @                                                      �?                                               @      @      @              �?               @       @                                              �?                                               @      @      @              �?              @      @                                                                                                      @                                      @      @                                              @              @      �?      �?                      9@      2@              @      @      6@      $@               @              @      �?      �?               @      �?      �?                      @      "@              �?      @      *@       @                               @              �?              �?                                      @      @                      @      @       @                              �?                              �?      �?      �?                      @       @              �?       @      "@      @                              �?              @              @                                      2@      "@              @      �?      "@       @               @              @      �?      @               @                                      .@      "@                      �?      @      �?                              �?      �?      �?              �?                                      @                      @              @      �?               @              @             @_@      :@     �X@       @      8@      @      >@     @]@     �d@      9@      7@      G@      e@     �]@      @      2@      .@      E@      (@      B@      (@      .@              @      @      @      >@     �S@      @      $@      ,@     �D@      B@              @       @      @       @      8@      @      (@              �?              @      .@     �H@               @      @      ;@      $@              @               @              0@      @      (@                              @      (@     �G@               @      @      8@      @              �?                              (@       @       @                              @      @      :@              �?      @      ,@       @              �?                              @       @      @                                       @      5@              @              $@      @                                               @                              �?                      @       @                      �?      @      @               @               @                                                                      @      �?                      �?      �?      �?               @                               @                              �?                              �?                               @      @                               @              (@       @      @              @      @      @      .@      >@      @       @      @      ,@      :@              @       @      @       @      (@      @       @                       @              @      :@                      @      $@      0@              @              �?      �?      @       @      �?                       @              @      8@                      @       @      .@              �?                              @      �?      �?                                               @                      �?       @      �?               @              �?      �?              @      �?              @       @      @      "@      @      @       @      @      @      $@              �?       @      @      �?              @      �?              @      �?      @      "@       @      @       @      �?      @      �?              �?      �?      @      �?                                              �?                       @                       @      �?      "@                      �?                     @V@      ,@      U@       @      4@       @      8@     �U@     @U@      5@      *@      @@     �_@     �T@      @      &@      *@     �A@      $@      U@      ,@      P@      @      $@       @      ,@     �Q@     �S@      2@      (@      9@     �]@     �Q@      @       @      $@     �@@      "@     �S@       @     �I@      @       @              *@     @P@     �Q@      @      (@      ,@      Y@     �O@       @      @      @      >@      @      N@      @      B@      @      @              &@     �G@      M@       @      @      $@      N@      B@      �?      @              3@      @      3@      @      .@      �?      @               @      2@      *@      @      "@      @      D@      ;@      �?      @      @      &@      �?      @      @      *@      �?       @       @      �?      @      @      &@              &@      3@       @       @      �?      @      @       @      @      @       @               @       @              @      @      @              @      2@      @       @              �?       @       @       @      �?      @      �?                      �?       @              @              @      �?      @              �?      @      �?              @              4@      �?      $@              $@      0@      @      @      �?      @       @      &@       @      @      @       @      �?       @              .@      �?      @               @      ,@      @      @      �?      �?      @      @              @      @       @      �?       @              $@      �?      �?               @      @      @      @      �?      �?      @      @              @      @              �?                      @              @                      @      �?                               @                                       @              @              @              @               @       @       @                      @      @      @       @                                      @              @              @              @       @       @                      @      @               @                                                      �?              �?              @                                                      @                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ	'thG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         >                   �3@ K1f��?�	           ��@       !                    @ma��x��?|            �@                           �?��Q����?�           p�@                           @�7v~t�?�            �s@                           �?-D*m�?�            @k@                            @t<Z�ï�?H            �]@������������������������       �lY���D�?1            �S@������������������������       �o,x���?            �C@	       
                    @�Q�|�?@             Y@������������������������       �Z��Oԣ�?             ?@������������������������       �Vx�����?)            @Q@                          �1@��U���?A            �X@                           �?����W�?            �C@������������������������       �x�W��#�?             7@������������������������       �      �?             0@                            �?�G��s<�?%            �M@������������������������       ��X�C�?             <@������������������������       ��̿0�=�?             ?@                           �?ݙ�E6�?�             w@                           @P�t]Ec�?9            �U@                          �2@     ��?'             P@������������������������       �ˠT�x?�?             F@������������������������       ����(\��?             4@                          �1@�9����?             6@������������������������       ��������?             @������������������������       �      �?             0@                          �0@�t���E�?�            �q@                           @�in�=�?            �D@������������������������       �T�r
^N�?             <@������������������������       �&�q-�?             *@                             �?��!�z�?�            `n@������������������������       ����X��?H             \@������������������������       �E�p��,�?U            ``@"       /                   �0@��(��?�           І@#       *                    �?���`,�?J            �_@$       '                    �?f�Sc��?            �H@%       &                    @�s��g�?             ;@������������������������       �p=
ףp�?             $@������������������������       ��"�O�|�?             1@(       )                    @;n,�R�?             6@������������������������       �VUUUUU�?             "@������������������������       �޾�z�<�?             *@+       .                    @L�*:�?+            �S@,       -                    @Ϋ�gE#�?"             N@������������������������       �\")�i��?             7@������������������������       �P��a��?            �B@������������������������       �<ݚ)�?	             2@0       7                    �?�R��~�?z           ؂@1       4                   �1@����b��?�            �r@2       3                    @��[.��?D            �Y@������������������������       ����)�?#            �M@������������������������       ���m(�9�?!            �E@5       6                     @�����?}            �h@������������������������       ��3�R��?b             c@������������������������       ��W+J���?            �G@8       ;                    @��ي��?�            �r@9       :                    @L�9���?P            �`@������������������������       �o��L��??            �Y@������������������������       ��������?             >@<       =                    @�E�Z�o�?i            @e@������������������������       ����.��?3            �S@������������������������       ������?6             W@?       Z                    �?wLNĸ�?,           ��@@       K                    �?n~U�B[�?�           t�@A       H                   �?@'Fί���?           py@B       E                     �?�犴ʫ�?�            �w@C       D                   �4@�r����?P             ^@������������������������       ����.�6�?             7@������������������������       �I�/m��?A            @X@F       G                    �?2J	���?�            Pp@������������������������       �=x�u�m�?E             ]@������������������������       ���Mg�?`             b@I       J                    @�h��9�?             :@������������������������       �      �?              @������������������������       �B{	�%��?             2@L       S                    �?�7�wo�?�           0�@M       P                     @4)�/�?�            @t@N       O                     �?�������?g            @e@������������������������       ���,���?\             c@������������������������       ������H�?             2@Q       R                   �;@�G�R/��?e            @c@������������������������       �
FVʫ��?O            �^@������������������������       �     �?             @@T       W                   �8@vEX��x�?            |@U       V                     @xW��:��?�            p@������������������������       ��I�e�H�?F            @\@������������������������       �����H�?Y             b@X       Y                    @1�4����?z             h@������������������������       �5hUN��?7            �U@������������������������       �3+��?�?C            �Z@[       h                     �?���u��?D           ��@\       c                   �=@�-J��?�           ��@]       `                    @�\`Ȇ �?�           �@^       _                    �?�=$w��?           �{@������������������������       ��GBJ���?�            �k@������������������������       �>�&�?�             l@a       b                   �4@@�<��?�            @p@������������������������       �1�*���?!             I@������������������������       ��H*��?�            @j@d       e                    �?#�o�h�?             �J@������������������������       �     ��?
             0@f       g                   �@@"�u�)��?            �B@������������������������       �J��LQ�?             7@������������������������       �^N��)x�?             ,@i       p                    @�����?^           `�@j       m                    �?7�V�<f�?�            �s@k       l                   �:@W�)3��?x            �f@������������������������       �1�/5mv�?e             c@������������������������       ���O��O�?             >@n       o                     @�Sۛ)��?O            �`@������������������������       �$�n��?0            �T@������������������������       �|xV��f�?            �H@q       t                    �?����?�            @n@r       s                     @���Ͷ�?=            �V@������������������������       ���\m��?#            �J@������������������������       �E�r*e�?            �B@u       v                     @�Uo���?Z             c@������������������������       �h�H���?&             O@������������������������       �� �����?4            �V@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F        }@     @R@     �s@      C@     �U@      ;@     �W@     H�@      �@     �P@     �V@     �c@     ��@     0{@      *@      S@     �A@     �^@     �M@     �f@      (@      W@      @      "@              &@     �v@     r@      0@      9@      8@     �h@      `@              6@       @      >@      @     @Y@       @      H@       @      @               @     �]@     �a@      $@      1@      *@     @[@     �Q@              @       @      9@      @      H@      �?      @                              �?     �Q@     �R@      @      @      @      K@     �A@                              "@       @      9@      �?      @                              �?     �K@      G@       @      @      @     �D@      ;@                              @       @      3@               @                                      =@      7@       @      @      �?      .@      1@                              @              (@               @                                      9@      4@              @      �?      @      "@                                              @                                                      @      @       @                       @       @                              @              @      �?      @                              �?      :@      7@                       @      :@      $@                                       @       @                                              �?      @      @                      �?      $@      @                                       @      @      �?      @                                      6@      0@                      �?      0@      @                                              7@               @                                      0@      =@      @              �?      *@       @                               @               @               @                                      @      3@       @                      @      �?                                              @               @                                      @      $@                                      �?                                              �?                                                      �?      "@       @                      @                                                      .@                                                      (@      $@       @              �?      $@      @                               @              (@                                                      @               @              �?      @       @                                              @                                                      @      $@                              @      @                               @             �J@      @     �D@       @      @              �?     �G@     �P@      @      ,@      "@     �K@      B@              @       @      0@      @      4@      �?      "@              �?              �?      (@      2@       @       @      @       @      @               @               @              2@      �?      @              �?              �?      (@      &@               @       @      @      @               @              �?              *@      �?       @                              �?       @       @               @       @      @                                      �?              @               @              �?                      @      @                                      @               @                               @              @                                              @       @              �?       @       @                              �?              �?              �?                                                      �?              �?      �?                                      �?              �?              @                                              @      �?                      �?       @                                             �@@      @      @@       @      @                     �A@     �H@       @      (@      @     �G@      ?@              @       @      ,@      @      @       @                                              @      *@                              "@      @                                              @       @                                               @      @                              "@      @                                              �?                                                       @       @                                       @                                              ;@      @      @@       @      @                      ?@      B@       @      (@      @      C@      8@              @       @      ,@      @      1@              @              �?                      3@      7@      �?      @      @      .@      $@              �?       @      @      @      $@      @      ;@       @      @                      (@      *@      �?      @       @      7@      ,@              @              $@             @T@      @      F@       @       @              "@     �n@     `b@      @       @      &@     �V@     �L@              0@              @       @      6@               @               @                     �Q@      2@                              $@       @                                               @               @                                     �A@      @                              @                                                      �?               @                                      5@       @                              �?                                                                                                              @       @                              �?                                                      �?               @                                      ,@                                                                                              �?                                                      ,@      @                              @                                                      �?                                                      @      @                              �?                                                                                                              $@      �?                               @                                                      4@                               @                      B@      (@                              @       @                                              $@                               @                      ?@      &@                              @                                                      @                               @                      "@      @                              @                                                      @                                                      6@      @                              @                                                      $@                                                      @      �?                                       @                                             �M@      @      E@       @                      "@     �e@      `@      @       @      &@      T@     �K@              0@              @       @      9@       @      3@      �?                       @     @Y@      P@      @      @      @     �C@      ;@              @              �?              "@               @                               @     �F@      ;@                      @      &@      @                                              "@                                               @      >@      ,@                              �?      @                                                               @                                      .@      *@                      @      $@                                                      0@       @      1@      �?                              L@     �B@      @      @      @      <@      8@              @              �?              &@       @       @      �?                             �I@      >@      @       @       @      3@      3@                              �?              @              "@                                      @      @               @      �?      "@      @              @                              A@       @      7@      �?                      @     �R@     @P@              @      @     �D@      <@              (@              @       @      2@              .@                              �?      >@      2@              @      �?      8@      5@                                              1@              ,@                                      :@      ,@              @      �?      3@      @                                              �?              �?                              �?      @      @                              @      ,@                                              0@       @       @      �?                      @      F@     �G@                      @      1@      @              (@              @       @       @               @                                      :@      ;@                      @       @      �?                                       @       @       @      @      �?                      @      2@      4@                              "@      @              (@              @             �q@     �N@     @l@      A@     �S@      ;@     �T@     �g@     0t@      I@     @P@     �`@     �x@     0s@      *@      K@     �@@     @W@      J@     �_@      =@     �]@      7@     �J@      1@      C@      E@     �[@     �@@     �D@     @T@     `d@     @c@      @      B@      7@     �H@      B@      E@      $@      A@      �?      ,@      @      @      3@     �J@      "@      5@      :@     �S@      E@              &@      "@      &@      0@      C@      $@     �@@      �?      "@      @      @      3@      J@      @      3@      2@     �S@      E@              $@      "@      $@      0@      *@      "@      @      �?       @      �?       @      @      ,@              @      @      B@      @              �?      @      @       @      �?              �?                                       @      @                              0@                                                      (@      "@      @      �?       @      �?       @       @      &@              @      @      4@      @              �?      @      @       @      9@      �?      :@              @       @      @      .@      C@      @      *@      .@     �E@     �A@              "@      @      @      ,@      $@      �?      @               @       @       @      $@      :@      �?       @       @      0@      "@              @      �?              "@      .@              3@              @              @      @      (@      @      @      @      ;@      :@              @       @      @      @      @              �?              @                              �?      @       @       @                              �?              �?                                              �?                                      @       @      �?                                              �?              @              �?              @                              �?                      @                              �?                              U@      3@     @U@      6@     �C@      ,@      ?@      7@      M@      8@      4@     �K@      U@      \@      @      9@      ,@      C@      4@      G@      "@      ;@      @      2@              1@      .@      =@              $@      1@      F@     �F@              @      @      5@       @      9@      @      1@       @      @               @       @      @              @      $@      7@      ;@              @       @      .@      @      4@      @      ,@       @      @               @       @      @              @      @      7@      7@              @      �?      .@      @      @              @                                              �?                      @              @                      �?                      5@       @      $@      @      *@              "@      @      6@              @      @      5@      2@              @      @      @      @      *@       @       @      @      @              @      @      6@              @      @      4@      1@                       @      @       @       @               @              @              @                                       @      �?      �?              @      �?              @      C@      $@      M@      0@      5@      ,@      ,@       @      =@      8@      $@      C@      D@     �P@      @      2@      "@      1@      (@      ;@      @     �F@      @      &@      $@      $@      @      1@      ,@      @      (@      4@      J@              @       @      &@      �?      5@       @      2@                              @      @       @      $@      �?      @      @      3@              @      �?       @      �?      @      @      ;@      @      &@      $@      @      �?      "@      @      @      "@      ,@     �@@                      �?      @              &@      @      *@      &@      $@      @      @      @      (@      $@      @      :@      4@      .@      @      (@      @      @      &@      @      @      @      @      "@      �?      �?      @       @      @              @      &@      @      @       @      @      @      @      @       @      "@      @      �?      @      @              @      @      @      5@      "@      $@      @      $@      @              @     �c@      @@     �Z@      &@      9@      $@     �F@     `b@     �j@      1@      8@      J@     �l@      c@      @      2@      $@      F@      0@     �W@      "@     �S@      @       @      @      2@      U@      c@      &@      .@      =@     �]@     �W@              &@      @      4@      @     @V@      "@     �P@      @       @      @      2@      U@     �b@      "@      .@      9@     @[@      T@              "@      @      3@      @     �M@      @     �I@      �?      �?      @      ,@      C@     �Y@      @       @      ,@     �Q@      J@              @              .@              7@      @      >@                              @      .@     �N@       @      @      @      @@     �A@               @              @              B@      @      5@      �?      �?      @      @      7@     �D@      @      @       @     �C@      1@              @              (@              >@      @      0@      @      @              @      G@     �H@       @      @      &@      C@      <@              @      @      @      @      @              �?               @                      $@      @              @       @      1@      @              �?                              7@      @      .@      @      @              @      B@     �F@       @      @      "@      5@      9@              @      @      @      @      @              &@                                              �?       @              @      "@      .@               @      �?      �?      �?      @              @                                                                      �?       @      @               @                      �?      @               @                                              �?       @              @      @      &@                      �?      �?                              @                                              �?       @                      @      @                      �?                      @               @                                                                      @      �?      @                              �?             �N@      7@      =@      @      1@      @      ;@     �O@      N@      @      "@      7@     @\@      M@      @      @      @      8@      (@      H@      ,@      ,@      @      @      @      "@     �A@      D@      @      @      @     �P@      ;@       @      @      @      @      (@      6@      ,@      @       @      @      @      "@      1@      ;@      �?      @      @     �A@      .@              @      @      @      @      5@      @      @       @      @      @      "@      1@      8@      �?       @       @      <@      .@              @       @      �?      @      �?      "@                              �?                      @              @      �?      @                      �?       @       @              :@              @      @      @       @              2@      *@       @               @      ?@      (@       @      �?               @      @      1@              @       @      @                      2@      "@       @                      3@      @      �?                                      "@              �?       @               @                      @                       @      (@      @      �?      �?               @      @      *@      "@      .@              $@              2@      <@      4@      @      @      2@     �G@      ?@      @       @      �?      3@              �?      @      @               @              @      4@      @       @       @      @      9@      ,@              �?      �?                      �?      �?      @               @                      ,@      @      �?              @      .@      "@                                                      @      �?                              @      @      @      �?       @      �?      $@      @              �?      �?                      (@      @      $@               @              .@       @      ,@      �?       @      ,@      6@      1@      @      �?              3@              @       @      @              @              @      @      @      �?       @      @      *@      �?      �?                      @              @      @      @              @              "@      @      @                       @      "@      0@      @      �?              *@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKqhnh4h7K ��h9��R�(KKq��hu�B�         4                   �3@�$�/�~�?�	           ��@                            @V;sq'��?z           ��@                           �?y>У��?z           ��@       	                   �0@޹P)a�?�            �p@                           �?�q�q�?             B@                            �?:J�����?             :@������������������������       �b���i��?             &@������������������������       ����ĳ��?	             .@������������������������       ���Q��?             $@
                            �?�*Y`��?�            @m@                            �?�B����?|             j@������������������������       �Y��sd�?E             ]@������������������������       ��x�W��?7             W@                          �2@M�h���?             :@������������������������       ���"e���?             "@������������������������       �躍`3�?             1@                          �1@��t)0�?�           ��@                          �0@��I���?�            v@                           @�a!���?V             `@������������������������       �PE�Y�?C            �Y@������������������������       �PS!����?             :@                            �?����S`�?�             l@������������������������       �s�n_Y��?c            �c@������������������������       �6c����?(             Q@                           @��0�z"�?�             w@                           @��n�kD�?�            �p@������������������������       �<�T<:��?�            �j@������������������������       ��8���?)             M@                           �?����x��?<            �X@������������������������       �Ό��i�?            �G@������������������������       �N�f��?             �I@        +                    @޷�L���?            �x@!       $                   �0@����`��?�            �r@"       #                    @      �?             @@������������������������       �)O���?
             2@������������������������       ����>4��?	             ,@%       (                   �2@.��B��?�            �p@&       '                    �?�����?�            �g@������������������������       ���+�D��?8            �R@������������������������       ��s-s��?J            �\@)       *                    �?CW���?0            @S@������������������������       �S��d�?             >@������������������������       �5v��?�?            �G@,       1                    @��Z,`�?;            �X@-       0                   �2@x��<��?            �C@.       /                    �?��_�#3�?             =@������������������������       ��������?             1@������������������������       �      �?             (@������������������������       �>
ףp=�?             $@2       3                    @���0�B�?"            �M@������������������������       �>
ףp=�?             D@������������������������       ���|���?	             3@5       T                    �?^�3Q��?-           ��@6       E                    �?��v��?3           P�@7       >                   �;@�We�..�?           �z@8       ;                   �:@������?�            �t@9       :                    �??����?�             s@������������������������       ���4��{�?S             `@������������������������       �B>�٬��?l            �e@<       =                     @������?             ?@������������������������       ��T�x?r�?             6@������������������������       �VUUUUU�?             "@?       B                    �?��x���?2            �W@@       A                   �<@���'�?            �@@������������������������       �
ц�s�?             *@������������������������       ��(\����?             4@C       D                    �?����t��?              O@������������������������       ���.���?             6@������������������������       �      �?             D@F       M                    �?������?/           �}@G       J                    �?�*H~�?�            @m@H       I                    @Y�,�L�?�            �i@������������������������       �C�����?D             Z@������������������������       ��ߖ$��?D            @Y@K       L                   �7@��-�?             =@������������������������       �r�q��?	             (@������������������������       �paRC4%�?	             1@N       Q                    @�gw�e��?�            @n@O       P                   �4@-���+T�?b            �c@������������������������       �Ҿ봜��?            �D@������������������������       ��jC��l�?N            @]@R       S                    �?��X��?3             U@������������������������       ��O�3b��?'            �P@������������������������       �4%���?             1@U       d                   �:@�0@h��?�           L�@V       ]                    �?v��녤�?�           ,�@W       Z                    @X}す9�?]           ��@X       Y                    �?�˰.�L�?�            �q@������������������������       ���5 &��?/            @S@������������������������       �R��q�?�            �i@[       \                   �8@��N�o�?�            @o@������������������������       ��~h���?�            �i@������������������������       �؍����?            �F@^       a                    �?sj{�^��?�           ��@_       `                   �8@��y�}�?K            �]@������������������������       ��;�[AC�??            �V@������������������������       �T�<q,��?             =@b       c                    @O����?W            �@������������������������       �����$}�?5            @W@������������������������       ��2�7���?"           0~@e       j                    �?��ђ�?�            �x@f       i                   @A@(�(� �?Z            �b@g       h                    @&1��?R            �`@������������������������       ���4�i�?!            �N@������������������������       ��q�q�?1             R@������������������������       �v�f��?             1@k       n                   �>@���դ�?�            @n@l       m                    @b�D����?o             d@������������������������       ��cŭT��?T            @]@������������������������       �����!p�?             F@o       p                    @VhΖ�M�?2            @T@������������������������       �5�1	4O�?,            �Q@������������������������       ���!pc�?             &@�t�bh�h4h7K ��h9��R�(KKqKK��h��BC       �z@      R@     �u@      :@     �P@      ;@     �S@     �@     p�@     �T@     �U@     `b@     ��@     �z@      6@     �O@     �F@     �[@      K@      d@      &@     �T@      @      @              $@     �u@     �r@      5@      *@      B@     �l@     �[@              (@      @      ;@       @     @\@      @     �F@       @       @              @     �r@     �k@      .@      "@      =@     �b@     �P@              @      �?      (@      @     �F@      @      1@              �?                     �H@     �L@      @      @      ,@     �E@      4@              @              @      �?       @              �?                                      &@      *@                               @      �?                                              @              �?                                      @      (@                               @                                                      @              �?                                      @      @                                                                                                                                              @      "@                               @                                                      @                                                      @      �?                                      �?                                             �B@      @      0@              �?                      C@      F@      @      @      ,@     �D@      3@              @              @      �?     �B@      @      (@              �?                      ?@      C@      @      @      ,@      D@      0@              @               @      �?      3@      @      @                                      ,@      7@       @      @      @      <@      (@                               @              2@              @              �?                      1@      .@      @      �?      $@      (@      @              @                      �?                      @                                      @      @                              �?      @                              @                               @                                      @      @                              �?                                                                       @                                      @      @                                      @                              @              Q@       @      <@       @      �?              @     �o@     �d@      $@      @      .@     �Z@      G@              @      �?      @      @      @@       @      "@                              @     �a@     @W@              @      "@     �D@      0@                               @       @      3@              �?                                      K@     �B@                      �?      ,@       @                              �?              1@              �?                                     �G@      7@                      �?      *@                                      �?               @                                                      @      ,@                              �?       @                                              *@       @       @                              @     �U@      L@              @       @      ;@      ,@                              �?       @      "@              @                               @     �P@     �A@              @      @      3@      @                              �?       @      @       @       @                              �?      4@      5@                       @       @       @                                              B@              3@       @      �?              @      \@      R@      $@       @      @     �P@      >@              @      �?      @      �?      ;@              $@       @      �?                     @X@     �E@      @       @      @     �J@      3@               @              @      �?      6@              "@       @                             �T@     �B@      @       @      @      A@      "@               @              �?      �?      @              �?              �?                      ,@      @                              3@      $@                               @              "@              "@                              @      .@      =@      @              @      *@      &@              �?      �?                      @              @                                      "@       @      @                       @      @                                               @              @                              @      @      5@                      @      @      @              �?      �?                      H@      @      C@       @      @              @     �H@     �S@      @      @      @      T@      F@              @      @      .@      @     �E@      @      8@       @      @              �?      >@     �I@      @       @      @      O@     �C@              �?      @      .@      @      $@               @               @                      @      �?                              &@      �?                                               @                                                      @      �?                              @                                                       @               @               @                      �?                                      @      �?                                             �@@      @      6@       @      @              �?      9@      I@      @       @      @     �I@      C@              �?      @      .@      @      8@      @      3@      �?       @              �?      7@      ?@       @      �?      @     �D@      8@                      �?      "@      �?      (@               @                              �?      *@      ,@       @                      3@      @                              @              (@      @      &@      �?       @                      $@      1@              �?      @      6@      5@                      �?      @      �?      "@              @      �?      �?                       @      3@      @      �?      �?      $@      ,@              �?       @      @      @      �?                                                      �?      &@                      �?      @       @                              �?      @       @              @      �?      �?                      �?       @      @      �?              @      @              �?       @      @              @              ,@                               @      3@      ;@               @       @      2@      @              @                               @              &@                                      "@      @               @      �?      @       @                                               @              $@                                      @      @                              @                                                       @              @                                      @      @                                                                                                      @                                      �?      �?                              @                                                                      �?                                       @       @               @      �?               @                                              @              @                               @      $@      5@                      �?      (@      @              @                               @              @                              �?      $@      $@                              @      @              @                              �?                                              �?              &@                      �?      @                                                     �p@     �N@     �p@      6@     �M@      ;@      Q@     �k@      t@     �N@     �R@     �[@     �x@      t@      6@     �I@     �D@     �T@      G@     �\@      @@      S@      @      1@      &@      .@      V@      c@      @@      6@      8@      `@     @^@      @      ,@      &@      7@      .@      L@      &@      G@      @      0@       @      "@      5@      I@      1@      .@      ,@      J@     �M@      @      "@       @      3@      (@      G@       @      >@       @      &@      @      @      5@     �C@      &@      @      ,@      I@     �G@       @      @      @      2@      @      E@       @      >@       @      "@      @      @      5@     �@@      "@      @      &@     �D@     �G@       @      @      @      2@      @      5@      �?      0@               @              @      (@      $@       @      @      @      4@      2@               @              "@      @      5@      @      ,@       @      @      @       @      "@      7@      @       @       @      5@      =@       @       @      @      "@              @                               @      �?                      @       @              @      "@                       @       @                      �?                               @                              @      �?              @      @                       @       @                      @                                      �?                              �?                      @                                                      $@      @      0@       @      @       @      @              &@      @      $@               @      (@       @      @      �?      �?      @      @       @      �?                                              @      �?      @               @      "@                                      �?                                                                      �?              @              �?      @                                      �?      @       @      �?                                              @      �?                      �?      @                                              @      �?      .@       @      @       @      @              @      @      @                      @       @      @      �?      �?      @      @      �?       @              @               @               @              @                      @              �?                               @              *@       @       @       @      �?               @      @                                       @       @      �?      �?      @      M@      5@      >@      @      �?      @      @     �P@     �Y@      .@      @      $@      S@      O@              @      @      @      @      ;@       @      (@                               @      A@     @Q@       @      @      @      F@      8@              �?               @              5@      @      $@                               @      :@     �O@       @      @      @     �D@      7@              �?              �?              &@      @      @                               @      @      A@       @              @      5@      *@              �?              �?              $@       @      @                                      5@      =@              @       @      4@      $@                                              @       @       @                                       @      @                              @      �?                              �?              @                                                               @                               @      �?                              �?                       @       @                                       @      @                              �?                                                      ?@      *@      2@      @      �?      @      @     �@@     �@@      *@      @      @      @@      C@              @      @       @      @      0@      $@      (@      �?      �?      @      �?      =@      :@      @      @       @      3@      4@               @       @      �?      @      @                                                      1@      �?              �?              "@      @                                      @      &@      $@      (@      �?      �?      @      �?      (@      9@      @      @       @      $@      .@               @       @      �?              .@      @      @       @                      @      @      @      @               @      *@      2@               @      �?      �?              .@      @      @                              @      @      @      @               @      "@      ,@               @              �?                              @       @                                              @                      @      @                      �?                     �c@      =@      h@      .@      E@      0@     �J@     �`@     @e@      =@      J@     �U@     �p@     �h@      2@     �B@      >@      N@      ?@     �^@      4@     `c@       @      1@      @      C@     �^@     �b@      1@     �@@      O@     `l@      a@       @      :@      4@     �F@      .@     �K@      @      M@      @      @      �?      0@     �R@      T@      @      0@      1@      Z@     �K@              &@      $@      (@      @      ?@      �?      B@      @      @      �?       @      3@      ?@              *@      $@     �O@      @@              &@      $@      @      @      (@      �?       @                      �?      �?      @       @              �?       @      9@      @              @      @      �?       @      3@              A@      @      @              @      *@      7@              (@       @      C@      9@              @      @      @       @      8@      @      6@               @               @     �K@     �H@      @      @      @     �D@      7@                               @              4@      �?      5@              �?              @     �H@     �F@      @              @      ?@      1@                               @              @      @      �?              �?              @      @      @              @      @      $@      @                                              Q@      .@     @X@      @      $@       @      6@      H@     �Q@      *@      1@     �F@     �^@     �T@       @      .@      $@     �@@      &@      .@      @      &@      �?      @      �?      �?      @      @       @       @      @      B@      *@              �?      @      @      @      $@      @      $@      �?      @              �?      �?      @      �?       @      @      5@      *@              �?      @      @      @      @              �?              �?      �?               @              �?              �?      .@                                               @     �J@      $@     �U@      @      @      �?      5@     �F@     @P@      &@      .@      D@     �U@     @Q@       @      ,@      @      =@      @      @       @      .@       @      �?               @      .@      ,@      @      @      @      $@      @                      �?      "@              G@       @     �Q@       @      @      �?      3@      >@     �I@      @      &@     �B@     @S@     �P@       @      ,@      @      4@      @     �@@      "@     �B@      @      9@      *@      .@      (@      3@      (@      3@      9@      E@      O@      $@      &@      $@      .@      0@      3@      @      0@      �?      *@              @      $@      $@              "@      @      ,@      :@      �?       @       @       @      @      1@      @      $@      �?       @              @      $@      $@              "@      @      ,@      7@               @       @       @      @      "@       @      @                                      @      @              @      @              &@               @              @      @       @      @      @      �?       @              @      @      @               @      �?      ,@      (@                       @      �?       @       @              @              @                                                                      @      �?                                      ,@      @      5@      @      (@      *@      (@       @      "@      (@      $@      3@      <@      B@      "@      "@       @      @      &@      *@       @      (@      @      "@      @      "@       @      @      @      "@      @      9@      @@      @      @      @      @       @       @       @       @      @      "@      @      @       @       @      @      "@      @      (@      ;@              @       @       @      @      @              @                              @               @      �?                      *@      @      @       @      @       @      �?      �?       @      "@      @      @      @      @              @      @      �?      .@      @      @      @      @      @      @      @      �?       @      @      @      @      @       @              @      @      �?      *@      @      @      @      @      @      �?      @                      @                              �?                                       @                                               @        �t�bub��(     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJU��4hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         :                    �?9{4�`��?�	           ��@                           �?p.]9�?           \�@                           �?jG�X*��?�           ��@       	                   �1@��l�ߦ�?�            pq@                            @�ܤ�?             E@                           �?�m۶m��?             <@������������������������       �����H�?
             2@������������������������       �p=
ףp�?             $@������������������������       ���>4և�?             ,@
                          �6@W�UM���?�            �m@                           �?G���U�?Q             a@������������������������       �08`�p�?             K@������������������������       �@+�*h�?3            �T@                          �7@B^tJ��??            @Y@������������������������       ��E��ӭ�?
             2@������������������������       ��py�[��?5            �T@                          �3@&a
���?           �z@                          �1@����_�?K             _@                            �?'�Tk��?            �F@������������������������       �Cu��?             5@������������������������       �9��8���?             8@                          �2@Yk'�ؿ�?2            �S@������������������������       �������?            �C@������������������������       �ףp=
��?             D@                           �?�h o��?�            �r@                          �;@��8r��?@            �X@������������������������       ��59���?5            @S@������������������������       �HN�zv�?             6@                           �?B�/O��?�             i@������������������������       ���!pc�?             &@������������������������       ��P�N �?~            �g@        /                   �=@���lp�?c           ��@!       (                    �?���d�#�?-           ��@"       %                   �1@,��>���?�            �s@#       $                     @��S�r
�?             <@������������������������       �k��\��?             1@������������������������       ��g���e�?             &@&       '                     �?��f�*�?�            0r@������������������������       ��x?r���?1             V@������������������������       ��{f��?�            `i@)       ,                    @C�XԀ�?i           ��@*       +                    @0
�p��?�            �u@������������������������       ��_���?�            �n@������������������������       �<�,���?C            �Z@-       .                   �2@�������?�            �j@������������������������       ���JÝ�?             G@������������������������       ��,y���?h             e@0       5                     @c[��V�?6            �X@1       4                   @A@�x�zrJ�?             K@2       3                     �?к����?            �B@������������������������       ��T�6|��?             *@������������������������       ��q�q�?             8@������������������������       �������?             1@6       9                    @�5��;��?            �F@7       8                   @@@K�]l���?             =@������������������������       �؉�؉��?             *@������������������������       �      �?             0@������������������������       �     ��?             0@;       Z                    �?��#X��?�           d�@<       K                    @WOc�!�?�            �@=       D                   �3@���7V�?           `{@>       A                     @bb�#�-�?r             f@?       @                    @ήՊz��?U            @a@������������������������       �}K�Zͺ�?=            �X@������������������������       �\���(\�?             D@B       C                    @��>;���?            �C@������������������������       ��zv�X�?             6@������������������������       �	6c����?             1@E       H                    @%�KG��?�            Pp@F       G                   �8@�����?i            `d@������������������������       �]�l� �?A            �Y@������������������������       �j���&P�?(            �N@I       J                   �:@��
��?B            �X@������������������������       �d�� z�?7            @T@������������������������       ��?�0�!�?             1@L       S                   �5@����<��?�           ��@M       P                     �?#+���?           @{@N       O                   �0@]��d�:�?�            p@������������������������       ��y�ʍ+�?             G@������������������������       �<(s}/��?�            `j@Q       R                   �1@���#�n�?t            `f@������������������������       ��q�1�?             H@������������������������       �F�Y��?U            ``@T       W                    @Xp�b��?�            �k@U       V                   �7@0E�f���?S            �a@������������������������       ��N�?�0�?(             Q@������������������������       ��;�ݩ0�?+            @R@X       Y                    @ҧS�i�?3            @T@������������������������       ����k���?             F@������������������������       ������?            �B@[       j                   �:@��ҋL��?�           ��@\       c                   �6@9B��/#�?p           H�@]       `                     @�%E���?�           ��@^       _                   �1@�v���?_           `�@������������������������       �pӟ�H�?U            @_@������������������������       �ϯ,�5�?
           �z@a       b                    @�ܤ�?j             e@������������������������       ����>�?S            �`@������������������������       �mo�<~'�?            �@@d       g                   �8@���2��?�            �n@e       f                     �?��9!��?h            �a@������������������������       ��}<Sv�?"             G@������������������������       �K�'��n�?F            @X@h       i                    �?|&�{&��??            �Y@������������������������       �w���<�?             ?@������������������������       ���-/e�?-            �Q@k       p                     �?cb�E�C�?b             d@l       o                   �>@�p=
ף�?             D@m       n                   �;@R�@��l�?             ;@������������������������       �������?             ,@������������������������       �g\�5�?             *@������������������������       ��1G����?             *@q       t                     @��h���?L            @^@r       s                   �=@������?3            �S@������������������������       ������*�?             H@������������������������       ���$�d��?             ?@u       v                    @ܶm۶m�?             E@������������������������       ��.sxQ��?             ;@������������������������       �B��S��?             .@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       �{@     �U@     0t@     �E@      S@      =@     @S@     �@     �@      R@     �[@      e@      �@     �}@      5@     @P@      H@      \@     �K@      h@      F@     �d@      9@      I@      2@      B@      `@     `f@     �A@     @Q@      W@     �l@      l@      4@     �C@      ?@      O@      F@      X@      (@      M@       @      ,@      @      3@      S@     �Y@      @      7@      =@     �[@     �U@      @      .@      "@      <@      *@     �E@      @      &@              @      �?       @      B@      K@      @       @      (@     �L@      <@                      �?      @       @      "@              @                                      *@      *@                      �?       @                                                      @               @                                      @      (@                      �?      �?                                                      @               @                                      @      @                      �?                                                                                                                       @      @                              �?                                                      @               @                                      @      �?                              �?                                                      A@      @      @              @      �?       @      7@     �D@      @       @      &@     �K@      <@                      �?      @       @      7@              @               @              �?      *@      :@      �?       @      @      D@      .@                               @              *@              @                                      @      .@                              &@      @                                              $@               @               @              �?       @      &@      �?       @      @      =@       @                               @              &@      @       @               @      �?      �?      $@      .@      @      @      @      .@      *@                      �?      @       @      @                                                              @      �?       @      @              @                                              @      @       @               @      �?      �?      $@      (@       @      @      �?      .@      $@                      �?      @       @     �J@       @     �G@       @      $@       @      1@      D@      H@              .@      1@     �J@      M@      @      .@       @      6@      @      ,@      �?       @                              @      >@      6@                      �?      2@      (@               @              "@      @       @               @                                      0@      @                               @      @                                              @                                                      &@       @                              @      �?                                              @               @                                      @       @                              @      @                                              @      �?      @                              @      ,@      2@                      �?      $@      @               @              "@      @      @      �?       @                              @      @       @                      �?      @                       @              @               @              @                                       @      $@                              @      @                               @      @     �C@      @     �C@       @      $@       @      *@      $@      :@              .@      0@     �A@      G@      @      *@       @      *@       @      <@      @      (@      �?      @              @      @      (@               @       @       @      &@      �?      @              @              3@      �?      (@      �?      @               @      @      $@                       @       @      "@      �?                      @              "@       @                                      �?               @               @                       @              @                              &@      @      ;@      �?      @       @      $@      @      ,@              *@      ,@      ;@     �A@      @      "@       @      @       @                      @                                                                                      @                               @              &@      @      7@      �?      @       @      $@      @      ,@              *@      ,@      ;@      >@      @      "@       @      @       @     @X@      @@     @[@      7@      B@      .@      1@      J@     @S@      ?@      G@     �O@      ^@     `a@      0@      8@      6@      A@      ?@     @X@      =@     @Y@      .@      :@       @      1@      J@     @S@      :@     �B@     �I@      ^@      a@      @      3@      .@      <@      ;@      D@      @     �@@      @      $@      �?       @      6@      =@      @      &@      1@     �L@      A@              @      @      "@      4@      "@                                                      @                              @      (@      �?                                               @                                                      @                              @      "@                                                      @                                                                                              @      �?                                              ?@      @     �@@      @      $@      �?       @      3@      =@      @      &@      ,@     �F@     �@@              @      @      "@      4@      @      @      (@      @      @      �?               @      @              �?      @      3@      @               @      �?      @      @      8@      �?      5@              @               @      &@      8@      @      $@      $@      :@      <@              @      @      @      .@     �L@      6@      Q@      (@      0@      @      "@      >@      H@      5@      :@      A@     �O@     �Y@      @      (@      "@      3@      @     �F@      &@      C@      $@      ,@      @      @      1@     �C@      0@      $@      .@     �D@     �O@      �?      @      "@      @      @      =@       @      5@      @      $@       @      @      (@      ?@      "@      @       @      ?@      G@      �?      @      "@      @      �?      0@      @      1@      @      @      �?              @       @      @      @      @      $@      1@              @                       @      (@      &@      >@       @       @      @      @      *@      "@      @      0@      3@      6@     �C@      @      @              *@      @      @              @                                      (@      @                       @      @      $@               @              �?              @      &@      ;@       @       @      @      @      �?       @      @      0@      1@      3@      =@      @      @              (@      @              @       @       @      $@      @                              @      "@      (@              @      (@      @      @      @      @              �?      @      @      "@      @                                      @      $@               @              @      @      @                      �?       @              "@      @                                      @      @               @              @       @      @                      �?      �?                      @                                      @                                      �?              @                              �?              "@                                               @      @               @               @       @       @                              �?      @                                                              @                               @       @                               @      @       @      �?      @                              @      @       @              �?      (@              @      �?      @               @      @       @      �?      �?                              @       @       @              �?      @              �?              �?               @       @                      �?                              @       @                      �?                                                              @       @      �?                                                       @                      @              �?              �?                                               @                                       @                              @               @      �?      @     �o@     �E@     �c@      2@      :@      &@     �D@      x@     �x@     �B@      E@      S@     �w@     �o@      �?      :@      1@      I@      &@     �]@      1@     �P@       @       @      �?      &@     �n@     �l@      &@      4@      @@     �g@      [@              "@      @      5@      �?      J@      $@      6@       @      @      �?      "@     @Q@     �[@      @      @      ,@      Q@      J@               @      �?      $@              2@      �?      �?      �?                       @      K@     �I@              @      @      :@      "@                              @               @      �?      �?      �?                       @     �F@     �F@              @      @      .@       @                              @              @      �?      �?      �?                       @      B@      :@              @      @      $@      @                               @              �?                                                      "@      3@                      �?      @      @                               @              $@                                                      "@      @                       @      &@      �?                                              @                                                       @      @                               @                                                      @                                                      �?      @                       @      @      �?                                              A@      "@      5@      �?      @      �?      @      .@     �M@      @       @      @      E@     �E@               @      �?      @              2@       @      4@      �?      @      �?       @      &@      >@               @      @      9@     �@@               @               @              *@      @       @      �?       @      �?              @      9@                      @      3@      1@                               @              @      @      (@              �?               @      @      @               @      �?      @      0@               @                              0@      �?      �?              @              @      @      =@      @               @      1@      $@                      �?      @              .@      �?      �?              @              �?      @      ;@      @               @      (@      "@                      �?       @              �?                                              @      �?       @      �?                      @      �?                               @             �P@      @      F@               @               @      f@     @^@      @      .@      2@     �^@      L@              @       @      &@      �?      I@      �?      7@               @               @     �a@     �R@       @      "@      *@     �T@      8@              @               @              D@      �?      @                               @     �P@      H@       @      @      (@      L@      (@               @              @              "@                                                      5@       @                               @                                                      ?@      �?      @                               @      G@      D@       @      @      (@      H@      (@               @              @              $@              0@               @                     �R@      ;@              @      �?      :@      (@              �?              @              @              �?                                      :@       @                              $@                                                      @              .@               @                     �H@      3@              @      �?      0@      (@              �?              @              1@      @      5@                                     �A@      G@      @      @      @      D@      @@              @       @      @      �?       @      @      .@                                      7@      D@      @      @      @      6@      .@              �?       @      �?      �?       @       @      �?                                      &@      6@                              ,@      *@                       @              �?      @       @      ,@                                      (@      2@      @      @      @       @       @              �?              �?              "@       @      @                                      (@      @      �?      @       @      2@      1@              @               @               @               @                                      &@       @                       @      *@      &@                              �?              @       @      @                                      �?      @      �?      @              @      @              @              �?             �`@      :@     �V@      0@      2@      $@      >@     �a@      e@      :@      6@      F@     �g@     @b@      �?      1@      ,@      =@      $@      ]@      2@     �R@      .@      .@       @      :@     `a@      d@      (@      2@      @@     @f@     �]@      �?      *@      @      1@      @     �V@      &@      M@      ,@       @      �?      1@     @]@     �`@       @      ,@      8@      \@     �W@              @      @      @      @     �R@      @      E@       @       @      �?      *@     @Y@     �Z@       @      $@      3@     @S@     �Q@              @      @      @      @      0@                                               @      B@     �A@              �?      @      7@       @                                      �?      M@      @      E@       @       @      �?      &@     @P@      R@       @      "@      0@      K@      O@              @      @      @       @      0@      @      0@      @      @              @      0@      <@              @      @     �A@      8@                              �?       @      *@      @      0@      @      @              @      (@      .@              @      @      ;@      6@                              �?       @      @       @                      �?                      @      *@                               @       @                                              :@      @      1@      �?      @      �?      "@      6@      9@      @      @       @     �P@      9@      �?      @       @      (@      �?      9@      @      $@      �?      �?              @      $@      1@      �?      @      @      C@      (@      �?      @              @      �?       @       @      @      �?                              @       @              @      @      @      @              @               @              1@      @      @              �?              @      @      .@      �?               @      ?@      "@      �?                      @      �?      �?      �?      @              @      �?      @      (@       @      @      �?      @      <@      *@              @       @      @                              �?              @      �?       @      @       @      @                      @      @               @       @                      �?      �?      @              �?              @      @      @              �?      @      9@      "@               @              @              3@       @      .@      �?      @       @      @      �?       @      ,@      @      (@      $@      ;@              @      @      (@      @      @              �?              �?      @                               @              �?      @      @                      @      �?       @      @                                      @                              �?              �?       @      @                      @               @      @                                      @                              �?              �?      �?       @                                                                                                                                              �?      @                      @               @      �?              �?              �?                                      @                      �?      �?                              �?              .@       @      ,@      �?       @       @      @      �?       @      @      @      &@      @      4@              @      �?      &@       @      (@      @      *@      �?      �?                              @      @      @      @      @       @              @      �?       @      �?      &@      @      @              �?                               @      @      @               @      @              @              @      �?      �?      �?      @      �?                                      @       @              @      @      @                      �?       @              @      @      �?              �?       @      @      �?       @                      @       @      (@                              @      �?      @                              �?              @      �?      �?                      @              &@                               @      �?              @      �?                       @      �?              �?                      @       @      �?                              �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ-
thG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmK{hnh4h7K ��h9��R�(KK{��hu�B�         @                    �?�8��g��?�	           ��@       !                   �7@s���)�?           0�@                          �1@�H�����?�           4�@                            @Bb��c>�?q             g@                           �?/y0��k�?@             Z@                            �?333333�?             D@������������������������       �+7����?             7@������������������������       ��P�n#�?             1@	       
                     �?     ��?%             P@������������������������       �(��&y��?             =@������������������������       �p�
���?            �A@                          �0@�P���?1            @T@                           @
ףp=
�?             9@������������������������       �0�����?             ,@������������������������       �*L�9��?             &@                           �?և���X�?$             L@������������������������       ��2�tk~�?             2@������������������������       �]��N��?             C@                           �?Q�����?           ��@                           �?�=%�II�?�            0u@                          �6@��:���?S            �a@������������������������       �a�,�q�?H            @\@������������������������       �N�7��?             =@                            �?����R�?w            �h@������������������������       �z-SO�w�?#            �N@������������������������       ��ɜoB�?T             a@                           @̯����?F           �@                           �?i��`��?�            `t@������������������������       ���@t�?Z            �a@������������������������       �#5@����?s             g@                             @JoN�w�?y            `g@������������������������       ��s7��?B            �X@������������������������       �]t�E�?7             V@"       1                   �=@�-i���?�           ��@#       *                    �?���:��?=           �~@$       '                   �:@k�=F?��?j             e@%       &                    @7�A�0�?:             V@������������������������       ��^��"��?+             Q@������������������������       ����Q��?             4@(       )                    @>
ףp=�?0             T@������������������������       ��r
^N��?"             L@������������������������       �      �?             8@+       .                    �?|H+�N�?�            pt@,       -                   �9@Z��P���?Z            �`@������������������������       ����:�0�?+            @P@������������������������       ����l��?/            �Q@/       0                   �8@UUUUU	�?y             h@������������������������       ��}�AV7�?!            �H@������������������������       �l!M�q�?X            �a@2       9                   �>@��8���?\             b@3       6                     �?�}<Sv�?             G@4       5                    �?9��8���?             8@������������������������       ��9����?             &@������������������������       �g\�5�?             *@7       8                    �?&ޏ���?             6@������������������������       �      �?              @������������������������       �I�$I�$�?             ,@:       =                    @������?C            �X@;       <                     @w�J���?$            �I@������������������������       �     ��?             @@������������������������       �/�s��?             3@>       ?                     @�a��d�?            �G@������������������������       �:߄*�u�?             A@������������������������       ��K8��?             *@A       ^                    �?���k��?�           z�@B       O                   �2@��Z&?�?�           x�@C       J                    @<,�s��?�            �t@D       G                   �0@>W����?�            �p@E       F                    �?�1y)�+�?-            �O@������������������������       ����Q��?             D@������������������������       ����C4�?             7@H       I                     @��V_!�?�            �i@������������������������       ��d���?q            �d@������������������������       �^����T�?            �C@K       N                    @R7�f��?'            @P@L       M                     �?iQT����?            �E@������������������������       ����d�?             ;@������������������������       �     ��?             0@������������������������       ��ˠT��?             6@P       W                   �8@W��ٯ��?�           ��@Q       T                   �7@���vQ{�?[           ��@R       S                    @L߆�{b�?5           `}@������������������������       �*St�ó�?@            �X@������������������������       �DA�Ezu�?�            @w@U       V                    @����"��?&             O@������������������������       ��T�l��?            �@@������������������������       ��c�Α�?             =@X       [                     �?�>��E��?u            �g@Y       Z                   �:@�	��-��?E            �[@������������������������       �гY����?             I@������������������������       ��X�%��?'             N@\       ]                    @�@�f�l�?0            �S@������������������������       ��6��D�?             5@������������������������       �y�ǋ��?$            �L@_       n                   �5@>��G~�?�           |�@`       g                    @���ؠ�?�           �@a       d                     @���Z�?           �|@b       c                    �?���M�)�?�            �v@������������������������       �q�i��?r            �f@������������������������       �(��yL�?l             f@e       f                    @k�%�?9            �X@������������������������       ���X��?             <@������������������������       �ihx�ҙ�?(            �Q@h       k                    @��ԇ}��?�            �n@i       j                    @.�袋.�?3             V@������������������������       �d���?             ;@������������������������       �s����)�?             �N@l       m                   �0@~��#���?m            �c@������������������������       �T�r
^N�?             ,@������������������������       �rH��7�?f             b@o       v                    @ b+Rq�?$           �}@p       s                   �9@X�I� ��?�            �q@q       r                    �?�������?_            `c@������������������������       �����|��?             F@������������������������       �tO�s�?D            �[@t       u                     �?��^-#�?K            �`@������������������������       �t|��?%            �Q@������������������������       �q�g+��?&            �N@w       x                     �?�t/�F��?z            �g@������������������������       ���'����?             G@y       z                     �?�E�����?^             b@������������������������       �>@�?��?            �E@������������������������       � �����?C            @Y@�t�bh�h4h7K ��h9��R�(KK{KK��h��BI       �}@     �T@     �s@      ;@      S@     �E@      X@     �~@     ��@      O@      V@     `e@     Ђ@     �y@      ,@     �R@     �C@     @a@     �Q@     `j@      E@     �d@      &@      G@     �@@      G@     @[@     @h@      =@      K@     @W@      n@     �h@      @     �D@      <@     �R@      K@     �a@      5@     �Y@      @      3@      3@      1@     �X@     �c@      *@      ?@     �G@     `d@     �\@              3@       @     �E@      0@      =@       @      @              @              �?     �B@      ?@      �?       @      $@      B@      5@                               @       @      *@               @               @              �?      :@      4@      �?              @      7@      @                                       @      @               @                                      $@      $@      �?              @      @       @                                               @               @                                       @      @                       @      @       @                                              @                                                       @      @      �?               @      �?                                                      @                               @              �?      0@      $@                      @      3@      @                                       @      @                                              �?       @      @                              "@      @                                              @                               @                       @      @                      @      $@      �?                                       @      0@       @      @              @                      &@      &@               @      @      *@      ,@                               @              &@       @      �?                                      @       @                                      @                                              $@       @                                               @                                                                                              �?              �?                                      @       @                                      @                                              @              @              @                      @      "@               @      @      *@      &@                               @              @                                                      �?      @                       @      @      �?                                               @              @              @                      @      @               @      �?       @      $@                               @              \@      3@     @X@      @      ,@      3@      0@      O@     �_@      (@      =@     �B@     �_@     @W@              3@       @     �D@      ,@     �F@      @      <@      �?      @              @      <@     @Q@       @      $@      .@      L@     �@@              "@       @      $@      $@      2@              *@                               @      2@      8@      @       @      @      >@      ,@              @              @      �?      "@              &@                               @      2@      5@      @       @      @      ;@       @              @              @      �?      "@               @                                              @       @              @      @      @                                              ;@      @      .@      �?      @              @      $@     �F@      @       @       @      :@      3@              @       @      @      "@      "@      @      "@      �?                      �?      �?      $@                      �?      ,@      @                              @       @      2@       @      @              @              @      "@     �A@      @       @      @      (@      .@              @       @              @     �P@      ,@     @Q@      @      &@      3@      "@      A@     �L@      @      3@      6@     �Q@      N@              $@      @      ?@      @      H@      (@      ?@      @      @      $@      @      8@      G@       @      "@      ,@      G@     �@@              "@      @      1@      @      2@      @      "@              @       @       @      3@      6@              @      @      :@      &@              @       @      @      @      >@      "@      6@      @      @       @      @      @      8@       @      @       @      4@      6@              @      @      $@              3@       @      C@       @      @      "@      @      $@      &@       @      $@       @      9@      ;@              �?      �?      ,@      �?      0@      �?      4@              �?               @      $@      @              @       @      $@      ,@              �?      �?      @      �?      @      �?      2@       @      @      "@      �?              @       @      @      @      .@      *@                              @             �Q@      5@      P@      @      ;@      ,@      =@      $@     �B@      0@      7@      G@     @S@     �T@      @      6@      4@      @@      C@     �O@      4@     �H@       @      3@       @      6@      $@      ?@      &@      $@      @@     @R@     �R@      @      ,@       @      1@      <@      <@      "@      (@              &@       @      @      @      @      @      @       @      @@      5@              @      @      "@      $@      "@      @      @              @       @              @      @       @      @      �?      6@      *@              @      �?       @      @      "@      @      �?              @       @              @       @      �?      @      �?      1@      *@               @      �?      @       @              �?       @                                               @      �?      �?              @                      �?              @       @      3@      @      "@              @              @       @       @       @      �?      �?      $@       @              �?       @      �?      @      @      @      "@              @              �?       @      �?       @      �?      �?      @      @                       @      �?      @      (@                                              @              �?                              @      @              �?                             �A@      &@     �B@       @       @      @      2@      @      9@      @      @      >@     �D@      K@      @      $@      @       @      2@      6@      @      0@              �?              "@              1@              �?      $@      2@      1@              @      @      @      "@      @              @                              @              (@              �?      "@      @      (@              @      @       @      @      1@      @      &@              �?              @              @                      �?      .@      @                              �?      @      *@      @      5@       @      @      @      "@      @       @      @      @      4@      7@     �B@      @      @       @      @      "@      @              @               @              �?      @      �?       @      �?       @      @      4@                              �?              "@      @      0@       @      @      @       @              @      @      @      2@      1@      1@      @      @       @      @      "@      @      �?      .@       @       @      @      @              @      @      *@      ,@      @       @      @       @      (@      .@      $@      @              @               @       @       @              @              @       @       @      @               @              $@       @                       @                       @       @              @                      �?              @              �?              @       @                      �?                               @              @                      �?               @                                       @                      �?                       @                      �?                                      �?              �?              @              @              @               @                                              @      �?       @      @              �?              @              @                                                                              �?      �?       @                      �?                                              @               @                                               @                      @                              @              @      �?      "@       @      @      @      @               @      @      $@      (@       @       @      @      @      (@      @       @      �?      �?      @              �?               @              �?      @      "@       @       @       @       @      @      �?      @      @      �?      �?       @              �?               @                       @      @       @       @      �?               @              @      �?                       @                                              �?      @      @                      �?       @      @      �?              @      @              @       @      @      @      @              �?              �?      @                      �?      �?      &@       @      @      @              @       @       @      �?       @              �?                      @                              �?      $@       @       @                      �?              @      @      �?                              �?                              �?              �?               @     �p@     �D@     �b@      0@      >@      $@      I@     x@      {@     �@@      A@     �S@     �v@      k@       @     �@@      &@     �O@      0@      _@      *@     �R@       @      @       @      "@     �k@     @m@      2@      2@      @@     �e@     @V@              $@      @      3@      @      E@      �?      2@                                     @[@     @V@      @       @      @      J@      (@                              �?             �@@      �?      2@                                     @X@      O@      �?       @      @      E@      "@                              �?              "@              @                                      ?@      $@               @               @                                                      @              @                                      3@      @               @              @                                                      @                                                      (@      @                              �?                                                      8@      �?      .@                                     �P@      J@      �?              @      A@      "@                              �?              3@      �?      @                                      L@      F@      �?              @      :@      "@                              �?              @               @                                      $@       @                               @                                                      "@                                                      (@      ;@       @               @      $@      @                                              @                                                      @      8@                       @      @      @                                                                                                       @      4@                       @              @                                              @                                                      @      @                              @                                                      @                                                      @      @       @                      @                                                     �T@      (@      L@       @      @       @      "@     �[@      b@      .@      0@      ;@     �^@     @S@              $@      @      2@      @      N@      @      D@               @       @      @      X@     @]@      (@      @      1@     @V@      L@              @      @      .@      �?      K@      @      @@               @       @      @     @T@     @Z@      "@      @      1@      V@      F@              @      @      *@      �?      (@      �?      @                       @              &@      <@      �?              @      4@      @                              @              E@      @      :@               @              @     �Q@     @S@       @      @      (@      Q@     �B@              @      @       @      �?      @               @                               @      .@      (@      @                      �?      (@              �?               @              @              @                                      *@      @      @                      �?      @                                              �?              @                               @       @      @                                      "@              �?               @              6@       @      0@       @      @              @      .@      <@      @      "@      $@      A@      5@              @              @      @      (@       @      *@       @                      @      &@      5@       @      @      @      &@      (@              @               @       @       @              @                              @       @      .@              @      �?      @       @               @              �?              $@       @      @       @                              "@      @       @       @      @      @      @               @              �?       @      $@      @      @              @                      @      @      �?      @      @      7@      "@               @              �?      �?              �?                      @                      �?       @              �?      �?      @      @              �?                              $@      @      @                                      @      @      �?       @       @      1@      @              �?              �?      �?      b@      <@     �R@      ,@      7@       @     �D@     �d@      i@      .@      0@      G@     `g@      `@       @      7@      @      F@      (@     �V@       @     �B@      @      @      @      2@     �a@      b@      @      $@      9@     �Y@     �Q@              (@      @      ,@      "@      O@      @      7@       @       @      @      ,@     @Y@     �U@       @      @      (@      S@      G@               @               @      @     �I@      @      1@               @      @      &@     @U@     �R@       @      @      $@      H@     �B@              @               @      @      2@               @               @      @      @      G@     �E@       @              @      2@      8@              @              �?      @     �@@      @      "@                              @     �C@      ?@              @      @      >@      *@              �?              �?              &@      �?      @       @                      @      0@      *@              @       @      <@      "@              @                       @      �?      �?      �?                              �?      @      @                       @      (@      �?                                              $@              @       @                       @      *@      @              @              0@       @              @                       @      <@       @      ,@      @      @              @      E@      M@      �?      @      *@      ;@      8@              @      @      (@      @      $@              @      @      �?              @       @      <@      �?      �?              @      3@                               @              @               @                                      @      @      �?                       @       @                                              @              @      @      �?              @       @      8@              �?              @      &@                               @              2@       @      @       @       @              �?      A@      >@              @      *@      6@      @              @      @      $@      @      @                              �?                       @                                                                                              *@       @      @       @      �?              �?      :@      >@              @      *@      6@      @              @      @      $@      @      K@      4@     �B@      @      2@      @      7@      6@     �K@      (@      @      5@      U@      M@       @      &@      @      >@      @      C@       @      0@      @      (@      @      &@      (@      E@       @      @      &@      C@     �E@      @      @      �?      2@       @      5@      @      @      @      @      �?      "@      @      B@      �?      @      @      :@      5@               @              @              (@      @      �?                      �?      �?       @      @                              @      "@               @                              "@       @      @      @      @               @      @      >@      �?      @      @      5@      (@                              @              1@      �?      $@      �?      "@      @       @      @      @      @       @      @      (@      6@      @      @      �?      .@       @      (@              @              @      �?              �?              @      �?      @      "@      ,@              @              "@              @      �?      @      �?      @       @       @      @      @       @      �?      @      @       @      @      �?      �?      @       @      0@      (@      5@       @      @              (@      $@      *@      @              $@      G@      .@       @      @      @      (@      �?      �?              @      �?                      @       @      �?      �?                      @       @              @      �?      @              .@      (@      ,@      �?      @              "@       @      (@      @              $@      D@      @       @       @       @      @      �?      @      @      @               @                      �?      @      �?              @      $@       @                       @      �?              (@       @       @      �?      @              "@      �?       @       @              @      >@      @       @       @              @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�zhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKuhnh4h7K ��h9��R�(KKu��hu�B�         >                    @C�5�ۍ�?�	           ��@       !                    �?�_�Q���?�           �@                           �?Y���
�?.           ��@                           �?�_��b�?�           ��@                          �1@&�ׁS��?�            Pq@                           @\����$�?            �C@������������������������       ��d�����?             3@������������������������       ��G�z�?             4@	       
                    �?N����?�            �m@������������������������       ����H�~�?:            @V@������������������������       �Ң�#�j�?b            �b@                            �?�|#ʯ�?�            t@                          �;@K����?=            �V@������������������������       �5eӏ��?3            @S@������������������������       ��>4և��?
             ,@                            @�������?�            �l@������������������������       �Y���_�?T            @^@������������������������       ���JMu�?G            @[@                           �?ማ��E�?�           h�@                          �2@�x=K^��?           p{@                          �0@�|�j��?7            �V@������������������������       ����(\��?             $@������������������������       �\���(�?0             T@                            �?c�ؔ���?�            �u@������������������������       �m�/K�]�?=             ]@������������������������       �~���l��?�             m@                           @#(��mX�?�           �@                          �:@���R:�?�            `r@������������������������       ���c%���?�            �n@������������������������       � �p?��?#            �H@                           �;@���}��?�            �s@������������������������       �r�Hǉ�?�            `p@������������������������       ��"��ǵ�?'            �K@"       1                   �4@+��&^>�?Z           ��@#       *                     @��(\h�?�            0q@$       '                   �0@�*;�1R�?{            �g@%       &                     �?�.v�P��?            �B@������������������������       ���ˠ�?             6@������������������������       ��h$���?	             .@(       )                    @�ZY2��?f             c@������������������������       ��b)0��??            �W@������������������������       �H���?'            �L@+       .                    @<�D�^��?1            �U@,       -                    �?R=6�z�?%            @P@������������������������       �$6M5��?            �D@������������������������       �r�q��?             8@/       0                    �?4և����?             5@������������������������       �ףp=
��?             $@������������������������       ��ˠT�?             &@2       9                    �?��l��?�            �p@3       6                     �?     r�?T             `@4       5                    @NI8d�?            �B@������������������������       ����(\��?             $@������������������������       ���k���?             ;@7       8                    @�v����?:            �V@������������������������       ���l���?%            �M@������������������������       �     ��?             @@:       =                   �?@ֶ�+{0�?Z            `a@;       <                     �?�ۏ��?Q            �^@������������������������       �\��[���?            �C@������������������������       �[T�D$��?7            �T@������������������������       �� =[y�?	             1@?       X                    @��rd��?J           �@@       K                   �0@=6\�?�           ��@A       F                    @Υ�,v�?B            @Y@B       E                    �?�7p��?            �E@C       D                    @8�Z$���?             :@������������������������       �*D>��?             *@������������������������       ��؉�؉�?	             *@������������������������       �/k��\�?             1@G       H                    @�5д>�?&             M@������������������������       ��m۶m��?             ,@I       J                     �?d�
��?             F@������������������������       �4և����?             5@������������������������       �K����?             7@L       S                   �7@��ы4j�?�           ,�@M       P                     @O�Vn;��?           Љ@N       O                    @��Y�`�?�           p�@������������������������       �BX����?           @z@������������������������       �Ӛ�H��?�            �p@Q       R                    �?]�l8b��?]            �a@������������������������       ��� ֤�?&            �L@������������������������       ���^d��?7            �T@T       W                   �@@����?�             j@U       V                    �?ƪ�6���?{             h@������������������������       ��s�����?7            �U@������������������������       � g���N�?D            �Z@������������������������       �      �?	             0@Y       h                   �8@�2�$��?k           X�@Z       a                   �6@����T�?           �|@[       ^                    �?&�����?�            �v@\       ]                    �?+����?w            �g@������������������������       ���2���?/            @S@������������������������       �����J.�?H            @\@_       `                   �2@���^=�?n            @e@������������������������       ����v��?(             O@������������������������       ��u0f���?F             [@b       e                    @�dm�Ƹ�?8            �X@c       d                     @�%y=d��?            �E@������������������������       �R?��yq�?            �A@������������������������       �      �?              @f       g                     @.~��zE�?!            �K@������������������������       ��Ł�r��?             C@������������������������       �|�l�]�?	             1@i       n                    �?θ�|C�?N             `@j       k                     �?cT!)��?             C@������������������������       ��q�q�?             (@l       m                   �:@o_Y�K�?             :@������������������������       �     @�?             0@������������������������       ��������?             $@o       r                     �?��8~�v�?9            �V@p       q                   �:@     ��?             @@������������������������       �0�����?             @������������������������       ��?�߾�?             9@s       t                    @OK�6��?$            �M@������������������������       ��T�6|��?             :@������������������������       �ڣ����?            �@@�t�bh�h4h7K ��h9��R�(KKuKK��h��BxE        {@     �S@     �s@      ;@     @S@      6@     �R@     Ђ@     ��@     @Q@     �V@      b@      �@     �z@      1@      R@      M@     �`@      N@     @m@     �H@     �i@      ,@      N@      4@      G@     �l@     �q@     �D@      N@     �X@     @v@      q@      $@      E@     �F@     �T@      G@     �f@     �@@     �b@      &@      K@      .@     �B@     �c@     �f@      =@     �J@     �T@     �p@     �i@       @      B@     �C@     �P@      F@     �S@      (@      G@              .@              "@     @P@     �U@       @      2@      8@     �^@      M@              &@      "@      5@      0@      A@      @      2@              @              @      G@     �J@      @       @      @      N@      2@              @      �?      @       @       @              @                                      0@      "@                               @                                                      @              @                                      @      @                               @                                                       @              �?                                      (@      @                                                                                      :@      @      ,@              @              @      >@      F@      @       @      @      M@      2@              @      �?      @       @      @      @      $@                                      (@      5@      �?      @      �?      2@      @               @      �?       @      @      5@      �?      @              @              @      2@      7@       @      @      @      D@      (@               @              @      @      F@       @      <@              (@              @      3@     �@@      @      $@      2@      O@      D@              @       @      ,@       @      @       @       @              @               @      &@      @               @      @      4@      $@               @      @      @       @      @       @      @               @              �?      &@      @                      @      4@      $@                      �?      @       @      �?              �?              @              �?                               @      �?                               @       @                     �B@      @      4@              @              @       @      <@      @       @      (@      E@      >@              @      @      "@      @      5@      �?       @              @               @      @      1@       @      @      "@      5@      .@              @              @      @      0@      @      (@              @              �?       @      &@      @      @      @      5@      .@              �?      @      @       @     �Y@      5@     �Y@      &@     �C@      .@      <@      W@     @X@      5@     �A@      M@     �a@     �b@       @      9@      >@     �F@      <@     �K@      @      A@      @       @              .@     �J@     �I@              0@      2@     @R@     �H@       @       @      .@      0@      0@      1@      �?       @                              �?      ;@      3@                       @      &@      @               @              @                                                                      @      �?                               @      �?                                              1@      �?       @                              �?      5@      2@                       @      "@       @               @              @              C@      @      @@      @       @              ,@      :@      @@              0@      0@      O@      G@       @      @      .@      &@      0@      1@      �?       @       @      �?              @      &@      *@              "@      @      :@      @               @      @      @      @      5@      @      8@       @      @               @      .@      3@              @      (@      B@     �E@       @      @      &@      @      &@      H@      .@     @Q@      @      ?@      .@      *@     �C@      G@      5@      3@      D@     �Q@     �X@      @      1@      .@      =@      (@     �@@       @      4@       @      3@      @      @      ;@      <@      "@      @      &@     �A@     �F@      @       @      "@      3@      @      @@       @      2@      �?      @       @      �?      ;@      ;@      @      @       @     �A@     �C@      @      @      @      1@      �?      �?               @      �?      ,@       @       @              �?      @              @              @      �?      @      @       @       @      .@      @     �H@      @      (@      &@      $@      (@      2@      (@      (@      =@     �A@      K@       @      "@      @      $@      "@      .@      @      H@       @       @       @      "@      (@      1@      &@      $@      3@      A@     �H@              @      �?      "@      @                      �?      @      @      "@      �?              �?      �?       @      $@      �?      @       @      @      @      �?      @     �J@      0@     �K@      @      @      @      "@      R@     �X@      (@      @      0@     �V@     �P@       @      @      @      1@       @      =@      @      5@       @      �?      @      �?      J@      P@      @      �?       @     �E@      :@              �?      @      &@      �?      5@              1@       @      �?                      B@     �G@      @      �?      @      6@      3@              �?      @      "@      �?      @              @                                      @      1@              �?              @                                                                                                              @      &@              �?              @                                                      @              @                                       @      @                              �?                                                      2@              ,@       @      �?                      =@      >@      @              @      0@      3@              �?      @      "@      �?      "@              $@                                      7@      5@                      @      *@      "@              �?               @      �?      "@              @       @      �?                      @      "@      @                      @      $@                      @      @               @      @      @                      @      �?      0@      1@                       @      5@      @                               @               @      @      @                      @      �?      0@      $@                              0@      @                                               @                                      @              $@       @                              $@       @                                                      @      @                              �?      @       @                              @      �?                                                              �?                                              @                       @      @      @                               @                                                                              @                       @      @                                                                      �?                                               @                               @      @                               @              8@      &@      A@      �?      @       @       @      4@      A@      "@      @       @      H@      D@       @      @      @      @      �?      (@      "@      0@               @              �?      $@      3@              @      �?      =@      7@               @              �?               @      @      �?              �?              �?      �?      "@               @      �?       @      @                              �?                                                                              @                      �?      @                                                       @      @      �?              �?              �?      �?      @               @              @      @                              �?              $@      @      .@              �?                      "@      $@              �?              5@      1@               @                               @      @      *@                                      @       @              �?              "@      &@              �?                               @               @              �?                      @       @                              (@      @              �?                              (@       @      2@      �?      @       @      @      $@      .@      "@      @      @      3@      1@       @      @      @      @      �?      (@       @      0@      �?      @       @      @      $@      .@       @      @      @      1@      *@              @      @      @      �?      @              "@               @      �?      @      �?       @              @      �?      @      @                       @                      "@       @      @      �?      �?      �?              "@      *@       @              @      *@      "@              @      �?      @      �?                       @                                                      @                       @      @       @                                      i@      >@     @\@      *@      1@       @      =@     Pw@     �s@      <@      >@      G@      p@     @c@      @      >@      *@      I@      ,@     �]@      5@     �Q@      &@      @      �?      0@     �q@      n@      (@      7@      ?@     �e@     �W@      @      @      @      *@      @       @              @               @                      M@      7@                              @      �?                              �?              @                               @                      6@      (@                               @                                                       @                                                      0@       @                                                                                      �?                                                      @      @                                                                                      �?                                                      "@      @                                                                                      @                               @                      @      @                               @                                                      @              @                                      B@      &@                              @      �?                              �?                                                                      &@       @                              �?                                                      @              @                                      9@      "@                               @      �?                              �?               @              @                                       @      @                               @      �?                              �?              �?                                                      1@      @                                                                                     �[@      5@     �P@      &@      @      �?      0@     �k@      k@      (@      7@      ?@     @e@     @W@      @      @      @      (@      @     �W@       @     �G@      @                      &@     �i@     �f@       @      2@      7@     �a@     �P@               @       @       @      @     @T@      @      :@       @                      "@     �f@     �c@       @      (@      .@     @]@     �K@               @       @      @      @     �P@      @      1@       @                      "@     �W@     �T@      @      &@      .@     @Q@      B@               @      �?      @      @      .@      @      "@                                      V@     �R@      @      �?              H@      3@                      �?      @              *@      �?      5@      @                       @      7@      9@              @       @      7@      &@                               @      �?      @               @                                      2@      $@              @               @      @                              �?              "@      �?      *@      @                       @      @      .@               @       @      .@      @                              �?      �?      1@      *@      4@      @      @      �?      @      1@      A@      @      @       @      >@      ;@      @      @      @      @      �?      .@      (@      1@      @      @              @      1@      A@      @      @       @      >@      5@      @      @      @      @      �?       @      @       @               @              @      .@      "@      �?       @       @      (@      (@               @              @      �?      @      @      "@      @      @               @       @      9@       @      @      @      2@      "@      @      �?      @      �?               @      �?      @                      �?                              �?                              @               @                             @T@      "@     �E@       @      $@      �?      *@     @W@     �S@      0@      @      .@     @T@      N@      @      7@      @     �B@       @     �R@      @      5@       @      $@              @     �T@     �Q@      @       @      &@     @Q@     �F@      @      2@       @      ?@      �?     �I@       @      0@       @       @              @     �R@      O@      @       @       @      J@     �C@              0@      �?      0@      �?      4@               @                              @      J@     �B@      @       @      @      =@      4@              @              @              $@               @                                      :@      &@                      �?      &@      0@                                              $@              @                              @      :@      :@      @       @      @      2@      @              @              @              ?@       @       @       @       @               @      6@      9@                       @      7@      3@              *@      �?      &@      �?      $@       @       @                                      "@      "@                              "@      �?               @      �?      &@              5@              @       @       @               @      *@      0@                       @      ,@      2@              @                      �?      7@       @      @               @                       @      "@       @              @      1@      @      @       @      �?      .@              *@       @      @                                       @       @                       @      @      @                              @              *@              @                                       @      @                       @      @       @                              @                       @      �?                                              @                                      �?                                              $@              �?               @                      @      �?       @              �?      ,@      @      @       @      �?      "@               @              �?               @                      @      �?       @              �?      (@       @               @      �?      @               @                                                                                               @      �?      @                      @              @      @      6@                      �?      @      &@      @      $@      @      @      (@      .@              @      @      @      @              @                                      �?      "@      @      @              �?      @      @               @       @       @      �?                                                              @      �?                                       @               @                                      @                                      �?       @      @      @              �?      @      �?                       @       @      �?                                                      �?       @       @      @                      @                               @                              @                                                       @                      �?              �?                               @      �?      @       @      6@                      �?      @       @       @      @      @      @      @      (@              @      @      @      @      �?              @                              �?              �?      @               @       @      @                      @       @      @                      �?                                              �?                                      @                                              �?              @                              �?                      @               @       @       @                      @       @      @      @       @      2@                      �?      @       @      �?      �?      @      �?      @      @              @               @       @      @              $@                      �?                      �?      �?      @              @       @                                               @       @       @                              @       @                      �?      �?       @      @              @               @       @�t�bub�     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��<hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         6                   �3@W+��s��?�	           ��@                          �0@t��_�?t           ��@                           @ڂ^b{��?x            `g@                           @��m���?8            @S@                           �?�|гY��?&             I@                            �?ŕ�(�?             5@������������������������       ���8��8�?
             (@������������������������       ��n���?             "@	       
                     �?�#:9$A�?             =@������������������������       �      �?             0@������������������������       ��T�6|��?	             *@                           �?g�WH��?             ;@������������������������       �*�8�G��?             1@������������������������       �p=
ףp�?             $@                           �?�@�!���?@            �[@                           @n�r�X`�?*            �R@                            �?�?             N@������������������������       ��c�MwR�?            �B@������������������������       ��㙢�c�?             7@������������������������       �$߼�x�?             .@                            �?($;=�,�?            �A@������������������������       ��$I�$I�?	             ,@                           @�to@���?             5@������������������������       ��n���?             "@������������������������       �9��8���?             (@       )                     @~� �K��?�           ��@       "                    �?a�AC�?           x�@                           �?FB�ϊ��?�            �l@                           �?����F�?B            @[@������������������������       �\HY���?!            �K@������������������������       ��m(>g�?!             K@        !                   �2@ᣢ���?K            �^@������������������������       �tk�
��?5            �U@������������������������       ����&��?            �A@#       &                    @9�ߧP��?�           @�@$       %                    �?�ֈ/f�?j           Ё@������������������������       �	�«��?�            @s@������������������������       ��ۛ��.�?�            `p@'       (                    �?�x���?             G@������������������������       �
ףp=
�?             .@������������������������       �ؓo
�?             ?@*       1                    @q�'I>�?�            �v@+       .                    �?��|��0�?�            @q@,       -                    @����Z�?|            @g@������������������������       ��ϜRYA�?b            �a@������������������������       �yOҙ��?            �E@/       0                    �?�~�#��?:            �V@������������������������       ���,���?             C@������������������������       ��m��1�?$             J@2       3                    @9�b"p��?5            �V@������������������������       ����Hx�?             B@4       5                    @~*_�#�?              K@������������������������       ���%����?            �@@������������������������       �u���?	             5@7       V                   �7@*����?"           ��@8       G                     @���|hb�?>           ��@9       @                    @�S��?N           0�@:       =                    �?�=�'"�?           `z@;       <                    �?�"$/�?�            �q@������������������������       ���ǆM�?Y            ``@������������������������       ����	"P�?_             c@>       ?                     �?jћ��j�?T            `a@������������������������       �x9/���?"             L@������������������������       �1}|Zu�?2            �T@A       D                    @    p��?B            �@B       C                     �?���Jq�?�            �u@������������������������       ��}�se�?�            `m@������������������������       � |�����?E            �[@E       F                    �?��O1��?l            �d@������������������������       �{[����?/             S@������������������������       �쉵���?=            �V@H       O                    �?9�Ϻ���?�            `x@I       L                   �6@Q����?k            �c@J       K                   �5@n�$��}�?W             `@������������������������       ��x��?>            @X@������������������������       �     �?             @@M       N                     @����S��?             <@������������������������       �)O���?             2@������������������������       �R���Q�?	             $@P       S                   �5@��e�$	�?�             m@Q       R                    @�)O�?S             b@������������������������       �l����?A             [@������������������������       �����K�?             B@T       U                    @��L.N�?2            @V@������������������������       �      �?             L@������������������������       ����%��?            �@@W       f                   �?@�/��u^�?�           ��@X       _                   �8@�ٽC�.�?�           ��@Y       \                    @�.?��V�?�            �m@Z       [                    �?�?@!���?D            @Z@������������������������       �������?%             K@������������������������       �y�j�
�?            �I@]       ^                    @c����O�?\            �`@������������������������       �|�Pk��?E             Y@������������������������       �eTY��&�?            �@@`       c                    @�C�I�?�           �@a       b                    �?7/N�}S�?|           ��@������������������������       ��w�I��?�            �o@������������������������       ���Ly%��?�            Pw@d       e                     �?j�z�a��?{             i@������������������������       ���>4���?C             \@������������������������       �x]��g��?8            @V@g       n                    �?�^���?M            �^@h       k                   �@@�.��T��?+            �P@i       j                    @��*;�?             >@������������������������       �>
ףp=�?             4@������������������������       ��(\����?             $@l       m                    �?n�����?             B@������������������������       ��q�q�?             (@������������������������       ��8��8��?             8@o       r                   �A@/�����?"             L@p       q                    @�3_�?             E@������������������������       ��{�Pk�?             9@������������������������       ��?�0�!�?             1@������������������������       �����>4�?             ,@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       @@     �W@     �u@     �A@      R@      4@      R@     ��@     ��@     @P@     �U@     �a@     ��@     �{@      .@     @P@     �H@      a@      L@      f@      8@     �[@      @      "@              @     �s@      p@      $@      4@      F@     �l@     �^@              &@      @     �E@      $@      :@      @      @              �?                      T@      A@                              :@      "@                               @              *@      @      @                                      .@      7@                              *@      @                                              (@      @      �?                                      $@      "@                              &@      @                                              @                                                       @      @                              @                                                      @                                                      @      @                              �?                                                       @                                                      @                                      @                                                      @      @      �?                                       @      @                              @      @                                              @              �?                                      �?      @                              @      �?                                              @      @                                              �?      @                                      @                                              �?               @                                      @      ,@                               @      @                                              �?                                                      @      @                               @       @                                                               @                                              @                                      �?                                              *@              @              �?                     @P@      &@                              *@       @                               @              @              @                                      F@      "@                              (@                                                       @              @                                     �C@      @                              &@                                                                      @                                      9@      �?                               @                                                       @                                                      ,@      @                              @                                                      @                                                      @      @                              �?                                                      @                              �?                      5@       @                              �?       @                               @              @                                                       @                                                                               @               @                              �?                      *@       @                              �?       @                                              �?                                                      @      �?                              �?      �?                                              �?                              �?                       @      �?                                      �?                                             �b@      5@     @Z@      @       @              @     �m@     �k@      $@      4@      F@     `i@     @\@              &@      @     �D@      $@     �Y@      0@      J@      @      @              @     `j@     �d@      @      @      @@     �a@      Q@              @      �?      5@      @      D@      @      .@      �?                              D@      A@      �?      @      ,@      F@      7@               @              @      @      8@       @      @                                      <@      ,@      �?      �?      @      6@      @                              @              &@               @                                      ,@      @      �?              @      ,@      @                                              *@       @      @                                      ,@      @              �?               @      @                              @              0@       @      $@      �?                              (@      4@               @      &@      6@      1@               @              @      @       @               @                                      @      2@              �?       @      6@      &@                               @       @       @       @       @      �?                              @       @              �?      @              @               @               @      �?      O@      (@     �B@       @      @              @     `e@     �`@      @      @      2@     �X@     �F@              @      �?      ,@      @     �I@      (@      A@       @                      @     �d@     �^@      @      @      0@      V@      F@              @      �?      *@      @      3@      @      *@       @                      @     �X@      R@      �?      �?      @      K@      9@                              @              @@       @      5@                              �?      Q@      I@      @      @      "@      A@      3@              @      �?      @      @      &@              @              @              �?      @      $@                       @      $@      �?                              �?              @               @                                      @                                      @                                                      @              �?              @              �?      �?      $@                       @      @      �?                              �?             �H@      @     �J@              @              �?      <@      L@      @      *@      (@     �N@     �F@              @      @      4@      @     �C@      @      ?@              @                      3@      E@      @      $@      "@      J@      A@               @      @      2@      �?      4@      @      7@              @                      "@      9@      @       @      @      A@      :@               @      @      2@      �?      1@      @      ,@              @                      "@      3@      �?       @      @      =@      3@               @      �?      (@              @              "@                                              @       @              �?      @      @                      @      @      �?      3@               @              �?                      $@      1@       @       @      @      2@       @                                              (@               @                                      �?      @                      @      &@      @                                              @              @              �?                      "@      *@       @       @       @      @      @                                              $@              6@                              �?      "@      ,@              @      @      "@      &@              @               @       @       @              2@                                      @      @               @       @      �?       @                                               @              @                              �?      @       @              �?      �?       @      "@              @               @       @      @              @                              �?      @       @              �?              @       @              �?                              @                                                                                      �?      @      @              @               @       @     0t@     �Q@      n@      @@     �O@      4@     @P@     �j@     �s@     �K@     �P@     @X@     �w@     �s@      .@      K@      F@     @W@      G@      i@      1@     ``@      .@      7@      $@      5@     �b@      i@      1@      <@     �F@      k@      c@       @      5@      2@      F@      &@     �a@      @      W@      @      ,@              (@     @]@     �d@       @      9@      :@      c@      Y@              0@      &@      A@      @     �K@       @     �O@       @      @               @      @@     �P@      @      1@      $@     @R@     �J@              @      @      0@              F@             �D@      �?      @              @      2@     �A@      �?      1@      @      L@      =@              @      @      &@              5@              1@              @              �?      *@      2@              @      @      A@      @              @               @              7@              8@      �?      �?              @      @      1@      �?      &@      @      6@      6@              @      @      "@              &@       @      6@      �?      �?              �?      ,@      @@      @              @      1@      8@                              @              @       @      @      �?      �?              �?      @      *@                       @       @      @                              @              @              0@                                      "@      3@      @              �?      "@      3@                                              V@      @      =@      @      @              @     @U@     @X@      �?       @      0@     �S@     �G@              "@       @      2@      @      J@       @      2@       @                      @     @P@     �Q@      �?      @      (@      M@      A@              @      @      &@       @      >@              1@                                      C@      L@      �?      @      $@      B@      :@              @      @      @       @      6@       @      �?       @                      @      ;@      ,@              @       @      6@       @                              @              B@      @      &@      @      @              �?      4@      ;@              �?      @      5@      *@              @      @      @      @      2@              @                                      *@      5@              �?      �?      &@      @              �?               @              2@      @      @      @      @              �?      @      @                      @      $@      $@              @      @      @      @     �L@      $@     �C@       @      "@      $@      "@      A@     �B@      "@      @      3@     @P@      J@       @      @      @      $@      @      3@      �?      1@      �?      @      @      �?      5@      1@       @      @      @      A@      6@      �?       @      @      @              &@              0@      �?      �?      @      �?      4@      &@       @       @      �?      ?@      5@               @       @      @              "@              0@              �?      �?      �?      .@      $@       @       @      �?      4@      *@               @      �?      @               @                      �?               @              @      �?                              &@       @                      �?      �?               @      �?      �?               @                      �?      @              �?       @      @      �?      �?              �?                       @      �?      �?              �?                               @                              @      �?      �?                                                                      �?                      �?      @              �?       @                                      �?                      C@      "@      6@      @      @      @       @      *@      4@      @              0@      ?@      >@      �?      @      @      @      @      @@      @      .@      @      @      @      @      @      @       @              ,@      4@      2@                      @      @      �?      0@      @      ,@              @      @      @      @      @       @              &@      2@      ,@                      @      @              0@      �?      �?      @                               @       @                      @       @      @                                      �?      @      @      @      @      @      @      @      @      *@      @               @      &@      (@      �?      @      �?       @      @      @      �?                       @       @              @      (@      @              �?      &@      @              @      �?      �?       @               @      @      @      �?       @      @      �?      �?                      �?               @      �?                      �?       @     �^@     �J@     @[@      1@      D@      $@      F@      P@     @]@      C@     �C@      J@      d@     �d@      *@     �@@      :@     �H@     �A@      \@      J@     �Y@      *@      <@      @      D@     �O@     �[@      9@     �@@      E@     @c@     `c@      @      <@      7@     �G@      ;@      :@      @      >@       @      @              @      7@      <@      @      @      @      7@      J@      �?      @       @      (@      @       @      @      "@       @                      @      1@      0@       @                      *@      7@               @              @              @      �?      @                               @      $@      "@       @                       @       @               @                              @       @       @       @                      @      @      @                              @      .@                              @              2@      @      5@              @               @      @      (@      @      @      @      $@      =@      �?       @       @      @      @      0@      @      3@              @               @      �?       @       @      @      @      @      8@                       @       @      @       @               @              �?                      @      @      �?                      @      @      �?       @              @             �U@     �F@     @R@      &@      8@      @     �@@      D@     �T@      4@      <@      C@     ``@     �Y@      @      8@      5@     �A@      8@      T@      9@      L@      "@      6@      @      8@      8@     �N@      (@      4@      A@     �U@     �S@       @      5@      2@      <@      4@     �C@      1@      4@      @      @              $@      *@      C@      �?      @      @      C@      @@              @      @      $@      @     �D@       @      B@      @      .@      @      ,@      &@      7@      &@      0@      =@     �H@      G@       @      ,@      &@      2@      0@      @      4@      1@       @       @              "@      0@      6@       @       @      @      F@      9@      �?      @      @      @      @      @      @      $@      �?       @                      *@      1@      @      @       @      <@      ,@                       @       @      @      @      0@      @      �?                      "@      @      @      @      �?       @      0@      &@      �?      @      �?      @      �?      &@      �?      @      @      (@      @      @      �?      @      *@      @      $@      @      &@      "@      @      @       @       @       @              �?      @      (@       @      @                      @      @      @              @       @       @      @              @      �?                      @      @       @                              @      @       @              @              �?       @              �?      �?                      @       @                                      @      @                      @              �?                                                              @       @                                               @                                       @              �?      �?              �?      �?      @              @                      @      �?      @                       @      �?      �?              @      �?              �?              @              @                                                               @                                                              �?       @                                      @      �?      @                      @      �?      �?              @      "@      �?      @                      �?      �?      �?      @      @              @      @      @      �?      @               @      �?       @              @                      �?              �?      @      @              @      @      @      �?      �?               @      �?                                                              �?      @      @                      @      @      �?      �?               @               @              @                      �?                      �?                      @       @      �?                                      �?      @      �?      �?                              �?                                                       @               @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�"�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         8                   �1@J�j5��?�	           ��@                           �?0$ډ�/�?�           ��@                           @�b"�i�?�             q@                           �?��˶�?@            �Z@                           �?��_R�?#            �N@                          �0@�8��8��?             8@������������������������       ���1G���?             *@������������������������       �Y�����?             &@	       
                    �?$��0�?            �B@������������������������       �     @�?             0@������������������������       �>F?�!��?             5@                           �?��JÝ�?             G@                          �0@X��H��?             A@������������������������       ��C��2(�?             &@������������������������       ����Q��?             7@������������������������       ��8��8��?             (@                            �?�M�����?a            �d@                           �?2q�{��?             E@                           @����3��?             :@������������������������       �b�r���?             .@������������������������       ���ˠ�?             &@������������������������       �      �?             0@                           �?�I�p�?G            @_@                           @`����?/            �U@������������������������       �Uat�X��?            �J@������������������������       ��hJ,��?             A@                          �0@��d���?             C@������������������������       ��C��2(�?             &@������������������������       �~X�<��?             ;@       +                   �0@���D--�?�            v@       &                     �?C�8����?Q            �`@        #                    @�~$7q�?)             O@!       "                     �?�<J�L�?            �B@������������������������       ��������?             1@������������������������       ��Q����?
             4@$       %                    @^K�=��?             9@������������������������       ��'}�'}�?             .@������������������������       ����(\��?             $@'       (                    �?�7�V�?(            �Q@������������������������       �،A��_�?
             1@)       *                    �?N��:��?             K@������������������������       �VUUUUU�?             8@������������������������       ���ĳ���?             >@,       1                     �?��ɰ'�?�            �k@-       .                    �?�2�tk~�?'            �O@������������������������       �x�5?,�?             2@/       0                    @�k��?            �F@������������������������       �/�E���?             ?@������������������������       �d}h���?             ,@2       5                    @C>��s�?g            �c@3       4                    @hֵ!�?2            �S@������������������������       �j�'�ſ�?%             M@������������������������       ���[r��?             5@6       7                    �?�7���?5            �S@������������������������       ���pX��?             ?@������������������������       ��������?             �G@9       V                   �6@ ��v���?           ��@:       G                     @��P�4�?~           �@;       @                    �?��1/>��?)           h�@<       ?                    @�v_�vz�?�            Px@=       >                     �?�0���|�?�            �w@������������������������       ���>�?~            �h@������������������������       ����5�?o            �f@������������������������       ��q�q�?             (@A       D                    �?y~����?5           ��@B       C                   �3@l�w�T��?           �|@������������������������       �ߞ�����?�            @j@������������������������       �Z�J�R�?�            �n@E       F                   �4@]R�0��?           �|@������������������������       �e�/�F�?�            �r@������������������������       ����I�?]            �c@H       O                    @f�Fqn��?U           �@I       L                   �4@������?           �y@J       K                   �3@�����?�            �p@������������������������       �8���V��?r            `e@������������������������       �E��F��?=            �W@M       N                    @�$���?_            �b@������������������������       ����i�V�?;             V@������������������������       ���2Tv�?$             N@P       S                    �?r]�&�_�?G            �`@Q       R                    @�����?!             O@������������������������       �B�����?             :@������������������������       ��E��ӭ�?             B@T       U                    @&a�u�|�?&            �Q@������������������������       �{�G�z�?             D@������������������������       ��>�\��?             ?@W       d                    �?T�˹�c�?�           h�@X       ]                    �?�SHͰ��?�           ؆@Y       \                   �>@NR'��?l            �e@Z       [                     �?����+��?a            `c@������������������������       ��&V���?            �H@������������������������       �6y��D�?G            �Z@������������������������       �ZZZZZZ�?             1@^       a                   �8@�X2Q9��?h           x�@_       `                    @�0���?s             g@������������������������       �Pdl<)��?b            �c@������������������������       ��@�Y��?             =@b       c                     �?�o'���?�            `w@������������������������       �P�k|_=�?L            �^@������������������������       ����c��?�            `o@e       l                     �?ܦ5��?�           ��@f       i                   �>@|d���?�            `i@g       h                    @������?y             g@������������������������       ��9��(��?M            �^@������������������������       ��!͎�?,            �O@j       k                    @0�����?             2@������������������������       �R���Q�?             $@������������������������       �      �?              @m       p                    @C�8
�?,           @@n       o                    @v��[��?�            `n@������������������������       �G�
�5�?_             e@������������������������       ��lJ�Y �?/            �R@q       r                   �>@<��S|��?�            p@������������������������       ��WXH��?�            �m@������������������������       ���Hx��?
             2@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       p|@      P@     �u@      G@     @V@      @@     �R@     ��@      �@      N@     �R@     �g@     ��@     {@       @     @Q@      K@     @]@     �O@     @U@       @      ;@              @               @     �k@      `@      @      @      0@      X@      :@               @               @       @      A@              @              @              �?     �]@     �M@      �?       @      @     �A@      @                              �?       @      7@              @              @              �?     �@@      .@      �?       @      @      3@      �?                                       @      .@               @                                      7@       @      �?       @      �?       @      �?                                              "@               @                                      @      @      �?              �?                                                               @               @                                      @      @                                                                                      @                                                      �?      �?      �?              �?                                                              @                                                      0@      @               @               @      �?                                              �?                                                      $@                                      @      �?                                              @                                                      @      @               @              @                                                       @               @              @              �?      $@      @                       @      &@                                               @       @                              @                      @      @                              "@                                               @      @                                                              @                              @                                                      @                              @                      @      @                              @                                               @                       @                              �?      @                               @       @                                                      &@              @                                     �U@      F@                      @      0@      @                              �?              @                                                      0@      2@                      �?      �?                                                      @                                                      $@      $@                      �?      �?                                                      @                                                      @      @                                                                                                                                              @      @                      �?      �?                                                       @                                                      @       @                                                                                      @              @                                     �Q@      :@                       @      .@      @                              �?               @                                                     �J@      5@                              $@      �?                                              �?                                                      A@      "@                              "@                                                      �?                                                      3@      (@                              �?      �?                                              @              @                                      1@      @                       @      @       @                              �?                                                                      $@                                      �?                                                      @              @                                      @      @                       @      @       @                              �?             �I@       @      4@              �?              �?     �Y@     �Q@       @       @      $@     �N@      6@               @              @              :@              �?                                      N@      9@                      �?      .@      @                                              &@                                                      5@      4@                      �?       @      �?                                              @                                                      $@      0@                              @      �?                                              �?                                                      @      @                              @      �?                                               @                                                      @      "@                              @                                                       @                                                      &@      @                      �?      �?                                                       @                                                      "@      @                              �?                                                      @                                                       @      �?                      �?                                                              .@              �?                                     �C@      @                              @      @                                               @              �?                                      @       @                                                                                      @                                                     �@@      @                              @      @                                              @                                                      *@      @                              @                                                      @                                                      4@                                      @      @                                              9@       @      3@              �?              �?      E@     �F@       @       @      "@      G@      1@               @              @              "@       @                                              "@      *@                              8@      @                               @              @                                                      @      �?                              &@                                                      @       @                                              @      (@                              *@      @                               @              @                                                      @      "@                              @      @                              �?              �?       @                                                      @                              @                                      �?              0@              3@              �?              �?     �@@      @@       @       @      "@      6@      *@               @              @              @              $@              �?              �?      6@      3@               @      @      (@      @                                              @              $@              �?              �?      0@      @               @      @      $@      @                                              �?                                                      @      (@                               @                                                      &@              "@                                      &@      *@       @              @      $@      "@               @              @              @              @                                      $@      $@                               @      �?                                              @              @                                      �?      @       @              @       @       @               @              @              w@      O@     �s@      G@     @U@      @@     @R@     Pu@     0|@     �L@     �Q@     �e@     @@     py@       @     �P@      K@     @[@     �N@     �j@      .@     �d@      1@      8@      @     �A@     �p@     �s@      4@      =@     @R@     �s@     `l@             �A@      0@      P@      6@      e@      @     @\@      @      &@              9@     `i@      n@      (@      7@      K@     �i@     `d@              6@      @     �B@      (@      N@       @     �F@      �?      �?              @     �A@      F@      @      (@      6@     �P@      G@              &@      @      2@      $@     �M@       @     �E@      �?      �?              @     �A@     �E@      @      (@      6@     �P@      C@              &@      @      2@      $@      ;@       @      1@      �?      �?               @       @      7@      @      @      1@     �E@      8@              @      @      &@      @      @@              :@                              @      ;@      4@      �?       @      @      8@      ,@               @              @      @      �?               @                                              �?                                       @                                             @[@      @      Q@      @      $@              2@      e@     �h@      @      &@      @@      a@     @]@              &@      @      3@       @     �J@       @     �@@              �?              @     @S@     �]@      @      @      &@      T@      K@              �?       @      "@              0@              6@                                      I@      F@      @      �?      @      A@      :@                              @             �B@       @      &@              �?              @      ;@     �R@      �?      @      @      G@      <@              �?       @      @              L@      �?     �A@      @      "@              *@     �V@     �S@      �?      @      5@     �L@     �O@              $@       @      $@       @      A@              1@      @      @              @     �Q@     �P@      �?      @      *@     �B@      A@              "@       @      @      �?      6@      �?      2@              @              "@      5@      (@              @       @      4@      =@              �?              @      �?      F@      $@      J@      (@      *@      @      $@     �N@     �Q@       @      @      3@     @\@      P@              *@      "@      ;@      $@     �B@      $@      B@       @      $@      @      $@      =@     �N@      @      @      0@     �U@     �G@              $@      "@      3@      "@     �A@      @      4@      @      @      �?              4@      D@       @      @      (@     �N@     �@@              @      �?      (@      @      5@      �?       @      @      @                      ,@      ;@      �?      �?      @     �C@      8@              @      �?      &@      @      ,@      @      (@               @      �?              @      *@      �?       @      @      6@      "@                              �?       @       @      @      0@      @      @      @      $@      "@      5@      @       @      @      9@      ,@              @       @      @      @       @      @      @              @      �?               @      2@      @      �?              .@      &@              @       @      @       @               @      $@      @               @      $@      �?      @       @      �?      @      $@      @                      @       @      �?      @              0@      @      @                      @@      $@      �?      �?      @      ;@      1@              @               @      �?       @              @                                      0@      @      �?      �?      �?      *@      (@              @              @               @              @                                      ,@                                      @      �?                               @                              �?                                       @      @      �?      �?      �?      $@      &@              @              @              @              &@      @      @                      0@      @                       @      ,@      @                              @      �?      @              &@      @                               @      @                       @      $@      �?                               @      �?       @                              @                      ,@      @                              @      @                              �?             �c@     �G@     @c@      =@     �N@      <@      C@     @S@     `a@     �B@      E@      Y@     �f@     �f@       @      @@      C@     �F@     �C@     �T@      8@     �W@      (@     �C@      3@      7@      3@      I@      4@      ;@      P@      R@      S@      @      3@      >@      =@      ;@      A@      @      5@       @      @      @      @      @      $@      @      @      @      2@      1@       @      @      @      .@      @     �@@      @      4@      �?      @       @      @      @      "@      @      @      @      (@      1@       @      @       @      .@      @      $@                              �?               @      @      @      @      �?       @      @      @                      �?      &@              7@      @      4@      �?      @       @      �?       @      @       @       @      @      "@      (@       @      @      �?      @      @      �?              �?      �?       @       @      �?              �?              �?              @                              �?                      H@      1@     @R@      $@     �@@      .@      3@      *@      D@      ,@      7@     �L@      K@     �M@      @      0@      ;@      ,@      8@      9@      "@      :@       @      @      �?      @      @      3@       @      (@      5@       @      =@               @       @      @       @      .@      @      7@       @      @      �?      @      @      3@       @      "@      4@      @      :@               @      @      @      �?      $@       @      @                                      �?                      @      �?      �?      @                       @       @      �?      7@       @     �G@       @      <@      ,@      0@       @      5@      (@      &@      B@      G@      >@      @      ,@      3@       @      6@      @      @      6@      @      &@      @      @              $@      �?      @      @      .@      @               @      @       @      @      1@      @      9@      @      1@       @      &@       @      &@      &@      @      @@      ?@      8@      @      @      (@      @      1@     �R@      7@      N@      1@      6@      "@      .@      M@     @V@      1@      .@      B@     �[@      Z@      @      *@       @      0@      (@      0@       @      *@              �?      @       @      2@      6@      @      @      $@      B@     �G@              "@      �?      @       @      0@       @      "@              �?      @       @      2@      5@      @      @      @      B@     �E@               @      �?      @       @      *@       @      @              �?      @       @      @      $@       @      @      @      <@      9@              @      �?      @      �?      @              @                                      &@      &@      �?              �?       @      2@              @              �?      �?                      @                                              �?      �?              @              @              �?              @                               @                                                                      @              �?              �?              @                               @                                              �?      �?              �?              @                                             �M@      5@     �G@      1@      5@      @      @      D@     �P@      *@      &@      :@     �R@     �L@      @      @      @      "@      $@      B@      &@      0@       @      3@      @      �?      *@      7@       @      �?      0@      A@      B@              @      @      @      @      2@      @      ,@       @      ,@      @              (@      ,@      @              &@      1@      <@              @      @      @      @      2@      @       @              @              �?      �?      "@      �?      �?      @      1@       @              �?              �?              7@      $@      ?@      "@       @              @      ;@      F@      @      $@      $@     �D@      5@      @              @      @      @      7@      $@      6@      "@       @              @      ;@      E@      @      $@      "@      D@      1@      @              @      @      @                      "@                                               @                      �?      �?      @                                      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�,thG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKuhnh4h7K ��h9��R�(KKu��hu�B�         8                   �2@׊�
���?�	           ��@                           @f;��<��?{           ؏@                            @��"��X�?;           �~@                            �?,�6���?�            �s@                           �?+U�߼��?d             e@                           @(N:!���?,            �Q@������������������������       �o� 6 �?$            �M@������������������������       �j�V���?             &@	       
                   �0@������?8            �X@������������������������       �$��Z=;�?             6@������������������������       �T��g��?,            @S@                           �?u���?\            `b@                          �0@^�t�C��?,            �R@������������������������       �X�<ݚ�?
             2@������������������������       ��W5����?"            �L@                          �1@��a�2��?0             R@������������������������       ��ח���?            �B@������������������������       ��0f߻�?            �A@                           �?��/��?{            �e@                           �?��Β��?3            @R@                          �1@�?9Ҫ~�?"            �G@������������������������       ����Q��?             4@������������������������       ���F�� �?             ;@                           @���B���?             :@������������������������       ���
ц��?
             *@������������������������       �;�;��?             *@                          �0@�!���?H            �Y@������������������������       ��q-��?
             *@                          �1@��x��?>            @V@������������������������       �<�bj*R�?             �G@������������������������       ��Sy'��?             E@        /                    �?���*�d�?@           ��@!       (                    @�{D (�?�            �k@"       %                     @��Z�L�?H            �^@#       $                   �1@R�8	��?.             S@������������������������       ���8���?             H@������������������������       �T�r
^N�?             <@&       '                    �?����?             G@������������������������       ��W��H��?             1@������������������������       �x�-�?             =@)       ,                     �?���&S�?@             Y@*       +                    �?h���I�?             7@������������������������       �B{	�%��?             "@������������������������       �^N��)x�?	             ,@-       .                    @XӨ*��?0            @S@������������������������       �h��|?5�?             I@������������������������       ��.sxQ��?             ;@0       1                    �?�������?�             s@������������������������       �S��d�?             >@2       5                     �?�<��}�?�            @q@3       4                   �0@��L��?,            �Q@������������������������       �;�;��?             *@������������������������       ��,!�N�?$            �L@6       7                    @�|�T{�?~            �i@������������������������       ������?^            �b@������������������������       �E��ůs�?             �K@9       X                    �?��7����?           ��@:       I                    �?}��'�?7           4�@;       B                     �?��J��?T           x�@<       ?                    �?��|���?^             c@=       >                    �?��92���?%             M@������������������������       ���(\���?             4@������������������������       �"P7��?             C@@       A                   �:@������?9            �W@������������������������       ����?.            �S@������������������������       ��X�%��?             .@C       F                     @#��@!��?�            pw@D       E                   �8@ۤm�Z�?g            �c@������������������������       ��䘉�B�?K            �]@������������������������       ��(\����?             D@G       H                    @�������?�             k@������������������������       �R�ߦ5�?<            �V@������������������������       �����j��?S            �_@J       Q                     @���v�W�?�           ��@K       N                   �>@-�zΟ �?           �|@L       M                    �?��JX(��?           �z@������������������������       �c��:��?q            �h@������������������������       ��^�sK��?�            �l@O       P                    �?ڣ����?            �@@������������������������       �ƵHPS!�?             *@������������������������       ����Q��?             4@R       U                    �?$u
?l�?�            @s@S       T                    �?�d�����?2             S@������������������������       �     ��?
             0@������������������������       ��&���?(             N@V       W                   �4@Z0Rb�?�             m@������������������������       ���*�R��?$            �K@������������������������       ���D� f�?s             f@Y       f                    �?��m���?�           �@Z       _                    �?��*��?�           ��@[       ^                   �;@3��-��?�            �n@\       ]                   �4@�,�'UJ�?�            �l@������������������������       �҇����?8            �U@������������������������       ���;����?\             b@������������������������       ��������?	             .@`       c                   �8@]D#�,�?>           �@a       b                    @L?�Z�j�?�            �u@������������������������       ���~UZ��?+            @Q@������������������������       ���N�?�            �q@d       e                    �?$� ����?a            �c@������������������������       �      �?
             0@������������������������       �Ԭ▾�?W            �a@g       n                   �9@L��	]��?           ��@h       k                    �?�_���?�           0�@i       j                    @�ke���?s             h@������������������������       ��=��/�?            �D@������������������������       �(�@݈g�?W             c@l       m                   �8@��T#s�?           P|@������������������������       ��_@��z�?           �y@������������������������       ��������?             D@o       r                    @�.WL��?y            `i@p       q                   �;@xJLCe��?3            �T@������������������������       ���pX��?             ?@������������������������       �o_Y�K�?#             J@s       t                   �>@v���� �?F             ^@������������������������       ���\ju��?6            @V@������������������������       ������?             ?@�t�bh�h4h7K ��h9��R�(KKuKK��h��BxE        @      T@     �t@     �A@      S@      A@     �U@     0�@     x�@      Q@     �Q@     @d@     H�@     �{@      &@     �P@     �F@      `@     �J@     �`@      &@     �N@      @      @              &@     Pp@      k@      "@      "@      9@     @f@      Q@              @      @      0@      @     @R@      @      @@      @      @              @     �S@     �Z@      @       @      0@     �W@      D@              �?      �?      (@      @     �G@              3@               @               @      R@     @S@      @      @      "@     �J@      .@              �?              @      @      <@              "@                                      <@     �C@      @      @      @      C@      @              �?              @      @      .@               @                                      .@      1@              @      �?      *@      @                              �?              ,@               @                                      *@      "@              @      �?      *@      @                              �?              �?                                                       @       @                                                                                      *@              @                                      *@      6@      @              @      9@      @              �?               @      @       @                                                      @      (@                               @      �?                                              &@              @                                       @      $@      @              @      7@      @              �?               @      @      3@              $@               @               @      F@      C@      �?      @      @      .@       @                              �?               @              @                                      >@      5@               @      @      @      @                                                                                                       @      $@                                                                                       @              @                                      6@      &@               @      @      @      @                                              &@              @               @               @      ,@      1@      �?      �?      �?      (@      @                              �?               @              @               @              �?      $@      @      �?      �?      �?       @      �?                              �?              @               @                              �?      @      *@                              $@       @                                              :@      @      *@      @      @              �?      @      =@       @       @      @      E@      9@                      �?       @      �?      @              @                              �?      @      .@       @              @      8@      $@                              @              @              @                              �?       @       @       @              @      $@      "@                              @               @               @                                              @       @               @      @      @                                               @              �?                              �?       @      @                       @      @      @                              @              @                                                      �?      @                              ,@      �?                                              �?                                                      �?      �?                              "@      �?                                               @                                                              @                              @                                                      3@      @      $@      @      @                      @      ,@               @      @      2@      .@                      �?      @      �?      @      �?                                               @      �?                                       @                                              (@      @      $@      @      @                       @      *@               @      @      2@      *@                      �?      @      �?      @              @              @                       @      @                      @      (@       @                      �?      @              @      @      @      @                                      $@               @              @      @                              �?      �?      N@      @      =@                               @     �f@     �[@       @      �?      "@     �T@      <@              @       @      @      �?      4@       @      6@                              @     �W@      B@              �?      @      <@      @              �?               @              2@       @      4@                                      E@      1@              �?      @      2@      �?                                              @       @      @                                      A@      .@              �?      �?      ,@                                                      @       @      @                                      6@      (@              �?      �?      @                                                      @                                                      (@      @                              $@                                                      (@              1@                                       @       @                       @      @      �?                                              �?              "@                                      @      �?                              �?                                                      &@               @                                      @      �?                       @      @      �?                                               @               @                              @     �J@      3@                      �?      $@      @              �?               @              �?                                              @       @      @                      �?      @       @                                                                                                      @                              �?      �?                                                      �?                                              @      �?      @                              @       @                                              �?               @                              �?     �F@      .@                              @      @              �?               @                                                              �?     �A@      "@                               @      @                                              �?               @                                      $@      @                              @      �?              �?               @              D@      @      @                              @     �U@     �R@       @              @     �K@      5@               @       @       @      �?       @                                                      �?       @                              @      @                                              @@      @      @                              @     �U@     �P@       @              @     �H@      ,@               @       @       @      �?      @      �?                                      �?      0@      <@                              (@      @                       @      �?               @                                                      @      @                                                                                      @      �?                                      �?      &@      6@                              (@      @                       @      �?              ;@      @      @                              @     �Q@      C@       @              @     �B@      $@               @              �?      �?      7@      @      @                              @      M@      5@                      @      9@      @                              �?      �?      @              @                                      (@      1@       @                      (@      @               @                             �v@     @Q@     �p@      @@     �Q@      A@      S@     p@     pw@     �M@     �N@      a@     p{@     @w@      &@     �O@      E@     @\@     �G@      f@     �C@     @a@      0@      E@      :@      @@      P@     @_@      3@      ?@      R@     `e@      f@       @     �C@      =@     �L@      @@     @R@      &@      K@       @      ,@      �?      "@      D@     �Q@      @      $@      6@     @V@      Q@      @      .@      *@      2@      $@      1@      @      4@      �?       @               @      @      7@      �?      @      @     �B@      0@              @      @      "@               @      �?      @                                      �?      (@      �?              @      0@      @               @      @      �?              @              �?                                              $@                              @                              @                      @      �?       @                                      �?       @      �?              @      *@      @               @              �?              "@       @      1@      �?       @               @      @      &@              @       @      5@      "@               @               @              @              1@      �?       @              �?      @      "@              @       @      5@       @               @              @              @       @                                      �?               @                                      �?                              @              L@       @      A@      �?      (@      �?      @      A@      H@      @      @      1@      J@      J@      @      &@      $@      "@      $@      =@      @      (@               @               @      4@      ,@      �?      @      @      7@      8@              @      @       @      @      =@              "@                              �?      3@      $@      �?      @      @      6@      (@              @               @       @              @      @               @              �?      �?      @              �?      �?      �?      (@                      @              @      ;@      �?      6@      �?      $@      �?      @      ,@      A@       @       @      *@      =@      <@      @      @      @      @      @      1@      �?      "@              @                      @      "@       @      �?      @      0@      (@       @      @              @              $@              *@      �?      @      �?      @      $@      9@              �?      "@      *@      0@      �?              @      @      @     �Y@      <@      U@      ,@      <@      9@      7@      8@      K@      .@      5@      I@     �T@     @[@      @      8@      0@     �C@      6@      P@       @      L@      @      (@      @      *@      4@      ?@       @      1@      ?@     �K@      P@      �?      2@      &@      ;@      .@      P@       @     �I@      @      &@      �?      &@      4@      >@      @      ,@      8@     �K@      P@      �?      0@      @      8@      ,@      @@      @      (@      �?      "@      �?      @      "@      3@      �?      @      $@      A@      :@              @      @      @      (@      @@      @     �C@      @       @              @      &@      &@      @       @      ,@      5@      C@      �?      (@       @      3@       @                      @              �?       @       @              �?      �?      @      @                               @      @      @      �?                      @              �?               @                              @       @                                               @                               @                       @                      �?      �?              @                               @      @      �?      �?     �C@      4@      <@      $@      0@      6@      $@      @      7@      @      @      3@      ;@     �F@      @      @      @      (@      @      ,@      @      "@              @              �?      @      @      @              @      @      $@               @      �?      @      @                                                              �?      �?      @              �?              @               @      �?              �?      ,@      @      "@              @              �?      @       @                      @      @      @                              @       @      9@      1@      3@      $@      &@      6@      "@              4@      @      @      (@      4@     �A@      @      @      @      "@      @      ,@      @      @                                              @                      @      $@      "@                               @              &@      ,@      .@      $@      &@      6@      "@              1@      @      @       @      $@      :@      @      @      @      �?      @     �g@      >@     �`@      0@      =@       @      F@      h@     @o@      D@      >@     @P@     �p@     `h@      @      8@      *@      L@      .@     �W@      $@      F@      @       @               @      ^@     �b@      &@      6@      4@      `@     �X@              &@      �?      4@      @      5@      @      .@              �?               @      =@     �P@      �?      @      @      L@     �A@              @              �?              4@      @      .@              �?                      =@     @P@      �?      @      @     �I@      A@                              �?              "@              @                                      1@      1@                       @      4@      1@                                              &@      @      &@              �?                      (@      H@      �?      @      @      ?@      1@                              �?              �?       @                                       @              �?                              @      �?              @                             @R@      @      =@      @      @              @     �V@     �T@      $@      0@      .@     @R@     �O@               @      �?      3@      @     �L@              2@      @                      @     �Q@      Q@      @      @      @      I@      C@              �?      �?      2@              ,@              @      �?                              @      ,@                      @      .@      @                              @             �E@              *@       @                      @      P@      K@      @      @       @     �A@      ?@              �?      �?      .@              0@      @      &@       @      @                      5@      ,@      @      "@      "@      7@      9@              @              �?      @              �?      �?               @                       @      �?                              @                                                      0@      @      $@       @      @                      *@      *@      @      "@      "@      4@      9@              @              �?      @     �W@      4@     @V@      &@      5@       @      B@     @R@     �Y@      =@       @     �F@     `a@     @X@      @      *@      (@      B@      (@      V@      (@     @R@      $@      &@       @      9@      Q@     @V@      (@      @      ?@     �[@     �M@              &@      @      4@      &@      0@      �?      ,@              �?       @      "@      ;@     �A@      @      �?      (@      ;@      8@              @      @      @       @      @      �?      @                       @              �?      "@                              "@      @               @               @              &@               @              �?              "@      :@      :@      @      �?      (@      2@      4@              @      @      �?       @      R@      &@     �M@      $@      $@              0@     �D@      K@      "@      @      3@     �T@     �A@              @       @      1@      @      R@       @     �K@      $@      $@              ,@      C@      H@      "@      @      2@      Q@      ?@              @       @      1@      @              @      @                               @      @      @               @      �?      .@      @                                              @       @      0@      �?      $@      @      &@      @      *@      1@      �?      ,@      =@      C@      @       @      @      0@      �?       @      @      @      �?      @      @              �?      �?       @      �?      "@      (@      7@       @              �?      @              �?      @      �?              @                      �?                              �?       @      (@                                              �?      @       @      �?              @                      �?       @      �?       @      @      &@       @              �?      @              @      �?      *@              @       @      &@      @      (@      "@              @      1@      .@      �?       @      @      &@      �?      @      �?      @               @       @      &@       @      "@      @               @      0@      &@      �?       @      @      &@      �?                      "@              @                       @      @      @              @      �?      @                                        �t�bub��     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ唞mhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmK{hnh4h7K ��h9��R�(KK{��hu�B�         @                     @^jӚ�?�	           ��@       !                   �5@�[N@Y�?�           ��@                           �?��G/"�?�           �@                            �?w��1D�?�            �y@                           �?�WZ�?�            �k@                           �?X���?.            @S@������������������������       ��Kh/���?             B@������������������������       �����#E�?            �D@	       
                    �?{�	)r��?W            �a@������������������������       �)栤�?%             O@������������������������       �)��I�?2            @T@                           @��V����?x            �g@                           @�b���?k            �d@������������������������       �P�n#��?X             a@������������������������       ���X��?             <@                           �?�g���u�?             ;@������������������������       �*�8�G��?             1@������������������������       ����(\��?             $@                           �?����]�?�           ��@                          �2@ڠ�Y��?c           H�@                          �0@O֦(�9�?�            0t@������������������������       ���y�T��?)            �R@������������������������       �X�'����?�             o@                            �?cV�Q��?�            `p@������������������������       � @���?l            �e@������������������������       ��2(&��?;             V@                           @�g+�f�?U            �@                           @l�h���?           pz@������������������������       �֔��@v�?�            �l@������������������������       �lS�$�?w             h@                           �2@X!�1�?Q            @^@������������������������       ��3��\{�?!            �H@������������������������       �<ݚ�?0             R@"       1                    �?&���?           $�@#       *                     �?���nN<�?H           �~@$       '                   �7@*ua��?�            Px@%       &                   �6@��>9��?V            �`@������������������������       ��d��0�?&             N@������������������������       ������?0            @R@(       )                    �?    �b�?�             p@������������������������       ��)�� <�?2            @T@������������������������       ��6���N�?v            �e@+       .                    �?�ψ<���?J            @Z@,       -                    @��a_j�?             C@������������������������       �q=
ףp�?             4@������������������������       �����K�?             2@/       0                    @D`(\00�?/            �P@������������������������       �ƿ:Gf0�?             =@������������������������       �q9W��S�?             C@2       9                   �:@ݶE�]�?�           ؆@3       6                   �6@�����?%           @~@4       5                    �?������?I            �\@������������������������       ���(\���?             D@������������������������       ���$���?0            �R@7       8                   �9@�2sܘ�?�             w@������������������������       ���<<X�?�            �r@������������������������       �{	�%���?*             R@:       =                    �?y�l�x��?�            �n@;       <                   �=@������?!            �L@������������������������       ���&T���?             A@������������������������       �7����?             7@>       ?                    @0�z{�?y            �g@������������������������       ����k�?e            �c@������������������������       �     ��?             @@A       \                    �?	ʒ���?�           �@B       O                    @�J*���?�           (�@C       H                   �1@�v��'�?X           0�@D       G                    �?p|���z�?-            @S@E       F                    �?�GcT!)�?             3@������������������������       �Y�����?             &@������������������������       �      �?              @������������������������       �>�����?             M@I       L                    �?1ϵI3�?+           �{@J       K                   �=@�a�a�?p             e@������������������������       �?�%n(��?h             c@������������������������       �l�l��?             .@M       N                    �?�G���?�            q@������������������������       �&ޏ��k�??             V@������������������������       �ڕ7g��?|             g@P       U                    �?��;�'�?q            �g@Q       R                   �9@��g�?0            �S@������������������������       ��.k���?             �I@S       T                   �;@�M[\!	�?             ;@������������������������       ��
t�F��?
             1@������������������������       �R���Q�?             $@V       Y                    @\�x�?A            @\@W       X                    �?TQm�?)            �R@������������������������       �+7����?             7@������������������������       �,�wɃ�?             J@Z       [                   �3@���)�c�?             C@������������������������       ��ˠT�?             &@������������������������       �J�_cV�?             ;@]       l                   �2@PU �DF�?           p{@^       e                    @3��|-��?[            `a@_       b                    �?�	A���?,            �R@`       a                   �1@�-Z�?             =@������������������������       �$�ɜoB�?
             1@������������������������       ��q�q�?             (@c       d                    @!��wy��?             G@������������������������       �     ��?             @@������������������������       �������?
             ,@f       i                    @     L�?/             P@g       h                    @��]�`��?            �C@������������������������       �������?             .@������������������������       ��q�q�?             8@j       k                    @ �o_��?             9@������������������������       �      �?              @������������������������       �|�l�]�?             1@m       t                    @���R߽�?�            �r@n       q                   �5@fn̙R��?{            �g@o       p                    �?@�/,��?C            @X@������������������������       �<�i$���?            �E@������������������������       ����u���?(             K@r       s                    �?&b�Ѧ�?8            @W@������������������������       �Spo��?             =@������������������������       �     �?'             P@u       x                    @5��>���?F            �[@v       w                   �6@�	4-���?"            �J@������������������������       ��F_��C�?             =@������������������������       �9��8���?             8@y       z                   �:@�q�q�?$            �L@������������������������       �ڼ�8��?            �E@������������������������       ����S�r�?             ,@�t�bh�h4h7K ��h9��R�(KK{KK��h��BI       �{@      R@     v@      B@     �P@      7@     �U@     @�@     ��@     �P@     @S@     �e@     8�@     �y@      &@     @Q@     �I@     @b@     �N@      r@      E@      m@      7@     �B@      @      O@     �|@     �}@      H@     �G@     @]@     Pz@     0q@      @      H@      ?@      Z@      D@      f@      .@      W@      "@      @      �?      3@     w@     �t@      (@      3@     @P@     �l@      `@              (@      @     �D@      (@     �P@      @     �C@       @       @              @      K@      N@      @       @     �@@      N@      G@              @              2@      @      ?@      @      7@       @       @               @      2@      <@      �?      @      4@      D@      :@              �?              *@      @      4@              @                              �?      @      .@                       @      &@       @                              @              (@              @                                      @      @                              $@      @                                               @              @                              �?              &@                       @      �?      @                              @              &@      @      0@       @       @              �?      .@      *@      �?      @      (@      =@      2@              �?              "@      @       @      @      @               @                      *@      @              �?      @      0@      @              �?                              @      @      *@       @                      �?       @       @      �?      @      @      *@      ,@                              "@      @     �A@              0@                              �?      B@      @@       @      @      *@      4@      4@              @              @      @      ;@              .@                              �?      B@      :@               @      *@      4@      ,@              @              @      @      7@              ,@                              �?      8@      7@               @      (@      .@      *@              @               @      @      @              �?                                      (@      @                      �?      @      �?                              �?               @              �?                                              @       @       @                      @                               @              @              �?                                              @       @       @                                                                      �?                                                              �?                                      @                               @             �[@      "@     �J@      @      @      �?      0@     �s@     �p@      "@      &@      @@     `e@     �T@              @      @      7@      @     �F@      @      7@      �?                      @      i@      b@      @      @      .@      X@     �A@                              $@              :@       @      @                              @     �`@     �U@               @      @     �E@      .@                              �?               @                                                     �C@      7@               @              @                                                      2@       @      @                              @      X@      P@                      @      D@      .@                              �?              3@       @      4@      �?                      @     @P@     �L@      @      �?      "@     �J@      4@                              "@              *@      �?      2@      �?                      �?      B@      ?@       @              @      E@      ,@                               @              @      �?       @                               @      =@      :@      �?      �?       @      &@      @                              �?             �P@      @      >@      @      @      �?      $@     �\@      _@      @       @      1@     �R@     �G@              @      @      *@      @      F@      @      9@      �?      �?      �?      @     �W@     @Y@      @      @      (@     �P@      C@              @       @      @      @      6@      @      .@      �?      �?      �?      @      D@     �I@      @      @      @     �D@      <@               @      �?      �?      @      6@              $@                                     �K@      I@       @       @       @      :@      $@               @      �?      @      �?      6@      �?      @      @       @              @      4@      7@              �?      @       @      "@              @      @       @       @      "@      �?                                      @       @      $@                              @       @               @       @      @              *@              @      @       @                      (@      *@              �?      @      @      @              �?      �?      �?       @     @\@      ;@     �a@      ,@      @@      @     �E@     �V@     �b@      B@      <@      J@     �g@     `b@      @      B@      :@     �O@      <@     �F@      *@      J@      �?       @              "@     �H@     �X@      @      .@      (@     @S@     @Q@              @      @      5@      @      B@      &@      B@      �?       @              "@      ?@     �U@      @      ,@      "@     �J@     �N@              @      @      3@      @      1@      @      &@              �?                      2@      >@                      @      <@      4@                              �?      �?      @              @              �?                       @      3@                              .@      "@                                              (@      @       @                                      $@      &@                      @      *@      &@                              �?      �?      3@       @      9@      �?      �?              "@      *@      L@      @      ,@      @      9@     �D@              @      @      2@      @      $@      @      �?      �?      �?              @      @      :@       @      @      �?      @       @                      @      @       @      "@      @      8@                              @       @      >@       @      "@      @      4@     �@@              @       @      .@      @      "@       @      0@              @                      2@      (@      �?      �?      @      8@       @              @               @              @      �?      @                                      @      @                      �?      &@       @              @                              @      �?      @                                              �?                      �?      @                      @                               @                                                      @      @                              @       @                                               @      �?      *@              @                      .@      @      �?      �?       @      *@      @                               @               @               @              @                       @                              �?      "@      @                                                      �?      @               @                      *@      @      �?      �?      �?      @      @                               @              Q@      ,@      V@      *@      8@      @      A@     �D@     �J@      ?@      *@      D@     @\@     �S@      @      =@      4@      E@      5@     �G@      "@      M@      @      0@       @      2@     �B@     �A@      .@      $@      5@     �X@     �K@      @      *@      @      6@      &@      1@       @      ,@      @       @              @      "@      @      @      @      @      (@      2@              @      @       @              @              @                                      @      @                      @       @      &@              �?       @                      $@       @      &@      @       @              @       @      @      @      @      �?      $@      @              @      �?       @              >@      @      F@      @      ,@       @      .@      <@      =@      (@      @      0@     �U@     �B@      @       @      @      ,@      &@      ;@      @     �C@      @      $@       @      .@      3@      8@      (@      @      &@     �R@      :@       @      @      @      @      @      @              @              @                      "@      @                      @      (@      &@      �?       @      �?       @      @      5@      @      >@      @       @      @      0@      @      2@      0@      @      3@      .@      7@              0@      *@      4@      $@      @      �?       @      @      @      �?      "@      �?      @      @      @       @       @      @                              @              @      �?       @              @              "@      �?      @      @      �?      �?       @       @                                              @                      @              �?                              @       @      �?              @                              @              ,@      @      <@      @      @      @      @      @      *@      "@              1@      *@      0@              0@      *@      0@      $@      $@      @      7@       @      @      @       @      @      *@      "@              .@      (@      *@              0@      (@      @      "@      @              @      �?                      @                                       @      �?      @                      �?      "@      �?     �b@      >@     @^@      *@      =@      0@      8@     @W@     @^@      3@      >@     �L@     @h@     @a@       @      5@      4@      E@      5@      V@      3@     �T@      &@      5@      .@      &@      C@      O@      *@      6@     �E@     �Z@     @W@      @      ,@      2@      <@      3@      Q@      .@     �E@      @      .@      &@      @      @@     �K@       @      4@      :@      Q@      S@       @      *@      0@      6@      .@      7@       @      �?              @                      .@      @               @              (@      @              �?      @                      @                                                       @      �?                              @      �?                                              @                                                      @                                      �?                                                       @                                                       @      �?                               @      �?                                              1@       @      �?              @                      @      @               @              "@      @              �?      @                     �F@      *@      E@      @      $@      &@      @      1@      I@       @      2@      :@      L@     @Q@       @      (@      (@      6@      .@      :@      @      *@      @      @      @              @      3@      �?       @      "@      5@      5@              @      @      (@      @      5@      @      *@      @      @      @              @      3@      �?       @      "@      4@      5@              @      @      (@      @      @                                      �?                                      @              �?                      �?      �?                      3@       @      =@      @      @      @      @      *@      ?@      @      $@      1@     �A@      H@       @      @      @      $@      $@       @              .@      �?       @      �?      �?      "@      ,@                      @      *@      "@              @      @       @      @      1@       @      ,@       @      @      @      @      @      1@      @      $@      $@      6@     �C@       @       @       @       @      @      4@      @      D@      @      @      @      @      @      @      @       @      1@     �C@      1@       @      �?       @      @      @      @      �?      @              @      �?      @       @      @              �?       @      :@      @              �?      �?      @      @      @              @                      �?      @       @      @              �?       @      (@      @              �?              @      @      @      �?      @              @                              �?                              ,@                              �?              �?      �?      �?                                                      �?                              *@                                              �?       @              @              @                                                              �?                              �?                      ,@      @     �@@      @      @      @              @      @      @      �?      "@      *@      *@       @              �?       @               @      @      7@              @                      @      �?       @      �?      @      &@       @       @              �?       @              @               @                                                       @      �?       @       @      �?                      �?      �?              @      @      .@              @                      @      �?                      @      "@      @       @                      �?              @              $@      @              @              �?       @      @               @       @      @                                              @              �?                                                      @                      �?      @                                              @              "@      @              @              �?       @                       @      �?       @                                             �O@      &@      C@       @       @      �?      *@     �K@     �M@      @       @      ,@     �U@     �F@      @      @       @      ,@       @      9@      �?      .@               @                      ;@      6@      �?      @      �?      A@      @              �?                              (@              *@                                      "@      (@               @      �?      8@       @                                               @               @                                      @      @                              $@      �?                                                              �?                                      @      @                               @                                                       @              @                                                                               @      �?                                              $@              @                                      @       @               @      �?      ,@      �?                                              "@               @                                      @       @               @      �?      @                                                      �?              @                                      �?                                       @      �?                                              *@      �?       @               @                      2@      $@      �?      �?              $@      @              �?                              @      �?       @                                      *@      @                              @      @              �?                              @      �?                                               @      @                              @      �?                                              @               @                                      &@      @                                      @              �?                              @                               @                      @      @      �?      �?              @                                                                                                                      @      �?      �?               @                                                      @                               @                      @                                      @                                                      C@      $@      7@       @      @      �?      *@      <@     �B@      @      @      *@     �J@      C@      @      @       @      ,@       @      <@      @      0@       @      @              @      5@      8@       @      @      @      @@      6@      @      @      �?      "@       @      *@       @      &@       @      @               @       @      $@               @       @      :@      "@                      �?      @               @      �?              �?      @                      @      @                              ,@      @                              �?              @      �?      &@      �?                       @       @      @               @       @      (@      @                      �?      @              .@       @      @              �?               @      *@      ,@       @      @      @      @      *@      @      @              @       @      ,@       @      �?              �?                              �?                       @              @              �?               @              �?              @                               @      *@      *@       @      @      @      @       @      @      @              �?       @      $@      @      @               @      �?      "@      @      *@      @              @      5@      0@      �?       @      �?      @              @       @       @                               @       @      *@       @              @      "@      (@                      �?                      @              �?                               @       @      @                      @       @      &@                                                       @      �?                                               @       @               @      @      �?                      �?                      @      @      @               @      �?      @      @              �?              �?      (@      @      �?       @              @              @      �?       @               @              @      @              �?                      &@      @      �?       @               @                      @      @                      �?       @                                      �?      �?                                      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJJ9hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKehnh4h7K ��h9��R�(KKe��hu�B         0                    �?��6��?�	           ��@                            @N??���?b           ��@                          �1@hS�z�?!           �@                           @ֻ�����?�             j@                           �?^��p��?j            �c@                            �?��S����?             ;@������������������������       �r�q��?	             (@������������������������       �I�7�&��?             .@	       
                    @��&+*�?Y             `@������������������������       �e�X��?6            �R@������������������������       �V���s�?#             K@                           @;�;��?&             J@������������������������       ����,�?             3@                          �0@^p�F�?            �@@������������������������       ���!pc�?	             &@������������������������       ���ճC��?             6@                            �?�������?�           ܐ@                          �7@\����?�           ��@                          �4@�`'��4�?Z           `�@������������������������       �\��"e �?�             r@������������������������       �UiAG��?�            �p@                           �?���.�?�            �p@������������������������       ��E����?(             R@������������������������       �6�\&�C�?q            @h@                           @��Cq�?�            p@                           @W�v����?g            �d@������������������������       ��v`���?W            @a@������������������������       ��S�����?             =@                           @���5�?7            �V@������������������������       ������?(            @P@������������������������       �S�!�uq�?             9@        /                    @E�5ï��?A           p@!       (                    �?�B�V�c�?&           p|@"       %                    �?q�����?�            q@#       $                    @
Rt�?�?.            @S@������������������������       �t�@��?&             N@������������������������       �Iє�?             1@&       '                    �?����\��?|            �h@������������������������       �=����?'            �K@������������������������       ��ȼ��?U            �a@)       ,                    @�w�[�?|            �f@*       +                   �:@     F�?W             `@������������������������       ��p%]^z�?Q             ]@������������������������       ��q�q�?             (@-       .                    @��3L���?%             K@������������������������       ���8��8�?	             (@������������������������       ��!͎�?             E@������������������������       �9��8���?             H@1       P                     @E;s�I��?=           ��@2       A                    �?")x���?�           ,�@3       :                   �2@1�8�#D�?y           H�@4       7                    �?�}����?G            �[@5       6                    �?����X�?            �A@������������������������       �x�"w���?             3@������������������������       �     ��?             0@8       9                    �?u#����?/             S@������������������������       ���k���?             6@������������������������       ���rᮾ�?              K@;       >                    �?�Nt�$t�?2           �}@<       =                    �?R�3�Y�?U            �a@������������������������       �������?!             L@������������������������       �XٙZ�?4            @U@?       @                   �<@w�s@���?�            �t@������������������������       ��R�c@�?�            �p@������������������������       �g���6W�?+            �P@B       I                   �5@��<1	9�?)           �@C       F                   �1@���2&�?>           Ѐ@D       E                     �?�u,*/�?^            `d@������������������������       ��Q�S�?D            @^@������������������������       ��2q�{�?             E@G       H                     �?�5��?�            pw@������������������������       ��f�	�?�            �p@������������������������       ��r��� �?A            �Z@J       M                   �6@\��"e��?�            �v@K       L                    @E�
��3�?3            @Q@������������������������       �x^�V��?%            �H@������������������������       ��(\����?             4@N       O                     �?������?�            0r@������������������������       �9��8���?x             h@������������������������       �a�����?@            �X@Q       ^                    @ףp=
�?�            �@R       Y                    @�89~��?~           ��@S       V                    �?D,���?�            w@T       U                   �5@l~X�<�?,             R@������������������������       ��)O�?             B@������������������������       �������?             B@W       X                   �9@�nF���?�            �r@������������������������       ��M��S��?�            �n@������������������������       ����{qg�?#            �I@Z       [                   �0@�i#���?�            �k@������������������������       �      �?              @\       ]                   �?@#�a���?�            �j@������������������������       �
7�Ȋ�?�            `i@������������������������       ��8��8��?             (@_       `                   �3@9��8�c�?             H@������������������������       �X�<ݚ�?             "@a       b                    �?>]6�I��?            �C@������������������������       ��q-�?             *@c       d                    @f�.y0��?             :@������������������������       �:߄*�u�?             1@������������������������       �B{	�%��?             "@�t�bh�h4h7K ��h9��R�(KKeKK��h��B�;       P}@     @U@     �s@      D@     �S@      5@     �T@     ��@     Ђ@      M@     �R@      b@      �@     �{@      ,@      O@      K@     �_@      N@      k@      >@     �`@      @      0@      @     �@@     �u@      s@      (@      ?@      J@     �r@     @g@      �?      8@      ;@     �G@      5@     `d@      3@     �U@      @       @              1@     pq@      o@      $@      6@     �@@     `i@     @_@              .@      &@     �@@      (@      1@      �?      @                               @     �Y@      J@              �?       @      6@      @                              �?              *@      �?      @                               @      U@      B@              �?       @      (@       @                                              @              @                                      "@      @                       @      �?      �?                                               @              @                                       @      @                              �?      �?                                               @                                                      @      @                       @                                                              "@      �?                                       @     �R@      =@              �?              &@      �?                                              @      �?                                       @      H@      &@              �?               @                                                      @                                                      ;@      2@                              @      �?                                              @              �?                                      2@      0@                              $@       @                              �?              @              �?                                      @      @                              @                                      �?              �?                                                      *@      &@                              @       @                                                                                                      @      @                               @                                                      �?                                                      "@      @                              @       @                                             @b@      2@     �T@      @       @              .@      f@     �h@      $@      5@      ?@     �f@     @^@              .@      &@      @@      (@      `@      .@      N@      @      @              ,@     �[@     ``@       @      4@      8@      b@     �W@              (@      $@      =@      (@     @W@      @     �B@       @      @              @     @V@      X@      @      "@      (@     �^@      O@              @       @       @              H@      @      $@       @                      �?     �O@      F@      @      @       @      K@     �A@              @              @             �F@      �?      ;@              @              @      :@      J@       @      @      @      Q@      ;@                       @      @              B@       @      7@      �?       @              "@      6@     �A@       @      &@      (@      7@      @@              "@       @      5@      (@      0@      @      @              �?              @      @      0@       @      @      �?      @      @                      �?      @              4@      @      3@      �?      �?              @      1@      3@              @      &@      2@      ;@              "@      @      0@      (@      1@      @      6@              @              �?     �P@     @P@       @      �?      @      B@      ;@              @      �?      @              *@      �?      1@               @              �?     �H@      ;@       @      �?      @      9@      3@              @      �?      �?              *@      �?      1@               @              �?      :@      8@       @      �?      @      8@      1@              @      �?      �?                                                                      7@      @                              �?       @                                              @       @      @              �?                      1@      C@                       @      &@       @                               @              @       @      @                                      (@     �A@                              @      @                                              �?               @              �?                      @      @                       @      @      @                               @             �J@      &@      G@      @       @      @      0@     �Q@      L@       @      "@      3@      X@     �N@      �?      "@      0@      ,@      "@     �J@      &@      D@      @      @      @      "@     @Q@      J@      �?      "@      0@     �T@      N@      �?       @      *@      &@      @      @@      @      9@      @      @       @      "@      <@      >@              @      (@     �C@      E@      �?      @      *@       @      @      @      @       @                      �?              (@      "@              @      @       @      .@              @              �?              @      @       @                      �?              (@      @              @      �?      @      $@              @              �?               @                                                               @                      @      @      @                                              :@      @      1@      @      @      �?      "@      0@      5@              @      @      ?@      ;@      �?      �?      *@      @      @      .@      �?      @              �?                       @      @              �?              @      .@                              @      �?      &@       @      ,@      @      @      �?      "@      ,@      0@               @      @      8@      (@      �?      �?      *@      @      @      5@      @      .@              �?      �?             �D@      6@      �?      @      @      F@      2@               @              @      �?      1@      @      &@              �?      �?              ;@      1@              �?       @      C@      @              �?              �?      �?      1@      @      &@              �?      �?              ;@      .@                       @      >@      @                              �?      �?                                                                       @              �?               @                      �?                              @              @                                      ,@      @      �?       @       @      @      *@              �?               @               @                                                      �?      �?                                      @              �?              �?               @              @                                      *@      @      �?       @       @      @      @                              �?                              @              �?              @       @      @      �?              @      *@      �?              �?      @      @      @     �o@     �K@     �f@      A@      O@      2@     �H@      l@     �r@      G@     �E@     @W@     �s@     �o@      *@      C@      ;@     �S@     �C@     `g@      @@     �\@      2@      E@      @      C@      g@     `l@      A@      ;@     �M@     �k@     �c@      @      9@      4@      L@      ?@     �O@      .@      M@      @      8@      @      0@      D@      Q@      ,@      .@      ?@     �T@     �Q@      �?      1@      .@      :@      3@      0@              @                              �?      ,@      <@       @      �?       @      :@      @                              @      �?      &@                                              �?      @      @              �?      @      @      @                              �?               @                                                       @      @                       @      �?       @                                              @                                              �?      @      @              �?      �?       @      �?                              �?              @              @                                      "@      5@       @              @      7@       @                               @      �?       @              �?                                       @      "@      �?               @      @                                                      @              @                                      @      (@      �?              @      2@       @                               @      �?     �G@      .@      J@      @      8@      @      .@      :@      D@      (@      ,@      7@      L@     @P@      �?      1@      .@      7@      2@      ;@      �?      ,@              @              @      &@      2@       @       @      @      2@      5@      �?              @      @       @      $@                               @              @      @      (@               @       @      @      $@                      �?      �?       @      1@      �?      ,@               @              @      @      @       @               @      (@      &@      �?              @      @              4@      ,@      C@      @      4@      @      "@      .@      6@      $@      (@      3@      C@      F@              1@      &@      1@      0@      4@      $@      @@      @      .@       @      @      .@      1@       @      "@      (@      C@      D@              &@      �?      (@      ,@              @      @       @      @       @      @              @       @      @      @              @              @      $@      @       @      _@      1@      L@      &@      2@      @      6@      b@     �c@      4@      (@      <@     @a@     @V@       @       @      @      >@      (@     �S@      @      6@      �?       @              $@      _@     �\@       @      @      1@     �R@     �I@              @       @      @      "@      5@       @      @                              �?     �F@     �I@              �?      @      4@      (@                                      �?      .@       @      �?                                      ?@     �F@              �?       @      .@       @                                      �?      @              @                              �?      ,@      @                       @      @      @                                              M@      @      1@      �?       @              "@     �S@     �O@       @      @      *@      K@     �C@              @       @      @       @      E@      �?      &@      �?      @              "@      J@     �D@       @      @      *@      >@     �B@              @       @      @      @      0@      @      @               @                      ;@      6@                              8@       @                               @       @     �F@      &@      A@      $@      $@      @      (@      4@     �F@      2@      @      &@      P@      C@       @      @      @      7@      @      (@      �?      $@      @      �?                       @      @               @      @      @      (@              �?              @              $@      �?      @                                       @      @               @      @      @       @              �?              @               @              @      @      �?                              �?                      �?              @                                             �@@      $@      8@      @      "@      @      (@      (@      C@      2@      @      @     �N@      :@       @       @      @      3@      @      7@      @      3@       @      @              @      @      <@      "@      @      @      I@      0@               @      �?      (@      �?      $@      @      @      @      @      @      @      @      $@      "@              �?      &@      $@       @               @      @       @     �P@      7@     @Q@      0@      4@      &@      &@     �D@     �Q@      (@      0@      A@     @W@      X@      $@      *@      @      7@       @     �K@      6@     �L@      .@      4@      $@       @     �B@     @Q@      (@      ,@      >@     �V@     �W@      "@      *@      @      6@       @      C@      (@      ?@      &@      ,@       @      @      5@     �I@      $@      $@      2@     �L@      J@      �?       @      @      ,@      @      @       @       @              �?                      @      @      @      @      �?      4@      .@               @       @      @               @               @                                       @       @              @      �?      1@      @                      �?                       @       @                      �?                      @      @      @                      @      "@               @      �?      @              A@      $@      =@      &@      *@       @      @      .@     �F@      @      @      1@     �B@     �B@      �?      @      @      $@      @      @@      $@      :@      @       @      �?      �?      .@     �D@       @      @      0@      B@      ?@              @      @      @               @              @      @      @      @      @              @      @              �?      �?      @      �?      @      �?      @      @      1@      $@      :@      @      @       @      @      0@      2@       @      @      (@     �@@      E@       @      @      �?       @      @                                      �?                      @                                              �?                                              1@      $@      :@      @      @       @      @      $@      2@       @      @      (@     �@@     �D@       @      @      �?       @      @      .@      $@      9@      @      @       @      @      $@      2@       @      @      &@     �@@     �D@      @      @      �?       @      �?       @              �?                                                                      �?                      @                              @      &@      �?      (@      �?              �?      @      @       @               @      @      @       @      �?                      �?              @               @                                                                                                                      �?              @      �?      $@      �?              �?      @      @       @               @      @      @       @      �?                                       @              @                                      @                                              �?                                              @      �?      @      �?              �?      @      �?       @               @      @      @      �?      �?                                      @      �?       @      �?              �?                       @               @      @              �?                                                              �?                              @      �?                                      @              �?                                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�@vhhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKmhnh4h7K ��h9��R�(KKm��hu�B�         6                   �2@�<P���?�	           ��@                           �??`�� l�?�           ��@                            @t8vȿ��?\           ��@                           @z�s���?           y@                           @Dp�N���?_            `c@                            �?     ,�?N             `@������������������������       ����/]��?G            @\@������������������������       ��h$���?             .@	       
                     �?B{	�%��?             ;@������������������������       �"pc�
�?             &@������������������������       �     @�?             0@                           @$�����?�            �n@                          �1@�'ୡs�?�            `g@������������������������       ��o	��?U             ]@������������������������       ��	Mo�?.            �Q@                          �0@�����?%            �M@������������������������       �hE#߼�?             .@������������������������       ��!pc��?             F@                          �0@�4 ��;�?U            �`@                           @      �?             @@������������������������       �Iє�?	             1@������������������������       ��'}�'}�?             .@                           @��ͪ���?D             Y@                           @�1�L�?8            �T@������������������������       �_��"�O�?.             Q@������������������������       �{�G�z�?
             .@������������������������       �	6c����?             1@       +                    @� �e���?N           p�@       $                   �0@~t�M�?�            �w@       !                    @I��PK��?-            @P@                             @��-]W��?            �E@������������������������       ��I+��?             9@������������������������       ��^B{	��?             2@"       #                    @
�GN��?             6@������������������������       ��'}�'}�?             .@������������������������       �4և����?             @%       (                    @�f'���?�            �s@&       '                    @3hI�g�?�            �k@������������������������       �:l�A�?_            �b@������������������������       �0�����?/             R@)       *                   �1@n?���?5            @W@������������������������       ��(\����?             I@������������������������       ��|S�ݮ�?            �E@,       1                    @k5(ˋ�?^            @b@-       .                   �0@���(�?G            �\@������������������������       ��.�?��?             .@/       0                    �?l	��g��?<             Y@������������������������       ����y4F�?             3@������������������������       ����'F��?1            @T@2       3                    �?������?             ?@������������������������       �      �?              @4       5                     �?K����?             7@������������������������       ��G�z��?             $@������������������������       �
ц�s�?	             *@7       N                    �?R:�@��?           L�@8       G                   �?@d�=BP�?5           ��@9       @                    �?Tho�+�?           ��@:       =                   �;@&�����?�            �v@;       <                    �?����p��?�            �s@������������������������       ��Oqx��?J            @_@������������������������       �J�AI��?y            �g@>       ?                     �?���y� �?            �H@������������������������       �B{	�%��?             "@������������������������       �      �?             D@A       D                   �6@G���15�?$           ��@B       C                   �3@j �`��?�            �x@������������������������       ���,��.�?5            �T@������������������������       �3����l�?�            `s@E       F                    @!N���n�?4           �~@������������������������       �9G%�i�?-           P~@������������������������       ��n���?             "@H       I                    �?x�5?,�?1             R@������������������������       �      �?             (@J       M                   �@@ϊF�y�?*             N@K       L                    �?�L-���?             ;@������������������������       �ffffff�?             $@������������������������       ��������?             1@������������������������       ��wC�Ҁ�?            �@@O       ^                     @ ���Fd�?�           �@P       W                   �:@�A�Q�7�?
           �@Q       T                   �5@�`A:���?�           L�@R       S                    @�h`A�?h           ��@������������������������       �4�\�K2�?N           ��@������������������������       �-�R��?            �B@U       V                    �?!���T�?.           �}@������������������������       ���Y� ��?g            �c@������������������������       �     T�?�             t@X       [                   �=@юc:W�?t            �e@Y       Z                    �?�j��t�?E            �[@������������������������       ���g�g�?             �M@������������������������       ��$B`~�?%            �I@\       ]                    �?q�{%�?/            @P@������������������������       ���&��?             9@������������������������       ��������?             D@_       f                    �?�*+�D��?�            �s@`       c                   �9@���;vR�?[            �a@a       b                    @�0�" ��?J            �\@������������������������       ���ђ�?,            �N@������������������������       ���?Z�9�?             K@d       e                    @6|���t�?             :@������������������������       ��T�6|��?             *@������������������������       ��T�6|��?	             *@g       j                   �7@��e Ʊ�?k            �e@h       i                    @θ	j*�?@             Z@������������������������       ���;�V��?            �@@������������������������       ��Y:s��?,            �Q@k       l                   �>@pB躍�?+             Q@������������������������       �Э�*��?$             M@������������������������       �>
ףp=�?             $@�t�bh�h4h7K ��h9��R�(KKmKK��h��B�@        |@     �Q@     �u@     �A@     �R@     �A@     �Q@     `�@     ��@     �O@      U@     �c@     �@      {@      &@      P@      J@     @`@      O@     �`@       @     �J@      �?      @              $@     ps@      i@       @      @      5@      e@     �V@              $@       @      ?@      @     @R@              4@                              @      i@     �Y@      @      �?      $@     @S@     �B@              @              @             �H@              (@                               @     @d@      V@      �?      �?      "@      I@      ;@                                              8@              @                                     �H@      A@              �?      @      6@      &@                                              .@              @                                      G@      9@                      @      2@      &@                                              ,@              @                                     �E@      6@                      @      (@      &@                                              �?               @                                      @      @                              @                                                      "@                                                      @      "@              �?      �?      @                                                                                                               @      @                              @                                                      "@                                                      �?      @              �?      �?      �?                                                      9@              @                               @     @\@      K@      �?               @      <@      0@                                              .@              @                               @     �W@      E@                              4@      $@                                              (@              @                               @     �O@      9@                              "@       @                                              @                                                      @@      1@                              &@       @                                              $@               @                                      2@      (@      �?               @       @      @                                              @                                                      &@      �?                                                                                      @               @                                      @      &@      �?               @       @      @                                              8@               @                              �?      C@      ,@       @              �?      ;@      $@              @              @              @                                                      ,@      @                              @      @                                              @                                                      @      �?                              @      @                                              @                                                      "@       @                              �?                                                      1@               @                              �?      8@      &@       @              �?      6@      @              @              @              1@              @                              �?      7@      @      �?              �?      1@      @              @              @              .@               @                              �?      .@      @      �?              �?      1@      @              @              @               @              @                                       @       @                                                                                                      @                                      �?      @      �?                      @                                      �?             �M@       @     �@@      �?      @              @     �[@     �X@      @      @      &@     �V@     �J@              @       @      ;@      @     �H@       @      8@      �?      @              @      U@      O@      @      @       @     �S@      >@              @       @      "@       @      (@               @                                      8@      &@                              $@      @                              �?              "@                                                      *@      @                              $@      @                                              �?                                                      $@       @                               @      @                                               @                                                      @      @                               @                                                      @               @                                      &@      @                                      �?                              �?               @                                                      "@      @                                      �?                                              �?               @                                       @      �?                                                                      �?             �B@       @      6@      �?      @              @      N@     �I@      @      @       @      Q@      9@              @       @       @       @      @@       @      2@      �?      @              @     �B@      =@      @      @      @      L@      .@               @       @      @              8@       @      "@      �?      @              @      4@      6@      �?      @      @      ?@      *@               @       @      @               @              "@                                      1@      @      @      �?              9@       @                                              @      @      @                              @      7@      6@                      �?      (@      $@               @               @       @      @      @                                              @      3@                      �?      $@      @              �?               @              �?      @      @                              @      0@      @                               @      @              �?                       @      $@              "@                                      ;@     �B@      �?              @      *@      7@              @              2@       @       @              @                                      9@     �@@                       @      &@      .@              @              1@                                                                      @      "@                              �?                                                       @              @                                      4@      8@                       @      $@      .@              @              1@                               @                                              @                                       @                               @               @              @                                      4@      1@                       @      $@      *@              @              "@               @               @                                       @      @      �?              �?       @       @                              �?       @      @                                                                      �?              �?                                                               @               @                                       @      @                               @       @                              �?       @                                                               @      @                                      �?                              �?       @       @               @                                                                               @      @                                             �s@     �O@     pr@      A@     �Q@     �A@     �N@     Pq@     `y@     �K@     �S@     @a@     �y@     `u@      &@      K@      I@     �X@      M@     �b@      @@      c@      .@     �I@      @@      >@      R@     �`@      9@     �E@     @T@     �e@      d@       @      >@      C@      H@      G@     `b@      @@     �b@      $@      D@      ;@      =@      R@     �`@      7@      C@     �Q@     �e@     �c@      @      ;@      >@      G@      F@     �N@      @      >@              (@      @      @      6@     �F@      @      .@      0@     �I@      G@      @       @      $@      *@      (@     �G@      @      =@              "@      @       @      6@     �C@      @      $@      0@     �H@     �B@      @      @      $@      *@       @      0@       @      @               @              �?      $@      3@      @      @      "@      6@      (@              @      @      �?      @      ?@       @      7@              @      @      �?      (@      4@      �?      @      @      ;@      9@      @       @      @      (@      @      ,@              �?              @      �?       @              @      �?      @               @      "@              �?                      @      @                                                              �?                                      �?                                              @              �?              @      �?       @              @      �?      @               @       @              �?                      @     �U@      <@     �]@      $@      <@      4@      9@      I@     �U@      1@      7@     �K@      _@     �[@              3@      4@     �@@      @@     �L@      "@      J@      @      @      @      @      9@      @@       @      $@      8@     @R@     �G@              @       @      4@       @      *@              @      �?                              "@      (@      �?              @      &@      *@                      �?      @      @      F@      "@     �G@      @      @      @      @      0@      4@      @      $@      4@      O@      A@              @      �?      *@      @      =@      3@     �P@      @      6@      *@      6@      9@     �K@      "@      *@      ?@     �I@      P@              .@      2@      *@      8@      9@      3@     �P@      @      6@      *@      6@      9@     �K@      "@      &@      ?@      H@      P@              .@      2@      *@      8@      @                                                                               @              @                                                      @              @      @      &@      @      �?              �?       @      @      $@              @      @      @       @       @       @                                      @                                              �?      @                              �?                              @              @      @      @      @      �?              �?       @      @      @              @      @       @       @       @       @      @              �?      @      �?      @                              �?      @                      @               @      @                      @                                                                               @                      �?                      @                                      �?      @      �?      @                              �?      �?                       @               @      �?                      �?              @       @      @              �?              �?      �?      �?      @                      @              @       @       @     �d@      ?@     �a@      3@      4@      @      ?@     �i@     q@      >@     �A@     �L@     �m@     �f@      @      8@      (@     �I@      (@     �`@      7@     �^@      (@      1@      @      4@     �d@     `m@      9@      =@     �E@     �g@     �`@       @      1@      "@      @@      @     �^@      .@     @X@      "@      &@              .@      c@     �k@      *@      :@     �@@     `e@      [@      �?      *@      @      9@      @     �Q@      @      I@       @      @               @     �Y@      a@      @      (@      1@     @V@      I@              @      @      &@      @      P@      @     �F@       @      @              �?     �Y@     �_@      �?      &@      1@      T@      I@              @      @      &@      @      @              @                              �?              $@      @      �?              "@                                                      J@      &@     �G@      @      @              *@     �I@     @U@      @      ,@      0@     �T@      M@      �?       @       @      ,@      �?      0@      @      (@              �?              @      4@     �C@      @      �?      @      1@      6@              @              �?              B@      @     �A@      @      @               @      ?@      G@       @      *@      $@     @P@      B@      �?      @       @      *@      �?      (@       @      9@      @      @      @      @      (@      *@      (@      @      $@      4@      8@      �?      @      @      @      @      $@      @      0@      �?      @      �?      @      &@      $@       @      @      @      $@      "@      �?       @       @      @      @      @      @      @              @              @      &@      "@      �?      �?      @      "@      @                               @              @      @      &@      �?              �?       @              �?      @       @      �?      �?      @      �?       @       @      �?      @       @       @      "@       @      �?       @              �?      @      @              @      $@      .@               @       @      @               @               @                                      �?              �?                      @      $@               @                                       @      @       @      �?       @                      @      @              @      @      @                       @      @              ?@       @      4@      @      @              &@      D@      C@      @      @      ,@     �F@      I@      �?      @      @      3@      @      &@       @      @      �?      �?                      <@      2@      @      @       @      3@      4@              @      �?      "@              "@      �?      @      �?      �?                      <@      (@      @      @      @      ,@      3@              @      �?       @              @      �?      �?      �?      �?                      2@       @               @       @      "@      $@                      �?                       @              @                                      $@      @      @       @      @      @      "@              @               @               @      �?       @                                              @               @       @      @      �?              @              �?              �?              �?                                              @               @       @      �?      �?                                              �?      �?      �?                                              �?                              @                      @              �?              4@      @      *@      @       @              &@      (@      4@       @              @      :@      >@      �?               @      $@      @      *@      @      &@      @      �?              @      @      (@                      @      6@      .@                               @      @              �?       @              �?              �?      �?      @                              @      @                              @              *@       @      @      @                       @      @       @                      @      .@      &@                               @      @      @      @       @      @      �?               @      @       @       @               @      @      .@      �?               @       @       @      @       @      �?      @      �?               @      @      @                       @      @      ,@                       @       @       @              �?      �?                                      @      �?       @                              �?      �?                                �t�bub�2'     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJTX�nhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKyhnh4h7K ��h9��R�(KKy��hu�Bx         >                    @�
����?�	           ��@       !                   �4@p'�O��?`           n�@                           �?Ȣ�}|��?           h�@                          �1@�'�����?�            �s@                          �0@�@B���?H            �^@                           �?��>4և�?             E@������������������������       �-)���?             =@������������������������       �����W�?             *@	       
                    �?��(\���?0             T@������������������������       ��]1�[��?            �@@������������������������       �L�i��J�?            �G@                           �?m |�F��?�            �h@                           �?jq�QP��?y             e@������������������������       �6��Lz)�?T            �]@������������������������       �8�e�?%            �I@                           �?��F�� �?             ;@������������������������       ���8��8�?             (@������������������������       ��|�j��?	             .@                            �?p�?��?M           x�@                           @���g6i�?g            �d@                           �?Ztjط}�?.            @R@������������������������       ����C���?             ?@������������������������       �h5����?             E@                          �0@����%�?9            �W@������������������������       �B{	�%��?             "@������������������������       �x�)�J�?2            @U@                           @�!�{6�?�            �x@                            �?�����?�            �m@������������������������       �     ��?(             P@������������������������       ���0å�?h            �e@                            �?:ٱ���?V            @c@������������������������       ��'���s�?$            �N@������������������������       ��H6&��?2            @W@"       1                     @�<���J�?A           (�@#       *                   �<@�sW�1�?           H�@$       '                   �7@1�嶏��?�           ��@%       &                    �?�fP�[�?�            Pu@������������������������       �&��AX��?Y            �a@������������������������       �HP�s�?w             i@(       )                    �?��H���?�            �u@������������������������       �DaH�,�?Y            �_@������������������������       �5�(����?�            �k@+       .                   @A@��z�ք�?T             c@,       -                   �=@� 2�xj�?G            �`@������������������������       �������?            �C@������������������������       �
�	�)D�?3            �W@/       0                    @P7�Z�?             3@������������������������       ��(\����?             $@������������������������       ���"e���?             "@2       9                    �?�y��b�?9           �@3       6                    �?��B���?�             k@4       5                    @Ec�[���?            �E@������������������������       �     ��?             @@������������������������       ��zv��?             &@7       8                    �?��@b���?m            �e@������������������������       ��"���?V            �a@������������������������       ��K>7�5�?            �@@:       =                   �@@AD˩�m�?�            �r@;       <                   �5@�� P�?�            �q@������������������������       �F_x����?            �I@������������������������       ��A����?�             m@������������������������       ��θ�?             *@?       ^                     @�
��?1           H�@@       O                    �?,��Ŝ�?n           ��@A       H                    �?���#Ae�?�           �@B       E                   �4@�K�=[��?�            �p@C       D                    @|�0�W��?d            �e@������������������������       ���)�8�?(             Q@������������������������       ��u��'�?<            @Z@F       G                     �?H�~Z���?A             W@������������������������       ��\@˜��?             7@������������������������       �j'����?0            @Q@I       L                   �7@�Qw
A�?           �{@J       K                    @���{B�?�            Pu@������������������������       �Sez�h�?_            �c@������������������������       �����P�?r             g@M       N                    @�[ A��?D             Y@������������������������       �������?
             .@������������������������       ��_8���?:            @U@P       W                    @J�uU�~�?�           ��@Q       T                    �?ܼ���?�            �s@R       S                   �8@*0F%��?�            �j@������������������������       ��z����?t            `f@������������������������       �|L�Sw�?            �A@U       V                   �5@t��f|�?A            @Y@������������������������       ��h�*$��?&            �L@������������������������       ������?             F@X       [                   �6@�����s�?�            0v@Y       Z                    @v�P1�?�             m@������������������������       ��6v�Y��?i            �c@������������������������       ��&'h�?-            @R@\       ]                    @�	Q�?Q            �^@������������������������       ���OF6��?4            @T@������������������������       ��q�q�?             E@_       j                    @����ҕ�?�             s@`       c                    �?��^�u�?2            @T@a       b                    @"�O�|�?             A@������������������������       ����I��?             1@������������������������       ��P�n#�?             1@d       g                   �3@]�޾��?            �G@e       f                   �1@��JÝ�?             7@������������������������       �     ��?	             0@������������������������       �������?             @h       i                    @�q�q�?             8@������������������������       �     @�?             0@������������������������       �      �?              @k       r                   �2@n����?�             l@l       o                   �1@�m���?2            �R@m       n                   �0@     ��?             @@������������������������       �6�h$��?
             .@������������������������       �v�f��?             1@p       q                    �?nR�-��?             E@������������������������       �O��E��?             2@������������������������       ��������?             8@s       v                    @ٽÆM��?_            �b@t       u                   �4@N�7��?             =@������������������������       �U��6���?	             1@������������������������       ���8��8�?             (@w       x                    @(CiVX�?N            �^@������������������������       ���!ZA�?F            @[@������������������������       �ݾ�z�<�?             *@�t�bh�h4h7K ��h9��R�(KKyKK��h��B�G       p}@     �S@     �t@      ;@     �O@      :@     @V@     h�@     �@     �Q@      X@     �g@     �@     P}@      1@     �R@      D@     @a@      K@     �q@      H@     �k@      1@     �K@      9@      J@     �h@     0p@      K@     �P@      ]@     �s@      r@      (@     �G@      <@     �W@      F@     �_@      "@     �P@      �?      *@              &@     �b@     `b@      &@      $@      @@     �b@     @X@               @      �?     �A@      ,@     �F@      @      ,@              $@              @     @R@     �N@      �?      @      (@      B@     �@@              �?              (@      @      6@               @              @              @     �D@      .@      �?      �?      @      2@      @                                      @      ,@              �?                                      1@      @                              @       @                                              "@              �?                                      *@      �?                              @       @                                              @                                                      @      @                              �?                                                       @              �?              @              @      8@      &@      �?      �?      @      ,@      @                                      @      @              �?                                      ,@      @      �?               @      @      �?                                               @                              @              @      $@      @              �?      @      &@       @                                      @      7@      @      (@              @              �?      @@      G@              @      @      2@      <@              �?              (@              5@      @      "@              @              �?      9@      D@              @      @      1@      ;@              �?              &@              ,@      @       @              @              �?      2@      7@              @      @      (@      .@                              &@              @              �?                                      @      1@                      �?      @      (@              �?                               @       @      @               @                      @      @              �?      �?      �?      �?                              �?                              �?                                       @      @                              �?      �?                              �?               @       @       @               @                      @                      �?      �?                                                             @T@      @      J@      �?      @              @     �R@     �U@      $@      @      4@      \@      P@              @      �?      7@      &@      :@              "@      �?                              >@      =@              �?      @     �G@      "@                              @      @      "@               @      �?                              (@      "@                       @     �@@      @                                       @      @                                                       @       @                       @      (@                                               @      @               @      �?                              $@      �?                              5@      @                                              1@              @                                      2@      4@              �?      @      ,@      @                              @       @                                                              �?      @                                      �?                                              1@              @                                      1@      *@              �?      @      ,@      @                              @       @     �K@      @     �E@              @              @     �F@     �L@      $@      @      *@     @P@     �K@              @      �?      3@      @      A@      @      =@                              @      C@      8@      @      @      @     �E@      C@              @      �?      @      @      *@               @                               @      *@      @              �?       @      @      .@              @      �?              �?      5@      @      ;@                              @      9@      3@      @       @       @     �B@      7@              @              @       @      5@              ,@              @                      @     �@@      @      �?      "@      6@      1@              �?              .@      @      (@              @               @                      �?      2@      @              @      "@                      �?              @              "@              $@              �?                      @      .@      @      �?       @      *@      1@                              (@      @      d@     �C@     �c@      0@      E@      9@     �D@     �I@      \@     �E@     �L@      U@     �d@      h@      (@     �C@      ;@      N@      >@     �\@      :@     �\@      @      7@       @      :@      A@     �R@      ;@      A@      F@      \@     �Y@              4@      *@      J@      ,@     @W@      7@     �X@      �?      ,@      @      2@      A@     @P@      2@      :@      >@     �Y@     �W@              *@      @      A@      &@      O@      @      K@              @      �?      "@      6@     �C@       @      .@      .@      F@      D@              @       @      1@      @      7@      @      @@              @              @      *@      2@               @      $@      3@      (@                               @             �C@      @      6@               @      �?      @      "@      5@       @      *@      @      9@      <@              @       @      .@      @      ?@      0@     �F@      �?       @      @      "@      (@      :@      0@      &@      .@     �M@     �K@              $@      @      1@       @      (@      @      0@      �?                      @      @      *@              @      @      3@      <@              @      @      @      �?      3@      "@      =@               @      @      @      "@      *@      0@      @      (@      D@      ;@              @       @      $@      @      5@      @      .@      @      "@      @       @              "@      "@       @      ,@      "@      @              @      @      2@      @      5@      @      "@      @      "@      @       @              @      @       @      "@      "@      @              @      @      2@       @      "@              @              @               @               @                      @      �?       @               @               @       @      (@      @      @      @       @      @      @              @      @       @      @       @      @              @      @      0@                              @                                               @       @              @              �?               @                      �?                      @                                                       @               @              �?               @                                              @                                               @                      @                                                      �?     �G@      *@      E@      (@      3@      1@      .@      1@      C@      0@      7@      D@      K@     �V@      (@      3@      ,@       @      0@      8@      @      .@      @      @      @       @      "@      3@       @       @      ,@      B@      B@      @      @      "@      @      @                      @                      �?      @      @       @       @       @      @      $@      �?               @              �?       @                      @                      �?              �?       @       @       @      �?       @                       @              �?       @                                                      @       @                              @       @      �?                                              8@      @      &@      @      @      @      @      @      &@              @      $@      :@     �A@      @      @      "@      @      @      7@       @      @       @      @      @      @      @       @              @       @      1@      =@      @      @      "@      @      @      �?      �?      @      �?                              @      @               @       @      "@      @              �?                              7@      $@      ;@      "@      ,@      &@      @       @      3@      ,@      .@      :@      2@     �K@      "@      (@      @      @      $@      7@      $@      :@      "@      ,@      &@      @       @      3@      ,@      *@      8@      2@     �K@      @      (@      @      @       @      @      @      "@              @       @      @              �?      @              @      @       @                      @      �?              1@      @      1@      "@      "@      "@       @       @      2@      $@      *@      5@      (@     �J@      @      (@      �?      @       @                      �?                                                               @       @                      @                               @      g@      >@     �[@      $@       @      �?     �B@     `t@     �s@      0@      =@      R@     pp@     `f@      @      <@      (@     �E@      $@     �b@      4@     @V@      $@      @      �?      9@     �q@     �q@      ,@      5@      L@     �j@     �a@      @      2@      &@      @@      @      O@      @     �C@              @              $@      g@     �d@      @       @      4@     �^@     �P@               @      @       @      �?      1@       @      $@                               @     �U@     �S@      �?      @      "@     �C@      2@                                              @      �?      @                                     �S@     �D@                       @      6@      "@                                               @      �?                                              2@      7@                      @      .@      @                                              @              @                                      N@      2@                      @      @      @                                              $@      �?      @                               @       @     �B@      �?      @      �?      1@      "@                                              @                                              �?      �?      &@      �?      �?               @       @                                              @      �?      @                              �?      @      :@               @      �?      .@      @                                             �F@      @      =@              @               @     �X@     @V@      @      @      &@      U@      H@               @      @       @      �?     �A@       @      0@               @              @     @V@      T@      @       @      @      P@      =@                      @      @              ,@              @                              @     �J@     �B@      @      �?      @      2@      0@                      �?       @              5@       @      *@               @                      B@     �E@              �?      �?      G@      *@                       @      @              $@      �?      *@              �?              @      "@      "@      �?      @      @      4@      3@               @              �?      �?       @              @                                      @      �?                      �?      @                                                       @      �?      $@              �?              @      @       @      �?      @      @      1@      3@               @              �?      �?     �U@      .@      I@      $@      @      �?      .@      X@      ]@      "@      *@      B@     @V@     �R@      @      0@       @      8@      @     �D@       @      B@       @       @      �?      @      M@     �M@      @      @      &@      :@      A@              @      @      @       @      8@      @      *@              �?      �?      @      E@     �H@      @      @      $@      .@      ;@              @       @      @       @      8@      �?      $@                               @     �C@      H@      �?       @      @      (@      8@              @      �?       @      �?               @      @              �?      �?      �?      @      �?      @      @      @      @      @               @      �?       @      �?      1@      @      7@       @      �?                      0@      $@                      �?      &@      @                       @                      (@      @       @              �?                      ,@      @                              @      @                                              @      �?      .@       @                               @      @                      �?      @       @                       @                      G@      @      ,@       @       @              (@      C@     �L@      @      @      9@     �O@      D@      @      "@      @      4@       @     �A@      @      @       @      �?              @     �@@      F@              @      0@      ?@      8@              @      �?      *@       @      2@      @      @                              @      >@      :@              @      $@      =@      2@              @              @      �?      1@      @      �?       @      �?              �?      @      2@               @      @       @      @              @      �?      @      �?      &@      �?      "@              �?              @      @      *@      @              "@      @@      0@      @      @      @      @              @               @                              �?      @      &@      @              @      8@      ,@      @       @              @              @      �?      @              �?              @      �?       @      �?               @       @       @              �?      @      @             �A@      $@      6@              �?              (@      G@     �A@       @       @      0@     �I@     �C@       @      $@      �?      &@      @      0@       @       @              �?                      @      "@               @       @      4@      @                              @      @      @      �?      �?              �?                      @      @                              "@                                      @              �?              �?              �?                      @                                      "@                                      �?              @      �?                                              @      @                                                                      @              "@      �?      �?                                              @               @       @      &@      @                                      @      @              �?                                              @               @      @      @      @                                               @              �?                                               @               @      @       @      @                                              �?                                                              @                              @                                                      @      �?                                                                              @      @       @                                      @      @                                                                                      @      @       @                                      @       @      �?                                                                               @      @                                                      3@       @      4@                              (@     �C@      :@       @      @       @      ?@     �@@       @      $@      �?      @      �?      @              ,@                              �?      ;@      $@                       @      (@      �?              �?              �?      �?       @              �?                                      1@      @                              @                      �?                                              �?                                      &@      �?                               @                                                       @                                                      @      @                              @                      �?                               @              *@                              �?      $@      @                       @      @      �?                              �?      �?      �?              (@                              �?       @                                       @                                                      �?              �?                                       @      @                       @      @      �?                              �?      �?      .@       @      @                              &@      (@      0@       @      @      @      3@      @@       @      "@      �?      @              @                                                      @       @              @      �?              @                              �?              @                                                      �?      �?              @      �?              @                              �?                                                                      @      @                                       @                                              &@       @      @                              &@       @       @       @              @      3@      ;@       @      "@      �?      @              &@      @      @                              @       @       @       @              @      2@      :@      �?      "@      �?      @                      @       @                              @                                              �?      �?      �?                                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�ߚchG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         @                     @=h����?�	           ��@       !                    �?w�3SV�?�           t�@                            �?�X�u�o�?           ȓ@                          �1@��f��?S           �@                           @z�˼��?c             e@                           @�kn��?R            `a@������������������������       ����Z��?>            �Z@������������������������       ���$d�?            �@@	       
                    �?|�j�Y��?             >@������������������������       �R���Q�?             $@������������������������       ��z�G��?	             4@                          �7@r?kF���?�           ��@                           �?��}&���?F           8�@������������������������       �E~����?o            �e@������������������������       ���Ųl�?�            �u@                          �9@A���]��?�            q@������������������������       �q T���?B            �\@������������������������       �z&dx)�?h            �c@                           @-Q�XX9�?�            s@                          �5@R�5�`��?P             _@                           @Vp���<�?)            @P@������������������������       ��W�!l��?            �E@������������������������       �b���i��?             6@                           �?�r��bn�?'            �M@������������������������       ��7�A�?             6@������������������������       ��,y8"q�?            �B@                           @NE�Z��?u            �f@                          �3@Dܗ�V�?T            �`@������������������������       �������?2            @S@������������������������       ��pyU���?"            �K@                            @f�nOwA�?!            �H@������������������������       �9��8���?             >@������������������������       �窷uJ��?             3@"       1                     �?���p��?�            �@#       *                    �?�������?�           ̑@$       '                   �6@�Y�T�O�?�            �y@%       &                    �?rʃ����?�            @q@������������������������       �_���l�?�            `m@������������������������       �ĭ[F�?            �D@(       )                    �?[�FR"��?N            �`@������������������������       ��Q��Q��?@            �Y@������������������������       ��q�q�?             >@+       .                     �?��/�?�           ؆@,       -                    �?�%�!�?            z@������������������������       �ؚ�:�^�?�            `h@������������������������       ��c�A%�?�            �k@/       0                   �9@RKfw���?�            �s@������������������������       ��jf8D�?�            �o@������������������������       �\&p��?(             O@2       9                   �5@�'�"�s�?�            Pu@3       6                    @���|�O�?w             g@4       5                    �?m�w6�;�?             �G@������������������������       �0�����?             2@������������������������       �c��gS~�?             =@7       8                    @֔�4��?W            @a@������������������������       �Y�C��?H             \@������������������������       ��T�6|��?             :@:       =                    @qq>]6��?d            �c@;       <                    @M�4M�4�?R            �_@������������������������       �����$}�?>            @W@������������������������       ���@�S��?            �@@>       ?                    @t�@�t�?             >@������������������������       �     ��?
             0@������������������������       �����>4�?             ,@A       `                    �?)7~���?�           <�@B       Q                    �?~k ��I�?J           ��@C       J                    �?s�M>��?�            @r@D       G                   �4@)v8���?7            @V@E       F                   �1@�t��hj�?            �H@������������������������       ��}�+r��?             3@������������������������       �|�j�Y��?             >@H       I                    @\���(\�?             D@������������������������       ������?             ?@������������������������       ���"e���?             "@K       N                    �??�b��x�?|            `i@L       M                   �3@���(A�?$            �I@������������������������       �*L�9��?	             &@������������������������       ��(\����?             D@O       P                    @��KM�]�?X             c@������������������������       �     x�?'             P@������������������������       ��T�x?r�?1             V@R       Y                    �?���v��?�            �m@S       V                    @&ޏ��k�?9             V@T       U                   �7@���W��?            �A@������������������������       �|гY���?             9@������������������������       ���Q��?             $@W       X                   �2@N���9�?"            �J@������������������������       ��z6�>�?             9@������������������������       ����S�r�?             <@Z       ]                    @�f�^��?^            �b@[       \                   �:@7exwX�?<            @X@������������������������       �b]�N��?5            �T@������������������������       �4և����?             ,@^       _                    @[$��m�?"             J@������������������������       ��������?             D@������������������������       �r�q��?             (@a       n                   �9@�ٵ�ZD�?�           ��@b       i                    @�ӡ*��?Z           �@c       f                    @F5y9h��?           0x@d       e                    @Pݻ��?�            s@������������������������       ��eڄn��?�            �p@������������������������       �v�[��?            �A@g       h                    @������?9            �T@������������������������       �ԭ�a�2�?2             R@������������������������       ����Q��?             $@j       m                    @��%��1�?R            �_@k       l                   �6@�����?8            �V@������������������������       �q=	�?.            @S@������������������������       ���WV��?
             *@������������������������       ��2�tk~�?             B@o       v                   �@@z�m�(�?T            @_@p       s                    �?f� �o��?I            �Z@q       r                    �?9��8���?2             R@������������������������       �j�����?             3@������������������������       ���>����?#            �J@t       u                    @�.k���?             A@������������������������       �]��N��?             3@������������������������       ��������?             .@������������������������       ���a_j�?             3@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       �|@     �Q@     `v@      E@     �Q@      :@     @S@     X�@     `�@      M@     @Z@     @_@     ��@     �y@      1@      P@      J@     `b@      O@      t@     �D@     `l@      <@     �E@      ,@      K@      |@     `|@      D@      Q@     @T@     @{@     `q@       @     �F@      ?@      W@      B@      f@      3@     @S@      @      ,@              $@     0p@      p@      $@      9@      ;@     �i@     �\@              *@      $@      ;@      0@     `b@      0@     �M@      @      @              $@     @d@     @i@      @      5@      8@     �c@     @U@              $@      "@      8@      0@      6@              @                               @     �P@      G@               @      @      5@      �?                              �?              0@              @                               @     �N@      B@               @      �?      .@      �?                              �?              .@                                               @      G@      >@               @      �?       @      �?                              �?              �?              @                                      .@      @                              @                                                      @              �?                                      @      $@                       @      @                                                                      �?                                      @      @                       @      �?                                                      @                                                       @      @                              @                                                     @_@      0@      K@      @      @               @      X@     �c@      @      3@      5@      a@      U@              $@      "@      7@      0@     �X@      @      <@      �?      @              @     @T@      \@      @      &@      *@     �Z@     �A@              @      @      @      @      @@      �?      0@              @               @      1@      6@               @      @     �H@      "@              �?              �?      @     �P@      @      (@      �?                       @      P@     �V@      @      @      @      M@      :@              @      @      @      �?      :@      &@      :@      @       @              @      .@      F@      @       @       @      >@     �H@              @      @      2@      (@      @              1@                               @      @      7@              @      @      &@      >@              @      �?      @              3@      &@      "@      @       @               @      &@      5@      @      @      @      3@      3@              �?      @      &@      (@      >@      @      2@               @                     @X@      K@      @      @      @     �G@      >@              @      �?      @              0@       @      &@              @                      ;@      3@               @      �?      2@      1@              @      �?      @              @      �?      @                                      8@      &@               @              @      &@                              @              @              @                                      .@      "@               @               @      @                              @              �?      �?                                              "@       @                               @      @                                              $@      �?       @              @                      @       @                      �?      ,@      @              @      �?                      @      �?       @                                              @                              @                      @                              @              @              @                      @      @                      �?       @      @                      �?                      ,@      �?      @              @                     �Q@     �A@      @       @       @      =@      *@                                              @              @                                     �N@      5@      @       @       @      7@      &@                                               @                                                      F@      .@      @                      &@      �?                                              @              @                                      1@      @               @       @      (@      $@                                              "@      �?      @              @                      "@      ,@                              @       @                                              "@      �?      �?                                      @      "@                              @       @                                                              @              @                      @      @                               @                                                     �a@      6@     �b@      6@      =@      ,@      F@     �g@     �h@      >@     �E@      K@     �l@     `d@       @      @@      5@     @P@      4@     @[@      *@     @_@      0@      ;@      (@      @@      `@     �c@      5@      A@     �D@     �d@     �a@      @      <@      3@      I@      0@      K@      �?      :@              @      @      0@      I@     �M@       @      .@       @     @Q@     �O@      @      @      @      (@      @      F@      �?      &@               @      @      "@     �H@     �J@              "@      @     �D@      A@              �?      @      @      @     �B@              "@               @      @      @      F@     �I@              @      @      A@      8@              �?      @      @      @      @      �?       @                              @      @       @               @              @      $@                                              $@              .@              @              @      �?      @       @      @      @      <@      =@      @       @      @      @      �?       @              "@              @              @      �?      @      @      @      @      0@      5@      @       @       @      @      �?       @              @                                                      �?                      (@       @                      �?                     �K@      (@     �X@      0@      5@       @      0@     �S@     @X@      *@      3@     �@@     �X@     @S@              9@      *@      C@      (@      :@       @      L@      ,@       @      @       @     �G@      E@       @      *@      4@      N@     �G@              (@      "@      8@      @      (@      @      =@       @      @      @      @      @      "@      @      *@      $@      9@      :@              $@      @       @      @      ,@       @      ;@      @      �?              @      E@     �@@      @              $@     �A@      5@               @      @      0@       @      =@      @     �E@       @      *@      �?       @      @@     �K@      @      @      *@      C@      >@              *@      @      ,@      @      <@      @     �B@              @              @      >@     �I@      @      @      &@      >@      6@              @      @      *@      �?      �?      �?      @       @      "@      �?       @       @      @       @      �?       @       @       @              @      �?      �?      @      A@      "@      9@      @       @       @      (@      O@      E@      "@      "@      *@      P@      7@      @      @       @      .@      @      6@      @      (@              �?              @      K@      =@      �?              @     �C@      &@                              @       @       @              &@              �?              @      @      @                      �?      @      @                                              @                                               @      @       @                              @      @                                              @              &@              �?               @      @      @                      �?      @      �?                                              ,@      @      �?                                      H@      8@      �?               @      @@      @                              @       @       @      @      �?                                     �F@      7@      �?               @      7@      @                              @              @                                                      @      �?                              "@      @                              �?       @      (@      @      *@      @      �?       @       @       @      *@       @      "@      $@      9@      (@      @      @       @      &@       @      @      @      @      @      �?       @       @      @      *@      @      "@       @      9@      $@      @      @       @      "@       @      @      @      @      @      �?       @       @      @      (@       @       @      @      7@       @      @      @       @       @      �?      @                      �?                      @              �?      @      �?      @       @       @      �?                      @      �?      @       @      $@       @                              �?              @               @               @              �?               @              @      �?      @       @                              �?              @                                              �?              �?              �?      �?      @                                                                       @               @                              �?             `a@      >@     ``@      ,@      <@      (@      7@     @Z@     �`@      2@     �B@      F@      h@     @`@      "@      3@      5@     �K@      :@      N@      @     �L@       @       @      @       @      Q@      T@              .@      .@     �Y@     �J@      �?      &@      "@      6@      @      ?@      �?      @@      �?      @      @      @      :@     �D@              @      (@     �M@      <@      �?       @      "@      .@      @      "@              $@                       @              .@      .@               @      @      .@       @              @               @      @       @               @                                      ,@       @                      �?      @      @              �?               @              @               @                                      @      @                      �?      @                                                      @                                                      &@      @                              @      @              �?               @              �?               @                       @              �?      @               @      @      "@      �?              @                      @      �?               @                       @                      @               @      �?      @                      @                       @                                                              �?                               @      @      �?                                      �?      6@      �?      6@      �?      @      �?      @      &@      :@              @       @      F@      4@      �?      @      "@      *@      @      .@      �?      @               @                              @              �?              $@      "@      �?                      @              �?      �?                                                       @                                      @                              @              ,@              @               @                              �?              �?              $@      @      �?                       @              @              3@      �?      @      �?      @      &@      7@              @       @      A@      &@              @      "@      @      @      @              $@               @               @      @      (@              �?      @      @      @              @      @              �?      @              "@      �?      @      �?      @      @      &@              @       @      ;@      @              �?      @      @       @      =@      @      9@      �?      �?      �?      @      E@     �C@               @      @     �E@      9@              @              @      �?      *@      @      (@              �?      �?              $@      .@                              .@      .@              �?              �?              @       @       @                      �?              @      @                              @      "@              �?                              @       @                              �?              @      @                              @      @                                                               @                                                                               @      @              �?                               @       @      $@              �?                      @      &@                              "@      @                              �?              @              $@                                      @      @                               @                                                      @       @                      �?                       @      @                              @      @                              �?              0@       @      *@      �?                      @      @@      8@               @      @      <@      $@               @              @      �?      "@              @      �?                              :@      2@              @              6@      @               @              @      �?      "@              @      �?                              :@      *@              @              4@      @                               @      �?                      �?                                              @              @               @                       @              �?              @       @       @                              @      @      @              �?      @      @      @                              @              @      �?       @                                      @      @              �?      @      @      @                              �?                      �?                                      @              @                              �?       @                               @             �S@      7@     �R@      (@      4@       @      .@     �B@      K@      2@      6@      =@     �V@     @S@       @       @      (@     �@@      3@     @Q@      2@     @P@       @      ,@      �?       @     �A@     �H@      *@      2@      6@     @U@      P@      �?      @       @      8@       @     �K@      .@     �H@      @      *@      �?      @      :@      E@      @      &@      1@      R@     �F@              @      @      ,@      @      E@      &@     �C@      @      &@      �?      @      7@      C@      @      &@      (@      I@      C@              @      @      "@      �?      A@      &@      C@      @      &@      �?      �?      ,@      B@      @      &@      (@      G@     �@@               @      �?      "@      �?       @              �?                               @      "@       @                              @      @              �?      @                      *@      @      $@               @              �?      @      @      @              @      6@      @                      �?      @       @      (@      @      $@               @              �?       @      @      @              @      .@      @                      �?      @       @      �?      �?                                              �?                                      @                                                      ,@      @      0@      @      �?              @      "@      @      @      @      @      *@      3@      �?              @      $@      @      $@      @      *@       @      �?               @      @      @      @      @      @      "@      *@                      @      $@      @      "@      @      @       @      �?               @      @      @      @      @       @      "@      (@                      @      $@      @      �?               @                                                              �?      �?              �?                                      �?      @              @      �?                       @      @      @      �?      @       @      @      @      �?                                      $@      @      "@      @      @      @      @       @      @      @      @      @      @      *@      @      @      @      "@      &@      $@      @      "@      @      @      @      @       @      @      @       @      @      @      *@       @      @       @      "@       @      @      @       @      @       @      @      @              @       @       @      @      @      @       @      @       @      @      @       @       @       @              �?                                      �?              �?      �?       @              @      �?       @      �?      @       @      @      @      �?      @      @              @      �?       @       @       @      @       @       @      �?      @      @      @      �?      �?               @              @       @      �?      @                       @       @                              @       @      @      �?                       @                              �?      @                              @                               @       @                      �?                              @       @                                       @      @                               @                                               @      �?                                       @      @                      @               @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�P�)hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKuhnh4h7K ��h9��R�(KKu��hu�B�         8                   �3@^J�Ф��?�	           ��@                           �?r�/�Z�?q           ̕@                           �?�&e����?           p{@                           @1��*�?w             i@                           �?���V��?J            @_@                           �?J{�/L��?!             I@������������������������       �"�u�)��?            �B@������������������������       �����W�?             *@	       
                    �?����9�?)            �R@������������������������       �� 5���?            �@@������������������������       �>��t�?             E@                          �1@�h�*$��?-             S@                          �0@,�Œ_,�?             >@������������������������       ��h$���?             .@������������������������       ��A��S�?	             .@                           �?�;5r��?             G@������������������������       �؉�؉��?             :@������������������������       �H�z�G�?             4@                            @��c!��?�            �m@                          �2@�@�����?S            �_@                            �?�3�����??            @X@������������������������       �m��
I��?3            @T@������������������������       �      �?             0@                           �?v��`��?             =@������������������������       �
ц�s�?             *@������������������������       �     @�?             0@                          �0@�)x9��?K             \@������������������������       ����Դ�?	             3@                           �?%<�����?B            @W@������������������������       �:m���?             >@������������������������       �ğӯZ��?.            �O@        +                   �1@s7,�8R�?\           ��@!       (                    @v0f����?            {@"       %                    �?_�kt6��?�            �y@#       $                     @q��$�?�            �k@������������������������       ���3��?l            �e@������������������������       ��_�a	��?            �H@&       '                   �0@�� ���?y            `g@������������������������       �#]�6�?(            �N@������������������������       �d���M�?Q            �_@)       *                    �?���H�~�?             7@������������������������       �*L�9��?             &@������������������������       �9��8���?             (@,       3                    @"�OA6�?N           `�@-       0                    �?���ĮH�?3           `~@.       /                   �2@���.��?�            �j@������������������������       ��J��s��?F            �\@������������������������       ���ͪ���?<             Y@1       2                    @pB�M�?�             q@������������������������       �>?�Ï�?y            `g@������������������������       �w�m�d��?8            @U@4       5                    �?�8	���?             C@������������������������       �X�3�R�?             3@6       7                   �2@^Cy�5�?             3@������������������������       �j�V���?             &@������������������������       �      �?              @9       X                    �?vq7�h��?A           ��@:       I                    �?L7�%,�?           �@;       B                    �?췿E��?           `{@<       ?                   �4@9��҉�?m            �d@=       >                     �?\")�i��?             7@������������������������       ����Q��?             $@������������������������       ��T�6|��?             *@@       A                    @z�:+��?^            �a@������������������������       �������?J             \@������������������������       ����;\I�?             =@C       F                   �<@C�ş���?�             q@D       E                   �7@�TF�Rn�?�             m@������������������������       �y�����?S             a@������������������������       ���a����?9            @X@G       H                   �?@�����?            �D@������������������������       ��+\&p�?             ?@������������������������       ��G�z��?             $@J       Q                    �?lS��~F�?�           `�@K       N                   �7@�9!x��?�            0s@L       M                   �5@>�&�?_            �b@������������������������       ��5τ���?7            �W@������������������������       ��$I�$I�?(             L@O       P                   �9@ԐO{���?`            �c@������������������������       �b�B���?&            �P@������������������������       ���S���?:            �V@R       U                     @�HtfQ�?6           �}@S       T                     �?\�����?�            �n@������������������������       �Z�#L��?d            `b@������������������������       ��xFƑ��?B            �X@V       W                   �@@?���b�?�            `l@������������������������       �Y�I�:�?�            @k@������������������������       ���E���?             "@Y       f                    �?��5�_�?;           P�@Z       a                    @K�a��?�            �x@[       ^                    @El<�1��?�            �j@\       ]                    �?X��%��?x            �e@������������������������       �Ǽ�����?A            �Y@������������������������       ��tk~X��?7             R@_       `                   �5@��a_j�?             C@������������������������       �������?             *@������������������������       ���+e��?             9@b       e                     @�b���f�?k             g@c       d                   �;@D�=��?\            �c@������������������������       �����?S            `b@������������������������       �r�q��?	             (@������������������������       ��<pƵ�?             :@g       n                   �:@�����{�??           8�@h       k                   �5@������?�           p�@i       j                   �4@���m��?�            �s@������������������������       � SoU_��?h            �d@������������������������       ��Rro-�?[            `c@l       m                    �?#|ӂrT�?           �x@������������������������       ���8��8�?             8@������������������������       ��O��,O�?�            pw@o       r                    �?%>L�S#�?u             g@p       q                     �?Q�a�r��?*             N@������������������������       ����(\��?             4@������������������������       �333333�?             D@s       t                     @�D�$�?K            @_@������������������������       ���u>�?7            �V@������������������������       ����:��?            �A@�t�bh�h4h7K ��h9��R�(KKuKK��h��BxE       �y@      W@     �t@      C@     �T@      ?@     �V@     ��@     ��@     �L@     �P@     @d@     p�@     �|@      $@      L@      L@     @[@     �J@     �e@      2@     @V@      @      $@              &@     �t@     �q@      @      $@     �E@      m@     @]@              $@      @      A@       @     �Q@      @     �A@      �?      "@              @      M@     @R@      @      @      ,@     @V@      F@              @       @      2@      @      :@              "@                              @     �B@     �C@      @               @      F@      3@              @               @       @      1@              �?                              @      =@      8@      �?              @      8@      "@              �?              @       @      (@                                                      "@      @      �?              @      "@      @              �?                              (@                                                      @      @      �?              @      @      @              �?                                                                                      @      �?                      �?      @       @                                              @              �?                              @      4@      1@                       @      .@      @                              @       @      @                                                      @      @                              $@      @                              @               @              �?                              @      .@      (@                       @      @                                               @      "@               @                                       @      .@       @              �?      4@      $@               @              �?              �?              @                                      @      "@                              @      @                                                              @                                      �?      @                               @      @                                              �?              @                                       @      @                               @                                                       @              �?                                      @      @       @              �?      0@      @               @              �?              @              �?                                      �?      @       @                      $@      @                                              @                                                      @      �?                      �?      @                       @              �?              F@      @      :@      �?      "@              �?      5@      A@       @      @      @     �F@      9@              �?       @      $@      @      5@              .@      �?      @              �?      (@      9@              �?      @      7@      $@                              @       @      2@              @              @              �?      $@      6@                      @      6@       @                              @       @      ,@              @              @                      @      3@                      @      4@       @                              @       @      @                                              �?      @      @                      �?       @                                                      @               @      �?                               @      @              �?              �?       @                               @                              @                                       @       @                                       @                                              @              �?      �?                                      �?              �?              �?      @                               @              7@      @      &@              @                      "@      "@       @      @       @      6@      .@              �?       @      @      �?      @      @                                              @      �?                               @      @                                              2@              &@              @                      @       @       @      @       @      4@      (@              �?       @      @      �?      &@              @               @                      �?      @              �?              @      �?                       @      �?      �?      @               @              @                      @      @       @       @       @      0@      &@              �?               @             �Y@      ,@      K@      @      �?              @     @q@     �j@       @      @      =@      b@     @R@              @      @      0@      @     �H@      @      (@                              @     �b@     �[@              �?      0@     @P@      4@              �?              @             �F@      @      (@                              @      b@      [@              �?      .@      O@      ,@              �?              �?              :@      �?      @                              �?     �W@      K@                      @     �@@       @                                              *@      �?      @                              �?     �U@      D@                      @      7@      �?                                              *@               @                                      "@      ,@                              $@      �?                                              3@       @      @                               @     �H@      K@              �?      &@      =@      (@              �?              �?              (@               @                                      4@      $@                       @      &@      @                                              @       @      @                               @      =@      F@              �?      "@      2@       @              �?              �?              @                                                      @       @                      �?      @      @                              @               @                                                      @      �?                      �?      @                                                       @                                                              �?                                      @                              @              K@      &@      E@      @      �?              @      `@     �Y@       @      @      *@     �S@     �J@              @      @      (@      @     �I@      &@      D@      @                      @     �^@     �V@       @      @      *@     �P@      J@              @      @      (@      @      :@              7@       @                       @      H@     �D@                       @      >@      A@              @       @              �?      ,@              0@                               @      =@      4@                              3@      (@               @                              (@              @       @                              3@      5@                       @      &@      6@              �?       @              �?      9@      &@      1@      @                       @     �R@     �H@       @      @      &@      B@      2@               @       @      (@       @      0@      &@      @       @                       @     �N@      @@       @      @      @      7@      "@                      �?      $@       @      "@              $@       @                              *@      1@               @      @      *@      "@               @      �?       @              @               @              �?                      @      (@                              *@      �?                                               @              �?                                      @      �?                              &@                                                      �?              �?              �?                       @      &@                               @      �?                                                              �?                                       @       @                                                                                      �?                              �?                              @                               @      �?                                             �m@     �R@     �n@      ?@     @R@      ?@      T@      j@     �s@      I@     �L@     �]@     Pz@     �u@      $@      G@      I@     �R@     �F@      ]@      E@     @b@      1@     �I@      8@      H@      D@      [@      6@      E@     @R@      g@     �e@      @      :@      @@      C@      ?@      H@      (@      D@              1@      @      .@      *@     �L@       @      1@      ;@     @W@      H@              @      $@      &@      (@      4@      @      1@              @       @      @      @     �@@      @      @      @     �D@      &@              @       @       @      @      @                               @                      @      @                              "@                                                      �?                                                      �?      �?                              @                                                       @                               @                      @      @                               @                                                      1@      @      1@              �?       @      @      �?      =@      @      @      @      @@      &@              @       @       @      @      ,@      @      1@              �?       @      @      �?      ;@      @      @      @      3@      @              @       @       @       @      @                                              �?               @              @              *@      @                                      �?      <@      @      7@              ,@      �?      &@      @      8@      @      &@      8@      J@     �B@              @       @      "@      "@      <@      @      3@               @      �?      @      @      7@      @      @      0@      I@     �A@              @      @       @       @      *@      @      ,@              @              @      @      6@      @      @       @     �@@      (@              �?      @      @      @      .@      �?      @              @      �?              @      �?       @      @       @      1@      7@              @              @      @              @      @              @              @              �?              @       @       @       @                       @      �?      �?              @       @              @              @              �?                      @       @       @                       @              �?                       @              �?                                              @       @                                              �?              Q@      >@     �Z@      1@      A@      5@     �@@      ;@     �I@      ,@      9@      G@      W@      _@      @      3@      6@      ;@      3@     �A@      &@     �E@      �?      &@              2@      2@      8@              &@      0@     �F@      E@       @      @      &@       @      @      4@              8@              @              @      2@       @              @      $@      >@      .@      �?      @              @      �?      .@              $@              @                      .@       @              @       @      2@      &@               @              @      �?      @              ,@               @              @      @      @              �?       @      (@      @      �?      �?                              .@      &@      3@      �?      @              *@              0@              @      @      .@      ;@      �?       @      &@      @      @      @              @                              $@              $@                      @      @      3@               @      �?              @      "@      &@      ,@      �?      @              @              @              @      �?      $@       @      �?              $@      @       @     �@@      3@     �O@      0@      7@      5@      .@      "@      ;@      ,@      ,@      >@     �G@     �T@      @      ,@      &@      3@      *@      ;@      @      >@      @      $@              @      @      $@       @      @      0@      ;@      I@              &@      @      *@      @      2@      @      6@      @      @               @      �?      "@      @      @      @      .@      <@              @      @      @      @      "@               @       @      @              @      @      �?      @      �?      $@      (@      6@              @       @      @      @      @      (@     �@@      $@      *@      5@      "@       @      1@      @      "@      ,@      4@      @@      @      @      @      @      @      @      (@     �@@      $@      (@      5@      "@       @      1@      @       @      ,@      4@      @@      �?      @      @      @       @                                      �?                                              �?                               @                              @     �^@      @@     �X@      ,@      6@      @      @@      e@     `j@      <@      .@      G@     �m@     �e@      @      4@      2@     �B@      ,@     �B@      "@      @@              @      @      @     �R@      W@      @      @      &@     �H@      J@              &@              @      @      5@      @      8@               @      @       @      4@     �I@      @      @      "@      ?@      =@              @               @       @      3@       @      2@               @      @       @      2@      E@      @              "@      5@      :@              @              �?       @      (@       @      &@              �?       @              @      ?@                      @      ,@      0@              �?                              @              @              �?       @       @      &@      &@      @              @      @      $@              @              �?       @       @      �?      @                                       @      "@              @              $@      @                              �?                              @                                       @      @               @                      �?                                               @      �?      @                                              @               @              $@       @                              �?              0@      @       @              �?              �?     �K@     �D@      @               @      2@      7@              @               @       @      0@      @       @                              �?      K@      @@      @              �?      *@      1@              @               @       @      0@       @       @                              �?      K@      ;@      @              �?      &@      *@              @               @       @              �?                                                      @                               @      @                                                      @                      �?                      �?      "@                      �?      @      @                                             �U@      7@     �P@      ,@      3@      @      =@     �W@     �]@      5@      &@     �A@     `g@      ^@      @      "@      2@     �@@      $@     @Q@      *@      J@      (@      &@              7@     �U@      Z@      $@      "@      :@     �d@     @U@      @      @      $@      :@      @     �A@      @      7@      @      @              $@      C@     �N@      @      @       @      S@      =@               @      @      *@      @      &@      @      $@      @       @              @      0@      B@               @      @     �A@      6@               @      @       @       @      8@      �?      *@              �?              @      6@      9@      @      �?      @     �D@      @                              @       @      A@      "@      =@      "@       @              *@      H@     �E@      @      @      2@     @V@      L@      @      @      @      *@      @      @              @      @                               @                                      @                              �?                      <@      "@      9@      @       @              *@      G@     �E@      @      @      2@     �T@      L@      @      @      @      *@      @      1@      $@      .@       @       @      @      @       @      .@      &@       @      "@      6@     �A@       @       @       @      @      @      @      @      @      �?       @                      @       @      @       @      �?      (@      (@                              �?      �?      @      @      �?                                       @               @                      �?      @                              �?              �?       @      @      �?       @                      @       @      �?       @      �?      &@       @                                      �?      (@      @      &@      �?      @      @      @      �?      *@       @               @      $@      7@       @       @       @      @       @      (@      �?      &@      �?      @      @      @              "@       @              @      @       @               @       @      @      �?               @                      �?              @      �?      @                      @      @      .@       @                              �?�t�bub�2'     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��=RhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         :                   �5@�:F���?�	           ��@                           �?퉴����?:           ؠ@                           @F��zM�?�           ��@                           �?���@�?�           �@                           �?��GZ��?�            �q@                            �?UeEaM�?P             `@������������������������       �b|�MA<�?1            �S@������������������������       ��3�B�Q�?            �I@	       
                     �?����?Z             c@������������������������       ���^�?             I@������������������������       �_���'Z�?A            �Y@                           @��j[�H�?           �|@                           �?8H�l�S�?�            `w@������������������������       ��F�5��?W             c@������������������������       ���Uր�?�            �k@                            �?���g��?4            �T@������������������������       ��ˠT�?             6@������������������������       ��-o0@��?&            �N@                           @�Q�}e��?#             J@                          �2@���h�u�?            �D@                           �?�q�q�?             2@������������������������       �}��7�?             &@������������������������       �������?             @                             @#8̺�8�?             7@������������������������       �9��8���?             (@������������������������       �*L�9��?             &@������������������������       �*L�9��?             &@       +                    �?J�$����?T           X�@       $                    @7^�ֻ��?�           8�@       !                    @S֔5eM�?k            �e@                           �3@�w,C��?S            @a@������������������������       �~KfK!��?4            �V@������������������������       ��s�æ��?            �G@"       #                   �2@،A��_�?             A@������������������������       �O��E��?             2@������������������������       �     ��?	             0@%       (                     �?'LzӍ��?P           ؀@&       '                    @��[���?P            @_@������������������������       ������z�?>             X@������������������������       ���`���?             =@)       *                    @�UK��?            �y@������������������������       ��������?�             x@������������������������       ���(\���?             >@,       3                    @�f�b��?�           x�@-       0                    @ΰ� �?�            �u@.       /                    �?.@Rdv��?�            �o@������������������������       �����8�?c            �d@������������������������       ��t���?4            �V@1       2                    �?F/.�?7            @V@������������������������       �*;L]�?#             N@������������������������       ���-�?             =@4       7                    @wIT���?�            ps@5       6                    @��)V��?:            @V@������������������������       �{�G�z�?             4@������������������������       ���JÝ�?,            @Q@8       9                   �4@�����?�            �k@������������������������       ���]�M��?~             h@������������������������       ������?             =@;       V                    �?���_F�?]           t�@<       K                   �>@�����?"           �@=       D                     �?
,\&U�?�           ��@>       A                    @����G�?            Py@?       @                    �?#�(�B�?�            �p@������������������������       ����;è�??            @Z@������������������������       �Oh�/�?`            �c@B       C                    �?$~\	���?a            �a@������������������������       �S��d��?(             N@������������������������       �)��I�?9            @T@E       H                    �?�q�4�&�?�            �u@F       G                     @UUUUU��?B             X@������������������������       �V�Lt�<�?             3@������������������������       ����n��?4            @S@I       J                    @��R���?�            `o@������������������������       ��J����?n             f@������������������������       �KX̦��?1            �R@L       O                     �?J������?A            @[@M       N                    @N贁N�?             >@������������������������       ��;��KM�?             3@������������������������       �t�E]t�?             &@P       S                    @ ��Aa�?/            �S@Q       R                    @v��4��?            �A@������������������������       ��~Q$���?             1@������������������������       ����^B{�?             2@T       U                   @@@�4_�g�?             F@������������������������       �g\�5�?             *@������������������������       �@Q�f?��?             ?@W       f                    �?������?;            �@X       _                    �?��e����?�            0y@Y       \                   �9@�o�tH��?R            �a@Z       [                   �7@�k����?<            @Z@������������������������       �:m���?#             N@������������������������       �D��OS��?            �F@]       ^                    @��Kh/�?             B@������������������������       �      �?             (@������������������������       �9��8���?             8@`       c                    @~<!�$�?�            `p@a       b                     �?.��d��?'            @P@������������������������       �0�N�?            �E@������������������������       �fP*L��?             6@d       e                   �8@F�\wy��?            �h@������������������������       ��B�c�I�?B            @Y@������������������������       �r�qW�?=             X@g       n                     @���
a��?C           �~@h       k                    @&�p���?
           �y@i       j                    @��I�j��?�            �s@������������������������       �������?�            �p@������������������������       ��C��2(�?             F@l       m                   �8@r�qw�?A             X@������������������������       �I��D��?#             K@������������������������       ��0�0�?             E@o       r                   �>@Il�py��?9            �T@p       q                    @L���?3            @R@������������������������       ��>���T�?            �A@������������������������       ��Ł�r��?             C@������������������������       �R���Q�?             $@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       @|@     @X@     0u@      D@      T@      =@     @U@     Ѐ@     `�@      F@     �U@     @b@     ��@     �{@      (@      M@     �N@      `@      H@      r@      ?@     @e@      @      9@      @     �@@      z@      x@      $@      <@      N@      x@     `j@              3@      ,@     �K@      &@     �\@      1@     �T@      �?      0@      @      ,@     @W@      Z@      @      2@      >@     �b@     �T@              @       @      C@      @     �Y@      1@     �Q@      �?      .@      @      ,@     @W@      Y@      @      0@      ;@      b@     �R@              @       @      A@      @      =@      @      .@              �?               @     �F@     �D@      @      @      ,@     �P@      8@              @      @      (@      @      .@              @                              @      B@      ;@               @      @      8@      "@              @              �?      �?       @               @                              @      5@      (@                      @      3@      @                                      �?      @              �?                                      .@      .@               @              @       @              @              �?              ,@      @      (@              �?              @      "@      ,@      @      @      $@      E@      .@                      @      &@       @       @      @      @                              @      @      @                      @      4@                                      @              (@      �?      @              �?                      @      $@      @      @      @      6@      .@                      @      @       @     @R@      (@      L@      �?      ,@      @      @      H@     �M@      �?      "@      *@     �S@     �I@              @      @      6@      @      Q@      &@     �C@      �?      (@      @      @     �A@     �I@      �?       @       @      M@     �E@              @      @      4@      @      <@      @       @              @                      7@      7@              �?       @      >@      0@              �?              $@              D@      @      ?@      �?      @      @      @      (@      <@      �?      @      @      <@      ;@               @      @      $@      @      @      �?      1@               @                      *@       @              �?      @      5@       @                               @                              "@                                       @      @                      �?      @       @                              �?              @      �?       @               @                      &@      @              �?      @      2@      @                              �?              *@              (@              �?                              @               @      @      @      @              �?              @      �?      "@              (@                                              @               @      @       @      @              �?              @              @              @                                                              �?              �?      �?              �?              �?              @              @                                                              �?              �?                                      �?              �?              @                                                                                      �?              �?                              @              @                                              @              �?      @      �?      @                              @              @              �?                                              @              �?                       @                              �?                              @                                                                      @      �?      �?                               @              @                              �?                                                               @      @                                      �?     �e@      ,@     �U@      @      "@      @      3@     0t@     �q@      @      $@      >@     �m@      `@              (@      @      1@      @     �T@       @     �E@               @       @       @      h@     `e@      @      @      @     �`@     �G@              �?              @              4@       @      "@                       @              @@      M@       @               @     �A@      "@                              �?              1@       @      "@                       @              ?@      D@                      �?      :@      "@                              �?              &@              @                                      =@      8@                      �?      1@      @                                              @       @      @                       @               @      0@                              "@      @                              �?              @                                                      �?      2@       @              �?      "@                                                      �?                                                      �?      (@       @                       @                                                       @                                                              @                      �?      @                                                      O@      @      A@               @               @      d@     @\@      �?      @      @      Y@      C@              �?              @              "@      �?      @                              �?      =@      ?@      �?              �?      <@      .@              �?              �?              "@      �?      @                              �?      6@      3@                      �?      5@      *@              �?              �?                                                                      @      (@      �?                      @       @                                             �J@      @      ;@               @              @     ``@     �T@              @      @      R@      7@                              @              I@      @      ;@               @              @      ]@     @T@              @      @     �P@      7@                              @              @                                              @      .@      �?                      �?      @                                                     @W@      @      F@      @      @       @      &@     ``@     @[@       @      @      7@     �Y@     �T@              &@      @      (@      @      J@       @      3@       @      �?       @      $@     �T@      E@      �?       @       @      M@      M@               @              @              A@      �?      1@       @               @      @      R@      =@      �?       @      @      G@      C@                                              2@              @       @               @      �?     �I@      3@      �?       @      @      ;@      ;@                                              0@      �?      $@                              @      5@      $@                              3@      &@                                              2@      �?       @              �?              @      $@      *@                      �?      (@      4@               @              @              "@               @                              @      @      "@                              @      3@               @              @              "@      �?                      �?              @      @      @                      �?      @      �?                                             �D@      @      9@      @      @              �?     �H@     �P@      �?      @      .@      F@      8@              "@      @      "@      @      (@      �?      0@              @                      $@      8@      �?                       @      "@                       @       @              @              @                                      @       @                              @                                                      @      �?      $@              @                      @      6@      �?                      @      "@                       @       @              =@      @      "@      @       @              �?     �C@     �E@              @      .@      B@      .@              "@      @      @      @      1@       @      @      @       @              �?     �B@      C@              �?      ,@      A@      ,@              "@      @      @      @      (@      �?       @                                       @      @               @      �?       @      �?                                      �?     @d@     �P@      e@      A@     �K@      6@      J@     �^@     �i@      A@     �M@     �U@     @o@     @m@      (@     �C@     �G@     @R@     �B@     �S@      C@      Z@      5@     �C@      0@      >@      >@     @P@      0@     �A@     �K@      Y@     �Z@      @      :@      @@      B@      ;@     �R@      A@      W@      2@      =@      $@      5@      >@     �N@      $@      <@     �F@     �X@      Z@       @      6@      8@      ?@      3@      I@      6@     �F@      @      .@              ,@      7@      <@      @      4@      .@     �J@      J@              2@       @      7@      $@     �C@      ,@     �@@      @      (@              @      ,@      2@      @      &@      (@      :@      @@              $@      @      1@      @      .@      �?      2@      @      @              @       @      "@              @      @      @      2@              @       @      @      @      8@      *@      .@      �?      "@              �?      (@      "@      @      @      @      6@      ,@              @      @      &@       @      &@       @      (@       @      @              "@      "@      $@              "@      @      ;@      4@               @      �?      @      @      @      @      @              �?               @       @       @               @       @       @       @              �?              @              @       @      @       @       @              @      �?       @              @      �?      3@      (@              @      �?      @      @      8@      (@     �G@      (@      ,@      $@      @      @     �@@      @       @      >@     �F@      J@       @      @      0@       @      "@      @       @      (@              @              �?      @      .@      �?      @      @      9@      @              �?      @      @      @      �?              @              �?                              @                      �?      @                                       @       @      @       @      "@               @              �?      @      (@      �?      @      @      3@      @              �?      @      @       @      3@      $@     �A@      (@      &@      $@      @      �?      2@      @      @      :@      4@     �G@       @      @      *@       @      @      2@      @      8@       @      &@      @              �?      0@       @      �?      7@      (@      ?@       @              &@       @      @      �?      @      &@      @              @      @               @      @      @      @       @      0@              @       @              �?      @      @      (@      @      $@      @      "@              @      @      @      $@       @       @      @      @       @      @       @              @      �?      �?               @      @                       @      �?      @                               @              @                      @      �?      �?              �?                               @      �?      @                               @              @                                                      �?      @                                       @                                              �?              @              &@       @      $@      @       @              @      @      @      @       @       @      @       @       @      �?       @      @                              �?      �?      �?              @      @      @      @       @      �?      �?       @       @      �?      @      @                              �?      �?      �?                       @      �?               @      �?      �?      �?       @              �?                                                                      @      �?      @      @                              �?              �?      @      �?              &@       @      "@      @      �?              �?      �?       @      �?              �?      @              @              �?                      @               @      �?                                              �?              �?                                      �?      �?              @       @      @       @      �?              �?      �?       @                              @              @                      U@      <@     @P@      *@      0@      @      6@      W@     `a@      2@      8@      ?@     �b@      `@      @      *@      .@     �B@      $@     �C@      "@      4@      @      "@              @     �P@     �S@      @      (@      $@      N@      N@              "@       @      "@      @      (@      @      @              �?                      ,@      C@      @      @      @      8@      9@              @                              $@      @      @              �?                      @      9@      @      @      @      4@      7@                                              @      @       @              �?                       @      *@      �?              @      0@      ,@                                              @      �?      @                                      @      (@       @      @              @      "@                                               @      �?      �?                                       @      *@                      �?      @       @              @                              �?              �?                                      @      �?                      �?                              @                              �?      �?                                              @      (@                              @       @                                              ;@      @      ,@      @       @              @     �J@     �D@      @       @      @      B@     �A@              @       @      "@      @      @      �?      &@      �?      @                      "@      @               @              "@      (@              �?                              @      �?      @               @                      "@       @               @              @      $@              �?                                              @      �?      @                              @                              @       @                                              4@      @      @      @      @              @      F@      A@      @      @      @      ;@      7@              @       @      "@      @      @              �?                              @      @@      4@              �?       @      $@      ,@              �?       @      @      @      0@      @       @      @      @                      (@      ,@      @      @      @      1@      "@              @               @      �?     �F@      3@     �F@      "@      @      @      3@      9@      N@      (@      (@      5@     �V@      Q@      @      @      *@      <@      @      D@      *@     �F@      @      @      @      ,@      6@     �G@      $@      (@      4@     �S@     �G@      @      @      (@      9@       @      <@      &@      :@      @      @      @      (@      3@     �F@      @      (@      &@     �P@      B@      @      @      @      1@              ;@      @      7@      @      @      @      $@      ,@     �B@      @      &@      &@     �H@      B@      �?      @      @      0@              �?      @      @                               @      @       @              �?              1@               @                      �?              (@       @      3@       @                       @      @       @      @              "@      (@      &@              �?       @       @       @       @              $@       @                      �?              �?      �?              @      (@      @              �?      @      @              @       @      "@                              �?      @      �?       @              @              @                      @      @       @      @      @               @      @      �?      @      @      *@       @              �?      (@      5@       @              �?      @      @      @       @               @      @              @      @      (@                              (@      5@      �?              �?      @      @      @                       @      �?              �?       @      @                              @      (@                               @      @      �?       @                       @              @      �?      @                              "@      "@      �?              �?      �?                      @                              �?                      �?       @              �?                      �?                                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJRFhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKyhnh4h7K ��h9��R�(KKy��hu�Bx         >                    �?*[�ކ�?�	           ��@                          �2@-�=�G��?o           ��@                            @��ŵp��?F           ��@                           �?]��*���?�            �x@                          �1@��K����?s            �h@                            �?����b��?P            �`@������������������������       ��(�	��?            �C@������������������������       ���C��?6            �W@	       
                    @     P�?#             P@������������������������       ���g���?             K@������������������������       ����(\��?             $@                           @B���?|            �h@                          �0@^�v�T��?@            �X@������������������������       ��θ�?
             *@������������������������       ��������?6            @U@                            �?@$,�o��?<            �X@������������������������       �:e��5��?             ?@������������������������       ��8g�;��?+            �P@                          �1@����u�?W            `a@                           �?M��w���?5            �U@                           @���{���?            �@@������������������������       �:/����?             ,@������������������������       ��W�3��?	             3@                           @z-�-�?$            �J@������������������������       ���[r��?             5@������������������������       �     ��?             @@                           @�)���?"            �J@                           @lv�"��?             E@������������������������       �hE#߼�?             >@������������������������       �r�q��?             (@������������������������       ���!pc�?             &@        /                    @Ŷ���I�?)           L�@!       (                    �?L�d;]��?           h�@"       %                    �?'��%��?M           ��@#       $                   �;@�s<x{�?^            �b@������������������������       �RcB�%U�?Q            @_@������������������������       ��]�`��?             :@&       '                     @�q�qM�?�             x@������������������������       �y`����?�            �j@������������������������       �����/�?g            `e@)       ,                   �7@Ux�n�?�            `s@*       +                   �3@)ڵ�z��?            �g@������������������������       �<�i$���?            �E@������������������������       �N������?d            `b@-       .                    @�gE#��?K             ^@������������������������       �/�s��?'            �L@������������������������       ���Sm��?$            �O@0       7                    @Yֿ��,�?           `|@1       4                    @�kl����?L             _@2       3                    �?�r-�3�?;            @X@������������������������       �     ��?             @@������������������������       ��2;���?)            @P@5       6                     @������?             ;@������������������������       ���y4F�?             3@������������������������       �      �?              @8       ;                     @lEQ��=�?�            �t@9       :                     �?y�_0���?�            pp@������������������������       �.A6l�+�?0            �T@������������������������       �p�K��?m            �f@<       =                    @۝����?)            �P@������������������������       �B�?���?             G@������������������������       ��%7)��?             5@?       ^                   �9@ 7J�O��?8           D�@@       O                    �?�/{�?!           ��@A       H                   �5@�6����?�            �@B       E                    �?�K&��?
           @y@C       D                    �?6��P^C�?^             c@������������������������       ���T��?              M@������������������������       �j�g'�?>            �W@F       G                   �4@r�5A�r�?�            �o@������������������������       ��Q�,�?�            �h@������������������������       �R�X;�U�?&             K@I       L                    @�I)���?�            �p@J       K                   �8@pvh�L��?f            `e@������������������������       �snt+g�?N            ``@������������������������       ���Q��?             D@M       N                    �?�������?=            @X@������������������������       �4{d�?            �C@������������������������       ��#:9$A�?#             M@P       W                   �3@ܼ�<�?t           P�@Q       T                    @��B��3�?            z@R       S                    @���s�?�            �s@������������������������       �ܔ2���?�            Pp@������������������������       ��n�B�$�?"            �L@U       V                     �?�Wi�:�?B            �X@������������������������       ��Œ_,��?             >@������������������������       �.Lj����?-             Q@X       [                    �?SJS\(7�?`           P�@Y       Z                    @j�����?g             c@������������������������       �o(T���?            �@@������������������������       ����ƅ��?N            �]@\       ]                    @������?�             y@������������������������       �
"�[��??            �X@������������������������       �./�<���?�            �r@_       l                   �>@#`�v׮�?           �{@`       g                    @^jC�C]�?�            t@a       d                    @m�@ l�?�            �q@b       c                    @ԛ�XOn�?�             n@������������������������       ��nk���?�            @k@������������������������       ���JÝ�?             7@e       f                    @���<��?            �F@������������������������       �p_�Q�?             9@������������������������       ���Q��?             4@h       i                   �;@�����?            �A@������������������������       ��������?
             .@j       k                     �?�������?             4@������������������������       �      �?              @������������������������       ���8��8�?             (@m       r                    �?(p��xh�?K            �]@n       q                     @     ��?(             P@o       p                     �?:m���?             >@������������������������       ��������?             4@������������������������       �
ףp=
�?             $@������������������������       �N�]��?             A@s       v                    @������?#            �K@t       u                    @l�l��?             >@������������������������       �ZZZZZZ�?             1@������������������������       ��T�6|��?
             *@w       x                    @F%u��?             9@������������������������       �ƵHPS!�?             *@������������������������       �      �?             (@�t�bh�h4h7K ��h9��R�(KKyKK��h��B�G       `{@      S@     Pt@      D@      R@     �@@     @S@     �@     �@     �Q@     @U@     `b@     ��@     z@      .@     �Q@     �G@      \@     �O@     �i@      4@      _@      @      7@       @      7@     �v@     �u@      0@      E@     �E@     @s@     �f@      @     �@@      8@     �A@      9@     �F@      @      >@                               @     �h@     �^@       @      �?      (@     �R@      @@                              @              >@      @      (@                               @      e@     �V@              �?      (@      I@      7@                              �?              1@      @      @                                     @Y@      B@              �?      @      5@      $@                                              $@      @      @                                     �Q@      2@              �?      @      2@      @                                              @              @                                      .@       @              �?       @       @       @                                              @      @       @                                     �K@      $@                      �?      0@      @                                              @                                                      ?@      2@                              @      @                                              @                                                      >@      (@                              @      @                                               @                                                      �?      @                                      �?                                              *@      �?      @                               @     �P@      K@                      "@      =@      *@                              �?              @      �?      @                              �?      9@      B@                      @      &@      $@                              �?                                                                      @      $@                                                                                      @      �?      @                              �?      6@      :@                      @      &@      $@                              �?              $@              @                              �?      E@      2@                      @      2@      @                                              �?                                                      *@      (@                              @                                                      "@              @                              �?      =@      @                      @      *@      @                                              .@              2@                                      ?@     �@@       @                      9@      "@                              @              (@              @                                      8@      9@       @                      1@       @                                              @              �?                                      $@      .@      �?                       @                                                      @                                                      �?      @      �?                      �?                                                                      �?                                      "@       @                              �?                                                       @              @                                      ,@      $@      �?                      .@       @                                              �?                                                      @       @                              (@                                                      @              @                                       @       @      �?                      @       @                                              @              ,@                                      @       @                               @      @                              @              @              ,@                                      @       @                              @      @                              @              @              @                                      @       @                              @      @                              @                              "@                                       @                                              �?                                                                                                       @      @                              �?                                       @             �c@      0@     �W@      @      7@       @      5@     �d@     �k@      ,@     �D@      ?@      m@     �b@      @     �@@      8@      <@      9@     �\@      (@     �O@      @      6@       @      5@     �P@     @a@      $@      4@      ;@     �a@     @[@      @      6@      5@      4@      5@     @Q@      @      H@       @      2@       @      1@      B@      Q@       @      2@      2@     @V@      M@      @      4@      4@      .@      4@      :@              0@                               @      @      :@              @             �A@      *@      �?      "@      �?      @      @      .@              .@                               @      @      4@              @              A@      &@      �?      @      �?      @      @      &@              �?                                              @                              �?       @              @                             �E@      @      @@       @      2@       @      .@      >@      E@       @      .@      2@      K@     �F@       @      &@      3@       @      ,@      @@      @      3@              @              (@      5@      2@       @      &@       @      @@      8@              "@      @      @      @      &@      �?      *@       @      (@       @      @      "@      8@              @      0@      6@      5@       @       @      (@       @      @     �F@      @      .@      @      @              @      >@     �Q@       @       @      "@     �J@     �I@               @      �?      @      �?      ?@      @      @              �?               @      4@     �I@      @              @     �C@      6@                      �?      @              @                                                       @      "@                      @      (@      @                              �?              :@      @      @              �?               @      (@      E@      @              @      ;@      1@                      �?       @              ,@      @      $@      @      @               @      $@      3@       @       @      @      ,@      =@               @               @      �?      @              @      @      �?                      @      (@      �?              @      &@      @               @              �?              @      @      @               @               @      @      @      �?       @              @      8@                              �?      �?     �F@      @      ?@              �?                     @Y@     @U@      @      5@      @     �V@     �D@              &@      @       @      @      @              4@              �?                      D@      *@      �?      @      �?      =@      @              �?       @       @              @              3@              �?                      3@      (@      �?      @      �?      <@      @              �?       @       @               @              @                                       @      @              �?      �?      *@                                                      @              0@              �?                      &@       @      �?       @              .@      @              �?       @       @               @              �?                                      5@      �?                              �?      �?                                                                                                      0@      �?                              �?      �?                                               @              �?                                      @                                                                                              C@      @      &@                                     �N@      R@      @      2@      @      O@     �B@              $@      �?      @      @      >@      �?       @                                     �J@     �P@      �?      .@      @     �G@      :@              @      �?      @      @      @               @                                      "@      9@      �?      @      �?      0@      .@              @              �?              8@      �?      @                                      F@     �D@              (@       @      ?@      &@              �?      �?       @      @       @      @      @                                       @      @       @      @              .@      &@              @              @               @       @       @                                      @      @      �?      @              @      "@              �?               @                      �?      �?                                      �?              �?                      $@       @              @              �?             @m@      L@      i@      A@     �H@      9@      K@     `j@     �p@      K@     �E@      Z@     �t@     `m@      (@     �B@      7@     @S@      C@      j@     �D@      c@      8@      :@      *@      D@     �i@      n@      9@      @@     �P@      r@     �e@              5@      (@      I@      1@     �U@      3@      U@      @      1@      $@      1@     �K@     �R@      *@      2@      A@     �Y@      V@               @      @      7@      "@     �M@      &@      I@      @      "@      �?      *@     �B@     �L@      @       @      4@      P@      B@              @      @      2@      @      :@      @      "@               @      �?       @      2@      =@              @      @      7@      @              @       @      @      @       @                              �?               @       @      ,@               @      @      "@      �?              @       @       @              2@      @      "@              @      �?              $@      .@               @              ,@      @                              @      @     �@@      @     �D@      @      �?              &@      3@      <@      @      @      ,@     �D@      >@               @      �?      (@       @      :@      @      >@      @      �?              @      ,@      7@       @      @      &@     �C@      8@              �?              $@       @      @      @      &@                              @      @      @      �?              @       @      @              �?      �?       @              <@       @      A@      @       @      "@      @      2@      1@      $@      $@      ,@      C@      J@              @      @      @       @      6@      @      3@       @      @      "@       @      .@      1@      @      @      @      8@      <@                       @      @              .@      �?      ,@       @      @      @       @      *@      &@      @      @      @      1@      <@                       @       @              @      @      @               @      @               @      @       @      �?              @                                       @              @      @      .@       @      �?               @      @              @      @      @      ,@      8@              @       @      �?       @      @              @                              �?      @              @      @       @      &@      @              �?                       @       @      @      "@       @      �?              �?                       @      @      @      @      5@               @       @      �?             �^@      6@     @Q@      1@      "@      @      7@      c@     �d@      (@      ,@     �@@     �g@     �U@              *@      @      ;@       @      G@      @      ?@       @       @              @     @Y@     @T@       @      @      0@     �P@      A@               @      @      @       @     �B@      @      :@      @      �?              @     @V@     �G@       @      @       @      J@      :@               @       @      @       @      B@      @      8@       @      �?              @      R@      E@      �?      @      @      E@      4@              �?      �?      @              �?       @       @      @                              1@      @      �?      �?      @      $@      @              �?      �?      �?       @      "@              @       @      �?               @      (@      A@                       @      .@       @                      �?      �?              @                                                      @      .@                       @      �?                              �?      �?              @              @       @      �?               @      @      3@                      @      ,@       @                                              S@      1@      C@      "@      @      @      2@     �I@     @U@      $@      $@      1@     @^@     �J@              &@       @      4@      @      2@      @      @      @      �?      @      @      ;@      =@       @              @      3@      8@              @               @      @      @      �?       @                      @      �?              "@                      �?      @      @                              �?              (@      @      @      @      �?              @      ;@      4@       @               @      ,@      4@              @              �?      @      M@      &@     �@@      @      @              ,@      8@      L@       @      $@      ,@     �Y@      =@               @       @      2@      @      &@      �?       @       @                      "@      @      6@       @      @       @      2@      $@                               @      �?     �G@      $@      9@      @      @              @      4@      A@      @      @      (@      U@      3@               @       @      0@       @      9@      .@      H@      $@      7@      (@      ,@      @      8@      =@      &@     �B@     �D@      N@      (@      0@      &@      ;@      5@      7@      $@     �@@      @      3@      @      $@      @      1@      3@      @      0@      B@     �K@      @      (@      "@      7@      ,@      4@      $@      ?@      @      3@      @      "@       @      .@      2@      @      .@     �A@     �E@      @      "@      @      6@      &@      .@       @      :@      @      2@      @       @       @      *@      $@      @      .@      :@      C@      @      @      @      4@      &@      ,@       @      5@      @      0@      @      @       @      (@      $@      @      *@      9@      @@      @      @      @      3@      &@      �?              @               @              @              �?                       @      �?      @                              �?              @       @      @              �?              �?               @       @      @              "@      @               @               @                       @      @                                               @      @      @               @      @                                              @                              �?              �?                      �?                      @      �?               @               @              @               @      �?                      �?      �?       @      �?              �?      �?      (@              @      @      �?      @                       @                              �?      �?       @                      �?              @              @                              @                      �?                                              �?                      �?      @                      @      �?      @                                                                                                              @                      @              �?      @                      �?                                              �?                      �?      @                              �?       @       @      @      .@      @      @      @      @      �?      @      $@      @      5@      @      @      @      @       @      @      @      �?              @      @      @      @      �?              @       @      @      ,@                      @      @       @      �?      @                      �?       @      @      �?      �?              �?              �?      &@                              @      �?      �?       @                      �?      �?              �?      �?                              �?       @                              @              �?       @                              �?      @                              �?                      @                                      �?                      �?              @       @               @                       @       @      @      @                      @              �?              @      �?      @      "@      �?              @      @      �?      @       @              @      @      @                              @                      @       @      �?              �?              �?       @      @              @      @      @                              �?                               @      �?                              �?              @              @      @       @                                                      @                              �?                       @                      �?      �?       @                              �?              �?              @                       @      @               @      @              @              �?                               @              �?              �?                       @                       @      @                              �?                               @                              @                              @                                      @                                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJo�#%hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKyhnh4h7K ��h9��R�(KKy��hu�Bx         <                    �?�"널�?�	           ��@       !                    �?�D���?            ��@                           @��:�l�?x           x�@                           �?=�n����?�            �p@                            �?��)z��?P            �`@                          �1@��f�W�?2            �U@������������������������       ���'s�	�?	             1@������������������������       �&e<g��?)            �Q@	       
                    �?��8����?             H@������������������������       ���d�7��?             A@������������������������       ��X�C�?             ,@                           �?{Wr�E�?[            �`@                          �7@�]^m>��?<             W@������������������������       ��۫�$a�?)            �N@������������������������       ��>U��p�?             ?@                            @9��8���?             E@������������������������       ���)x9�?             <@������������������������       �^N��)x�?             ,@                           �?%t�û�?�             t@                          �8@�nY<�?S            @`@                          �5@��:�ե�??            �X@������������������������       ��噮��?)            �O@������������������������       ������H�?             B@                          �<@5yy8,�?             ?@������������������������       �fP*L��?             6@������������������������       ������H�?             "@                            @�������?z             h@                            �?I�$I�$�?I             \@������������������������       �/�����?:            �V@������������������������       ��ܤ��?             5@                           �1@�p=
���?1             T@������������������������       �VUUUUU�?             "@������������������������       ���=��?+            �Q@"       /                   �3@�W�kH�?�           T�@#       *                    @�z*U��?�            �q@$       '                    �?�2c��?�             l@%       &                   �1@���g�y�?/            �R@������������������������       �     ��?             @@������������������������       �+#eV�?            �E@(       )                    @F�g!���?[            �b@������������������������       ��M}�A��?L            @`@������������������������       ��z�G��?             4@+       .                    @P7�Z�?!            �L@,       -                    �?T�Y��?            �B@������������������������       ���ˠ�?             &@������������������������       �h��9J�?             :@������������������������       ��p=
ף�?	             4@0       7                    �?��c5�n�?�           ؇@1       4                   �4@�n}:���?�            `j@2       3                     �?)O���?             B@������������������������       �躍`3�?
             1@������������������������       �3�R�f�?
             3@5       6                     @�+m|���?s            �e@������������������������       ��J�w��?C            �Y@������������������������       ��͗(Cj�?0            @R@8       ;                   @A@��z9Kq�?V           @�@9       :                    �?C⹥XY�?I           ��@������������������������       �AM�h�'�?�             j@������������������������       �v�]Y~X�?�            t@������������������������       �@��Z��?             7@=       \                   �3@�S�l���?�           ʡ@>       M                   �1@Px���1�?K           ��@?       F                   �0@�����?           0{@@       C                    @ �qa�?]            `c@A       B                     �?�Y�H�7�?%             N@������������������������       �=[y��?             A@������������������������       �B�����?             :@D       E                    �?F%^�4�?8            �W@������������������������       �R���Q�?             D@������������������������       �*L�9��?            �K@G       J                     @y�Y�n~�?�            �q@H       I                     �?�jR��?�            �k@������������������������       ���Q����?k             e@������������������������       �~�	�[�?"            �J@K       L                    @o� 6 �?$            �M@������������������������       �~�Q���?             C@������������������������       ���i��i�?             5@N       U                    @��=���?=           �@O       R                    @��1v�j�?�            �v@P       Q                    @]+Yt��?�            �p@������������������������       �Iϙ D�?�            @j@������������������������       �>�>��?(             N@S       T                     @��v�@�?=            �W@������������������������       �fffff��?6             T@������������������������       �$߼�x�?             .@V       Y                     �?,U�&��?S             b@W       X                    �?]W���V�?1            �U@������������������������       ��4_�g�?             6@������������������������       �     ��?$             P@Z       [                   �2@`-�����?"            �M@������������������������       ��zv��?             6@������������������������       ����Z��?            �B@]       j                    �?X,QO�m�?J           Д@^       e                    @     ��?            x@_       b                    �?j\��54�?�            `l@`       a                   �6@b�[��y�?L            �\@������������������������       ���k
~�?)            �N@������������������������       �@�9S˅�?#             K@c       d                   �:@�X���?M             \@������������������������       ���`�i��??            �V@������������������������       �ܶm۶m�?             5@f       i                   �:@��g�a�?h            �c@g       h                   �6@�����?]            �a@������������������������       ����|���?<             V@������������������������       �GKv��x�?!            �J@������������������������       �     ��?             0@k       r                   �7@�"}���?I           ��@l       o                     �?t6���h�?F           ��@m       n                    @D�3�0
�?�            @s@������������������������       �N�zv�?(            �P@������������������������       �-x�mV��?�            @n@p       q                    @S�m׈��?�            �k@������������������������       ��&5D�?2             Q@������������������������       �r��o.��?R            `c@s       v                     @@\{��*�?           z@t       u                    @9sQFV#�?�            �t@������������������������       ��a�a�?1             U@������������������������       �7���Y��?�            `o@w       x                    �?0f�[
�?/            �T@������������������������       �
ףp=
�?             4@������������������������       �B�9(���?!             O@�t�bh�h4h7K ��h9��R�(KKyKK��h��B�G       @|@     �T@     pu@     �D@     @T@      ;@     �Q@     �@     ��@      M@      T@     @f@     `�@     @{@      $@     �R@      C@     ``@      I@     @j@     �A@      h@      4@      K@      2@      A@     �[@     @f@      =@     �I@      V@     �n@      g@      @      D@      9@     �Q@     �E@     @W@       @     �O@              5@               @      B@     �V@       @      ,@     �B@      Z@     �L@              &@       @      3@      ,@     �A@      @      B@               @               @      0@      H@      @      @      ,@      M@      ;@              @       @      @       @      2@      �?      7@                              �?      @     �@@      �?      @      @      >@       @              @                      �?      &@              *@                              �?      @      <@      �?      @      �?      .@       @              �?                      �?       @              "@                                      @       @                                      �?                                              "@              @                              �?      �?      :@      �?      @      �?      .@      @              �?                      �?      @      �?      $@                                      @      @                      @      .@                      @                              @      �?      @                                      �?      @                      @      @                       @                                              @                                       @                                       @                      �?                              1@      @      *@               @              �?      "@      .@       @      @      "@      <@      3@              �?       @      @      �?      *@      �?      @               @              �?      @      &@       @      @      @      &@      1@              �?       @       @      �?      $@      �?      @              �?              �?      @      $@      �?       @      @       @      @              �?      �?              �?      @              �?              @                              �?      �?      �?              @      &@                      �?       @              @       @      @                                      @      @                       @      1@       @                              �?              �?       @      @                                      �?      �?                       @      *@       @                                              @              �?                                       @      @                              @                                      �?              M@      @      ;@              *@              @      4@      E@      @       @      7@      G@      >@              @      @      0@      (@      5@              @              @              �?      (@      9@      �?      @      "@      3@      ,@               @      �?      @      @      2@              @              @                      "@      8@      �?      @      "@       @      (@                      �?      @       @      (@              @              @                       @      &@      �?      �?       @      @      @                               @              @                                                      �?      *@              @      �?      �?      @                      �?      �?       @      @              @                              �?      @      �?                              &@       @               @              �?      @      �?              �?                              �?      @      �?                              "@      �?               @              �?       @       @               @                                                                               @      �?                                       @     �B@      @      4@              "@              @       @      1@      @      @      ,@      ;@      0@              @      @      (@      @      (@      @      (@              @              @      @      (@      @      @      *@      2@      @              @      @      @      @      &@      @       @              @              @      @      (@      �?      �?       @      2@       @              @       @      @      @      �?              @                              �?      �?               @       @      @               @                      �?      �?      �?      9@      �?       @              @                      @      @      �?      �?      �?      "@      (@                       @      @      �?      @                                                      �?                                              �?                              @              5@      �?       @              @                      @      @      �?      �?      �?      "@      &@                       @      @      �?     @]@      ;@     @`@      4@     �@@      2@      :@     �R@      V@      5@     �B@     �I@     �a@     �_@      @      =@      1@     �I@      =@      =@      @      <@      @      @                     �G@      B@      @      @      @      P@      ;@              �?      �?      3@      @      9@      @      9@      @      @                      9@      @@       @      @      @      M@      2@              �?      �?      .@      @      @      @      @                                      2@      .@                              7@      @                              @      �?      @                                                      *@      @                              &@                                                              @      @                                      @      &@                              (@      @                              @      �?      5@       @      6@      @      @                      @      1@       @      @      @     �A@      .@              �?      �?      $@      @      4@       @      5@      @      @                      @      .@       @      @       @      >@      $@                              "@      @      �?              �?                                               @              �?       @      @      @              �?      �?      �?              @              @                                      6@      @      @              �?      @      "@                              @              @               @                                      2@      @                      �?      @       @                              �?              �?              �?                                      @       @                              �?                                                       @              �?                                      (@       @                      �?      @       @                              �?              �?              �?                                      @              @                              @                              @              V@      6@     �Y@      1@      >@      2@      :@      <@      J@      .@     �@@      G@     �S@      Y@      @      <@      0@      @@      9@      G@      @      1@      @      $@      @      @      ,@      ,@       @       @      &@      :@      ;@      �?       @      @      *@      �?      $@                              �?                      $@      �?                      @      �?      @                              @              @                                                       @                              @              @                              @              @                              �?                       @      �?                       @      �?      �?                                              B@      @      1@      @      "@      @      @      @      *@       @       @      @      9@      6@      �?       @      @      $@      �?      =@      @      $@       @      @              @      @      "@       @              @      @      ,@              �?      �?       @              @      @      @      @      @      @              �?      @               @      �?      2@       @      �?      �?      @       @      �?      E@      .@     @U@      &@      4@      ,@      7@      ,@      C@      *@      ?@     �A@     �J@     @R@      @      :@      &@      3@      8@      E@      .@      U@      "@      4@      ,@      7@      ,@      B@      *@      =@      =@     �J@     @R@       @      :@      &@      3@      1@      1@      @      ?@      @      @      @      (@       @      1@              (@      @      7@      @@              @      @       @      (@      9@      &@     �J@      @      0@      $@      &@      @      3@      *@      1@      6@      >@     �D@       @      4@      @      &@      @                      �?       @                                       @               @      @                      @                              @     @n@     �G@     �b@      5@      ;@      "@      B@     �x@     `|@      =@      =@     �V@     Pw@     �o@      @     �A@      *@     �N@      @     �X@      "@     �H@       @      �?              @     pp@     �m@      @      "@     �B@     @`@     @Q@               @      @      *@      �?      E@      @      (@              �?              �?     �a@      `@              @      1@     �N@      0@              �?              @              .@              @              �?                     �O@      G@              @       @      2@       @                               @              @               @              �?                      2@      8@              @               @      �?                                                               @                                      @      1@              @              @                                                      @                              �?                      *@      @                              �?      �?                                              (@              �?                                     �F@      6@                       @      $@      �?                               @              @                                                      7@       @                              @                                                      @              �?                                      6@      ,@                       @      @      �?                               @              ;@      @      "@                              �?     �S@     �T@                      .@     �E@      ,@              �?              @              7@      @      @                              �?     �P@     �P@                       @      >@      *@                              @              .@      @       @                              �?     �H@      L@                      @      6@       @                              @               @      �?       @                                      2@      $@                      �?       @      @                                              @              @                                      &@      0@                      @      *@      �?              �?              �?                              @                                       @      *@                      @      @                                                      @                                                      @      @                       @      @      �?              �?              �?             �L@      @     �B@       @                      @     �^@     �[@      @      @      4@     @Q@     �J@              @      @      @      �?      E@              <@                              �?      Z@     @R@       @      @      ,@     �K@      B@                       @      @      �?      @@              8@                              �?     �O@      N@       @      @       @      G@      :@                       @       @              <@              1@                                     �M@      E@       @      �?      @     �A@      2@                       @      �?              @              @                              �?      @      2@              @      @      &@       @                              �?              $@              @                                     �D@      *@                      @      "@      $@                              �?      �?      @              @                                     �D@      *@                               @       @                              �?              @                                                                                      @      �?       @                                      �?      .@      @      "@       @                      @      2@      C@      @       @      @      ,@      1@              @       @      @              *@      @      @       @                      �?      ,@      0@      @              @      @      "@              @       @       @               @                                              �?       @      $@                              @       @              �?                              &@      @      @       @                              (@      @      @              @      @      @              @       @       @               @              @                              @      @      6@               @       @      @       @               @              �?                              @                                      @       @                              @      @                              �?               @              �?                              @      �?      ,@               @       @      @      @               @                             �a@      C@     @Y@      3@      :@      "@      =@     �`@     �j@      8@      4@     �J@     `n@     �f@      @      ;@      "@      H@      @      H@      *@      3@      @      @      @      @      K@     @X@      @      @      (@      F@     �L@              "@       @      @              9@      @      0@      �?      �?      @       @      2@     �P@      @      �?      &@      @@      >@              @       @      @              (@      @      "@                      �?       @      "@      C@      �?              @      1@      ,@              @              �?              @      �?       @                      �?       @      @      :@                      �?       @      @                              �?              @      @      @                                       @      (@      �?               @      "@       @              @                              *@       @      @      �?      �?       @              "@      <@       @      �?       @      .@      0@               @       @      @              "@       @      @              �?       @              "@      <@                      @      $@      ,@               @              �?              @                      �?                                               @      �?       @      @       @                       @       @              7@      @      @      @       @               @      B@      ?@      @      @      �?      (@      ;@              @              �?              7@              @      @       @               @      B@      ;@      @      @      �?      &@      7@              @              �?              2@              �?      @      �?                      1@      .@              �?      �?      "@      3@              @                              @               @              �?               @      3@      (@      @       @               @      @                              �?                      @                                                      @                              �?      @                                             �W@      9@     �T@      .@      7@      @      9@     @T@     �]@      2@      0@     �D@     �h@     �_@      @      2@      @     �E@      @      P@      $@     �A@      @      @              @      J@     @V@      @      @      6@     �a@     �L@       @      "@      @      .@      �?     �C@      @      :@      @      @              @      >@      O@      @      @      0@      M@      >@              "@      @       @      �?      $@      @      @      �?      @              �?      &@      �?       @               @      (@      &@               @      �?       @              =@      �?      6@       @      @              @      3@     �N@      �?      @      ,@      G@      3@              @       @      @      �?      9@      @      "@       @                      �?      6@      ;@       @       @      @      U@      ;@       @              �?      @              @              @       @                      �?      "@      "@              �?      @      2@      "@                      �?                      2@      @      @                                      *@      2@       @      �?      �?     �P@      2@       @                      @              ?@      .@     �G@      $@      0@      @      4@      =@      =@      *@      "@      3@     �L@     @Q@       @      "@      @      <@      @      <@      $@     �E@       @      (@      @      $@      :@      7@      *@       @      1@      I@      G@              @      @      8@      @      "@      �?      3@      @              �?              $@      @      @       @       @       @      @                      @      @              3@      "@      8@      @      (@      @      $@      0@      1@      @      @      "@      E@      E@              @              5@      @      @      @      @       @      @       @      $@      @      @              �?       @      @      7@       @      @              @      �?      �?      �?       @       @                              �?      @              �?              @       @              �?                               @      @       @              @       @      $@       @      @                       @      �?      5@       @       @              @      �?�t�bub�R     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�o�ChG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         8                    �?!	.)��?�	           ��@                           �?n(=s�$�?�           @�@                            �?�mD*��?l           0�@       	                    �?��t�'8�?d            `b@                           8@�:�Ń��?             E@                           �?d�ϙ�?             ;@������������������������       ���8��8�?             (@������������������������       ��������?             .@������������������������       �
ףp=
�?             .@
                          �7@�im��?E            @Z@                           @��ĳ���?(             N@������������������������       ��&5D�?
             1@������������������������       ��|S�ݮ�?            �E@                          �=@��ٯi\�?            �F@������������������������       �_������?            �A@������������������������       ��(\����?             $@                          �4@���y��?           0{@                           �?ڟ��+�?o            @f@                           @������?9            �V@������������������������       �_���D�?3            @T@������������������������       �ffffff�?             $@                            @�=C|F�?6            �U@������������������������       ��X�g�?             A@������������������������       �>α�
��?            �J@                           �?��e\���?�            p@                           @h�9��?:            �X@������������������������       ��n�MJ��?2             U@������������������������       ��'}�'}�?             .@                            �?�G��/�?_            �c@������������������������       �t|��?)            �Q@������������������������       �������?6            �U@        /                   �=@K���&*�?�           (�@!       (                   �3@�Y	l'��?U           @�@"       %                    @�ɲ���?�            Pq@#       $                   �1@
�J���?            @i@������������������������       �[�[��?1            �R@������������������������       ��3:�^��?N            �_@&       '                    �?���=��?/            �R@������������������������       ���i��i�?             5@������������������������       �� .E3�?!             K@)       ,                    �?��Sp��?�           ��@*       +                    �?����[�?�            �p@������������������������       �#8̺�8�?;             W@������������������������       ���6���?u            @f@-       .                   �8@dpt?�?�            Px@������������������������       ���t���?�            @o@������������������������       ���U�a�?T            `a@0       5                   �@@����%^�?>            �X@1       4                   @@@\���"�?&            �N@2       3                    �?Ukט��?            �F@������������������������       ��x�W�?             7@������������������������       ��#��Z=�?             6@������������������������       �      �?	             0@6       7                     �?������?            �B@������������������������       ��'}�'}�?
             .@������������������������       �h���eP�?             6@9       X                   �2@ZV�wC��?�           �@:       I                    �?��ZH���?�           `�@;       B                    @oa�+��?�            �q@<       ?                     @�7��W�?_            `b@=       >                     �?
���W�??            �X@������������������������       �~�Q���?             C@������������������������       �贁N��?#             N@@       A                    �?�V���?             �H@������������������������       �#����?             ;@������������������������       �fP*L��?             6@C       F                     �?������?J             a@D       E                    @�S�%
&�?/            @V@������������������������       ��֤����?            �H@������������������������       ��p=
ף�?             D@G       H                   �0@��8��)�?            �G@������������������������       �                     "@������������������������       �����U�?             C@J       Q                    @�ze�~�?           {@K       N                     �?�U����?�            `i@L       M                    @���,��?I            �[@������������������������       ��D��v�?8            �U@������������������������       ��(��0�?             9@O       P                    @?�)
;&�?8             W@������������������������       �����[��?             B@������������������������       �������?#             L@R       U                    �?Oa��[��?�            �l@S       T                    @      �?M             \@������������������������       ��q�q�?             8@������������������������       �n,�Ra��?>             V@V       W                    @��Ԃ���?E            �]@������������������������       ��������?!             N@������������������������       �z��sk��?$             M@Y       d                    �?=^}�t�?�           ��@Z       a                   �=@q���R��?<           �@[       ^                   �6@ 
Z.ҫ�?0            @\       ]                     @َ=�ͤ�?�            �r@������������������������       �n�m�<w�?�            �n@������������������������       �~h����?#             L@_       `                     �?2Tv���?|            `h@������������������������       �Gس����?D            @X@������������������������       ��������?8            �X@b       c                   �>@|�l�]�?             1@������������������������       �9��8���?             @������������������������       �������?             &@e       l                    �?�^�]���?�           ��@f       i                   �8@x�Q�WF�?1           �}@g       h                     �?{v�X��?�             v@������������������������       �Y�(%LL�?�            �i@������������������������       ������?c            `b@j       k                     @��ڎ���?K            @^@������������������������       �b�|���?@            �Y@������������������������       ����Hx�?             2@m       p                    @���l>��?�           ��@n       o                   �3@�hz-���?$           0|@������������������������       ��	�O��?-            �Q@������������������������       ����y��?�            �w@q       r                    @�������?a             b@������������������������       ��]���?:            @T@������������������������       ���s{��?'            �O@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       0y@     �T@     Pu@      @@      O@      ;@     �V@     �@      �@      N@     @Y@      f@     �@     �}@      &@     �Q@     �K@     @_@     �F@      e@      A@     @e@      1@      C@      3@     �C@      _@     @h@      ?@     �N@     �Y@     �l@     �i@      @      E@      E@     �N@      @@      Q@      &@     �B@      �?      (@       @      (@     �O@     �T@      (@      ?@      >@     �Y@      L@              6@      "@      6@      "@      1@      @      $@      �?      @      �?      @       @      4@       @      @      @     �B@      &@              @       @      @      @      @              @              �?                      @      *@              @               @      @                      �?      �?              @              @                                      @      @                              @      @                              �?               @               @                                       @       @                              @      �?                                               @              �?                                       @      @                              �?      @                              �?                                              �?                              @              @              @                              �?                      *@      @      @      �?       @      �?      @      @      @       @      �?      @      =@      @              @      �?      @      @       @              @      �?      �?                       @      @                      @      :@      @                              �?      @      �?              @                                      �?       @                              $@                                                      @               @      �?      �?                      �?       @                      @      0@      @                              �?      @      @      @       @              �?      �?      @       @      @       @      �?      @      @      @              @      �?      @              @      @                      �?      �?               @       @              �?      @      @      @              @      �?      @                               @                              @              �?       @                                               @                             �I@      @      ;@              "@      �?      "@     �K@     �O@      $@      ;@      7@     @P@     �F@              .@      @      0@      @      >@              @              @              �?      A@      9@      @       @      (@      5@      2@              @      @      @      @      *@              @               @                      :@      1@      @      @      @      $@      @              @               @      �?      *@               @                                      :@      *@      @              @      $@      @              @               @      �?                      �?               @                              @              @                                                                      1@                              �?              �?       @       @      @      @      @      &@      .@              @      @       @       @      @                                              �?      @      @      �?              @      @       @               @                      �?      ,@                              �?                      @      @       @      @      �?       @      @               @      @       @      �?      5@      @      8@              @      �?       @      5@      C@      @      3@      &@      F@      ;@               @      @      (@       @      $@      @      "@              �?      �?      �?      "@      9@              @       @      1@      @              @               @               @      @      "@              �?      �?      �?      @      9@              @       @       @      @              @               @               @                                                      @                                      "@      �?                                              &@       @      .@              @              @      (@      *@      @      ,@      "@      ;@      4@              @      @      $@       @      @              @              @              @       @      @      �?      "@      @      1@      $@               @                      �?      @       @      (@              �?                      $@       @      @      @      @      $@      $@              �?      @      $@      �?     @Y@      7@     �`@      0@      :@      1@      ;@     �N@     �[@      3@      >@      R@      `@     �b@      @      4@     �@@     �C@      7@     �W@      6@     @_@      ,@      3@      $@      ;@     �N@     �[@      *@      6@     �L@     �_@     �a@      �?      .@      6@     �A@      2@      A@      @      :@      �?                      @      A@      G@              @      "@      G@      E@               @      @      2@      @      8@      @      6@      �?                      @      3@     �C@              @      @      C@      7@                      @      *@      �?      ,@      �?       @                              �?      *@      "@                       @      2@      @                      @      �?              $@       @      ,@      �?                      @      @      >@              @      @      4@      2@                              (@      �?      $@              @                                      .@      @                      @       @      3@               @              @       @      @              �?                                      @      @                      �?       @      �?               @                              @              @                                      $@      @                       @      @      2@                              @       @      N@      3@     �X@      *@      3@      $@      7@      ;@     @P@      *@      0@      H@     @T@     @Y@      �?      *@      3@      1@      .@      ?@      @     �I@              @      �?      @      $@     �A@              @      1@     �D@     �@@      �?      @      &@      @      @      ,@      @      7@               @              @      �?      @               @      @      2@      &@      �?                       @      �?      1@      @      <@              @      �?      @      "@      =@              @      (@      7@      6@              @      &@       @      @      =@      (@      H@      *@      *@      "@      0@      1@      >@      *@      $@      ?@      D@      Q@              "@       @      *@      $@      7@      @      B@      @      @      @      @      ,@      6@      @      "@      1@      6@      H@              @       @      "@      @      @      @      (@      $@      @      @      $@      @       @      @      �?      ,@      2@      4@              @              @      @      @      �?       @       @      @      @                              @       @      .@      �?      @      @      @      &@      @      @      @      �?      @       @      @      @                              @      @      @      �?      @              @       @      @              @      �?      @       @      @      @                              @      @      @      �?       @              @       @      @              @      �?                       @                                              �?      @      �?       @              @              @               @              @       @      �?      @                              @       @                                      �?       @                                      �?                      �?                                      @                      @              �?      @                                      @              @                                      @      �?      &@                      @              @              @                       @                                                      @              "@                                                      �?                       @              @                                              �?       @                      @              @              @     @m@     �H@     `e@      .@      8@       @     �I@     z@      z@      =@      D@     �R@     pw@     �p@      @      <@      *@      P@      *@     �P@      @     �F@              @              $@     `k@     �d@       @      @      ,@     �Z@     �M@              @      �?      @      �?      3@              4@                              @      \@      O@      �?       @      @      A@      4@              @              �?              *@              0@                              @     �I@      >@      �?       @      @      7@      @              �?                              @               @                              @     �D@      :@      �?       @              *@       @              �?                              @                                                      "@      *@               @               @       @              �?                              @               @                              @      @@      *@      �?                      @                                                      @              ,@                                      $@      @                      @      $@       @                                              @              @                                      @      @                              @       @                                               @              @                                      @      �?                      @      @                                                      @              @                               @     �N@      @@                      �?      &@      0@               @              �?              @              �?                                      C@      8@                      �?       @       @               @              �?                              �?                                      ;@      *@                              @      @                                              @                                                      &@      &@                      �?      @      @               @              �?                              @                               @      7@       @                              @       @                                                                                                      "@                                                                                                              @                               @      ,@       @                              @       @                                              H@      @      9@              @              @     �Z@      Z@      �?      @      $@     @R@     �C@              �?      �?      @      �?      *@      @      2@                              �?     �L@      I@              @              E@      .@                                              $@      @      @                              �?      ?@      :@              @              9@      "@                                              @      �?      @                                      >@      5@              @              2@      @                                              @       @                                      �?      �?      @                              @       @                                              @              .@                                      :@      8@              �?              1@      @                                              �?              @                                      "@      @              �?              *@                                                       @              $@                                      1@      1@                              @      @                                             �A@       @      @              @              @      I@      K@      �?      �?      $@      ?@      8@              �?      �?      @      �?      9@              �?                              �?      ?@      ?@      �?              @      &@       @                                              @                                                       @      .@      �?                       @      �?                                              6@              �?                              �?      =@      0@                      @      "@      @                                              $@       @      @              @              @      3@      7@              �?      @      4@      0@              �?      �?      @      �?      @       @      @              @              @      @      $@              �?              0@      (@                              �?              @              �?                                      0@      *@                      @      @      @              �?      �?      @      �?     �d@      F@     �_@      .@      5@       @     �D@     �h@     �o@      ;@     �@@      N@     �p@     `j@      @      8@      (@      M@      (@      F@      0@     �A@       @      @      @      @     �O@      [@      @      @      4@     �V@     �U@              "@      @      "@       @     �E@      .@     �A@       @      @      @      @     �O@      [@      @      @      0@     �T@      U@              "@       @      "@       @      6@      �?      3@       @              @       @      F@      R@              �?      "@      N@     �M@              �?      �?      @      �?      3@      �?      2@                       @       @     �C@     @P@              �?       @     �E@     �F@                      �?              �?      @              �?       @              �?              @      @                      �?      1@      ,@              �?              @              5@      ,@      0@              @       @      @      3@      B@      @      @      @      6@      9@               @      �?      @      �?      "@              *@              @              @      *@      6@      @       @       @      (@      &@              @                              (@      ,@      @              @       @      �?      @      ,@               @      @      $@      ,@              @      �?      @      �?      �?      �?                                                                              @       @       @                      �?                      �?      �?                                                                              �?       @      �?                                                                                                                                      @      @      �?                      �?                     �^@      <@     �V@      *@      .@      @     �A@     �`@      b@      7@      <@      D@     @f@     @_@      @      .@      "@     �H@      $@      M@      *@     �@@      @      @              "@     �S@     �R@      @      0@       @      S@     �K@              "@      @      1@      @      F@      @      6@      @       @              @      Q@      Q@      @       @      @      L@     �B@              @      @      ,@             �@@      �?      "@       @       @              @      @@     �H@              @      @      >@      8@              @      @      @              &@       @      *@      @                      @      B@      3@      @      @       @      :@      *@              �?               @              ,@      $@      &@              @               @      $@      @       @       @      @      4@      2@              @              @      @      $@      $@      $@              @               @      $@      @       @      @      @      3@      1@              @              @              @              �?                                              @              �?              �?      �?               @                      @     @P@      .@      M@       @      "@      @      :@     �L@     @Q@      0@      (@      @@     �Y@     �Q@      @      @      @      @@      @      J@      (@      E@      @      @      �?      0@     �I@     �L@      .@       @      5@     �T@     �D@      @      @      �?      ;@      @      1@              @              @                      ,@      .@      @       @      �?      "@                                                     �A@      (@      B@      @      @      �?      0@     �B@      E@      &@      @      4@     @R@     �D@      @      @      �?      ;@      @      *@      @      0@      @       @       @      $@      @      (@      �?      @      &@      4@      =@      �?              @      @      �?      @      �?      *@      @      �?       @      @       @      @      �?              @      .@      &@      �?              @      @      �?      @       @      @              �?              @      @      @              @      @      @      2@                      �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�AiJhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKqhnh4h7K ��h9��R�(KKq��hu�B�         6                   �5@������?�	           ��@                            @�s>pi��?N           �@                           �?���&�?�           Ę@                           @�˰��?           @{@                           �?;�[�D��?	           �z@                          �3@��J���?r            �f@������������������������       ��!k\��?J            �[@������������������������       �����L��?(            �Q@	       
                   �2@3�l��N�?�            �n@������������������������       ��\L�k��??            @[@������������������������       ��'s�	U�?X             a@������������������������       ���"e���?             "@                          �2@%�&7ǧ�?�           ��@                            �?g��xqu�?_           Ё@                           @�}����?�            0y@������������������������       ����Zv�?�            Ps@������������������������       ��/"93��?7            �W@                           @��1H��?e            �d@������������������������       ��盢���?V            �a@������������������������       ���@����?             9@                           @���0�y�?j           �@                           @RDBF�E�?P            �`@������������������������       �d��E��?'             Q@������������������������       �h���eP�?)            �P@                           �?�k����?           �{@������������������������       ���� !��?x            `e@������������������������       ��G���?�             q@       )                    @u$K�;�?u           �@       $                    �?`�ĪW �?*            }@       !                    �?�H�y�?�            `t@                            �?������?G             \@������������������������       ����S�r�?             E@������������������������       ��.��D��?*            �Q@"       #                   �1@�n�Z�9�?�            �j@������������������������       �&K:�m��?!             K@������������������������       �H�z��?g             d@%       (                   �4@�������?[            @a@&       '                    @�#�]��?O            @^@������������������������       ��7�A�?8             V@������������������������       �,j�J��?            �@@������������������������       �|�l�]�?             1@*       /                    @�p��V�?K            @\@+       ,                    �?U��6���?             A@������������������������       �����>4�?	             ,@-       .                   �2@q=
ףp�?             4@������������������������       �r�q��?
             (@������������������������       �      �?              @0       3                    �?p��D׀�?2            �S@1       2                    @4{d�?            �C@������������������������       �c}h���?             <@������������������������       �}��7�?             &@4       5                   �2@\���(\�?             D@������������������������       ����Դ�?             3@������������������������       �����X�?             5@7       T                    �?[�KG?�?D           \�@8       E                    �?�`zf�P�?)           ��@9       >                   �6@���t-��?�            `r@:       =                     @c�/��b�?&             N@;       <                    @���[���?            �F@������������������������       �
ףp=
�?             4@������������������������       ���H�}�?
             9@������������������������       �[�[��?             .@?       B                    �?�.�{B��?�            @m@@       A                   �;@��I��I�?'             N@������������������������       ��� =�	�?             ?@������������������������       �c��gS~�?             =@C       D                    �?li#�,��?s            �e@������������������������       �,�ѳ��?&             Q@������������������������       ��R�:��?M            �Z@F       M                    �?|_�h�v�?i           X�@G       J                   �9@-"}�o��?\            `d@H       I                     @������?+            @R@������������������������       ����Hx�?             B@������������������������       �*e��}`�?            �B@K       L                     �?�P�a�r�?1            �V@������������������������       ���N8��?             E@������������������������       ��q�1�?             H@N       Q                    �?��t��f�?           �z@O       P                     @������?             K@������������������������       ��!pc��?             6@������������������������       �     ��?             @@R       S                    @���Ӕw�?�             w@������������������������       ���?��!�?n            @e@������������������������       �n4��@��?�             i@U       b                    �?g#�u��?           0�@V       ]                     @)C/Ap�?�            @n@W       Z                     �?�Sd�/;�?�             h@X       Y                    �?�Ft��?T            @`@������������������������       �K&:~��?0             S@������������������������       �ߍL�t��?$             K@[       \                    �?���5��?,            �O@������������������������       �+f��ӫ�?             5@������������������������       �*�s���?             E@^       a                   �:@|xV��f�?            �H@_       `                    @F��'s��?             A@������������������������       ��z6�>�?             9@������������������������       �~X�<��?             "@������������������������       ��A��S�?             .@c       j                    @zF���	�?�           ��@d       g                     @4���,��?M            �^@e       f                    @r�q�?>             X@������������������������       � *4>HR�?#            �I@������������������������       �ǿ��S��?            �F@h       i                   �7@���d�?             ;@������������������������       ��(\����?             $@������������������������       �躍`3�?	             1@k       n                    @:e%kn��?3           �@l       m                    @�$�F��?�            �v@������������������������       �q[� sA�?�            �r@������������������������       �bE'���?,            �Q@o       p                     @xA�@��?V            `a@������������������������       �p՘�}�?A            @Z@������������������������       �����.�?             A@�t�bh�h4h7K ��h9��R�(KKqKK��h��BC       P~@     �S@      t@     �A@     �P@      A@     �T@      �@     h�@     �P@     �T@     `c@     (�@     �z@      (@      Q@      K@      a@     �L@     �r@      6@      a@      $@      $@      @      B@     0{@     �x@      :@      ;@     �R@     x@     �f@              7@      *@     @P@      5@     �l@      0@     �U@      @      @              7@      w@     s@      .@      2@     �I@     �p@     ``@              *@      @      =@      0@      S@      @      >@      @      @              &@     �O@     �Q@      @      "@      3@     @S@      C@              @              (@      *@     �R@      @      >@      @       @              &@      O@     �Q@      @      "@      3@     @S@      A@              @              (@      (@     �D@       @      @                              @      ;@      :@      �?      @      @     �E@      (@              @                       @      ;@       @      @                                      6@      5@      �?      @      @      1@       @                                              ,@               @                              @      @      @               @      �?      :@      @              @                       @     �@@       @      7@      @       @              @     �A@      F@       @      @      ,@      A@      6@                              (@      $@      &@              @               @              �?      :@      4@       @              &@      6@      @                              @      �?      6@       @      0@      @                      @      "@      8@              @      @      (@      3@                              "@      "@       @                              �?                      �?                                              @                                      �?      c@      (@     �L@      @      @              (@     s@     `m@      (@      "@      @@     `g@     @W@               @      @      1@      @     @Q@      @      0@                              @     �g@      _@      @              $@      V@      F@              @      @      @      �?     �N@      @      $@                              @     �Z@     �Y@      @              "@      N@      =@              @      @      @      �?     �A@      �?      @                              @     �V@      T@       @              @      K@      8@              �?       @       @      �?      :@      @      @                                      .@      6@      �?              @      @      @              @       @      @               @      �?      @                                      U@      6@       @              �?      <@      .@                                              @      �?      @                                     �S@      0@       @              �?      5@      *@                                              @                                                      @      @                              @       @                                              U@      @     �D@      @      @              "@     �\@     �[@      @      "@      6@     �X@     �H@              @      @      (@       @      2@              @              �?              @      6@      C@                      @      ;@      *@                              @              �?               @                              �?      *@      5@                      @      4@      @                                              1@              @              �?               @      "@      1@                              @      @                              @             �P@      @     �A@      @       @              @     @W@     @R@      @      "@      3@      R@      B@              @      @      "@       @      3@      �?      (@                              @     �@@      @@               @      @      D@      2@              �?       @               @     �G@      @      7@      @       @               @      N@     �D@      @      @      ,@      @@      2@              @      �?      "@             �P@      @      I@      @      @      @      *@     �P@     @V@      &@      "@      7@     @^@      J@              $@      @      B@      @      L@      @      A@       @      @      @      @      D@     @Q@      $@      @      7@     �Z@      H@              "@      @      ?@      @      B@      @      =@              �?      �?      @      9@     �G@      "@      @      0@     �O@      C@              "@      @      <@      @      ,@      �?      @                                      $@      0@      @      @      @      6@       @              @      @      @      �?      @              �?                                      @      &@      �?                      "@       @               @              @              @      �?      @                                      @      @      @      @      @      *@      @              @      @      @      �?      6@      @      6@              �?      �?      @      .@      ?@       @      @      &@     �D@      >@              @              6@       @      "@       @      @                                      (@       @              �?              (@      @                                              *@      @      0@              �?      �?      @      @      7@       @       @      &@      =@      :@              @              6@       @      4@              @       @      @      @      �?      .@      6@      �?      �?      @     �E@      $@                              @      �?      4@              @       @      @      @              .@      6@      �?      �?      @     �A@      @                              �?      �?      0@              @      �?       @      @              *@      *@                       @      ;@      @                                      �?      @                      �?      �?                       @      "@      �?      �?      @       @      �?                              �?                              �?                              �?                                      �?       @      @                               @              &@              0@      �?                      "@      ;@      4@      �?       @              .@      @              �?              @      �?      �?              &@                                      "@      @              �?              @                                       @                              @                                      @      @              �?                                                                      �?              @                                      @      @                              @                                       @                              @                                      @      �?                               @                                                      �?              �?                                               @                               @                                       @              $@              @      �?                      "@      2@      ,@      �?      �?              &@      @              �?              @      �?      @              @                              @      "@      @      �?      �?              @       @                               @               @              @                                      "@      @              �?              @       @                              �?              �?                                              @                      �?                      @                                      �?              @               @      �?                      @      "@      @                              @       @              �?              �?      �?       @              �?                              @      @      �?                               @                      �?              �?      �?      @              �?      �?                      �?       @      @                              @       @                                             �g@     �L@     �f@      9@     �L@      =@     �G@     @\@     `h@      D@      L@     @T@     �l@     �n@      (@     �F@     �D@      R@      B@     @U@      8@     �Z@      .@      C@      4@      ;@      6@     �V@      ;@     �E@     �B@      Y@     �`@       @      7@      8@     �@@      9@      <@      @      A@       @      .@      @      @      $@     �E@      "@      .@      @      L@     �C@              @      @      @       @      @              @       @                              @      @      �?                      8@      @              �?      �?      �?      @      @              @       @                               @      @                              5@      @              �?      �?                      @               @       @                              �?      @                              @      @                      �?                                      �?                                      �?      @                              2@      �?              �?                                              @                                       @      �?      �?                      @      �?                              �?      @      7@      @      <@              .@      @      @      @      B@       @      .@      @      @@      A@              @      @      @      @      @      �?       @                              @       @      1@               @      �?      "@      @               @      �?               @      @      �?                                               @       @              �?      �?      @       @               @      �?               @      �?               @                              @              "@              @               @      @                                              2@       @      :@              .@      @      @      @      3@       @      @      @      7@      <@              �?      @      @      @      $@              @              �?       @              �?      *@      @      @      �?       @      .@              �?       @                       @       @      4@              ,@      �?      @      @      @      @      @      @      .@      *@                       @      @      @     �L@      5@      R@      *@      7@      1@      4@      (@      H@      2@      <@      ?@      F@     �W@       @      3@      2@      ;@      1@      A@      @      4@      @      @       @      @      @      .@      @      �?       @      .@      3@       @      @      @      "@       @       @       @       @      @      @      @       @      @      @       @                       @      .@              @      @                      @      �?      @                               @      @       @       @                      @      &@                                              @      �?      �?      @      @      @                      �?                              @      @              @      @                      :@       @      (@      �?      @       @      �?              (@      @      �?       @      @      @       @      �?              "@       @      (@      �?      �?      �?       @              �?              @      @                              @       @                      "@              ,@      �?      &@              �?       @                      @              �?       @      @                      �?                       @      7@      1@      J@      @      1@      "@      1@       @     �@@      *@      ;@      =@      =@     �R@      @      ,@      .@      2@      .@              �?      @              @      @               @      @      @       @               @      .@      �?      �?              �?      @              �?      @               @                                      �?       @              @      @              �?              �?                                              �?      @               @      @      @                      @      (@      �?                              @      7@      0@      G@      @      ,@      @      1@      @      >@      "@      9@      =@      5@      N@      @      *@      .@      1@      (@      .@      @      :@      @       @      �?      @      @      &@      @      @      0@      @      =@               @      @      "@      @       @      $@      4@      @      @      @      (@              3@      @      2@      *@      0@      ?@      @      @      "@       @      @      Z@     �@@     @S@      $@      3@      "@      4@     �V@      Z@      *@      *@      F@      `@      \@      @      6@      1@     �C@      &@     �@@      (@      *@              @      @       @      :@     �F@      @      @      &@      =@     �A@              &@       @      @       @      >@      @      *@              �?      @      �?      9@     �B@      @      @      @      9@      6@              @              @       @      3@              &@              �?                      3@      =@      @      @      @      1@      2@               @              @              &@              @                                      ,@      :@      �?       @       @      &@      @                                               @              @              �?                      @      @      @      �?       @      @      *@               @              @              &@      @       @                      @      �?      @       @      �?              @       @      @              @              @       @      @      �?                                              �?      @                       @      @      �?                                               @      @       @                      @      �?      @       @      �?              �?      �?      @              @              @       @      @      @                       @              �?      �?       @                      @      @      *@              @       @                      @      @                       @              �?      �?      @                       @      @      *@                       @                      �?       @                       @                      �?      @                       @       @      (@                                               @      �?                                      �?              �?                              �?      �?                       @                               @                                                      @                       @      �?                      @                             �Q@      5@      P@      $@      0@      @      2@     @P@     �M@       @      $@     �@@     �X@     @S@      @      &@      .@     �@@      "@      *@      @      4@      @                              3@      &@       @               @      (@      &@       @              &@      @              &@      @      4@       @                              1@      @       @              @      "@      @                      &@      @              $@       @       @      �?                              @      �?       @              @      @      @                      @      @              �?      �?      (@      �?                              (@      @                              @      @                       @                       @      �?              @                               @      @                      @      @      @       @                                       @                                                       @      �?                              @       @                                                      �?              @                                      @                      @               @       @                                      M@      1@      F@      @      0@      @      2@      G@      H@      @      $@      9@     �U@     �P@       @      &@      @      <@      "@      E@      ,@      8@       @      ,@      �?      0@     �D@     �F@      @      @      (@     �P@      I@               @      �?      (@      @      ?@      ,@      5@               @      �?      @      =@      C@      @      @      &@      P@     �E@              @              "@      @      &@              @       @      @              "@      (@      @               @      �?      @      @              @      �?      @              0@      @      4@      @       @      @       @      @      @      �?      @      *@      4@      0@       @      @      @      0@       @      .@              1@      @      �?               @      @      @      �?      @      &@      ,@      "@              �?      @      .@       @      �?      @      @              �?      @               @                               @      @      @       @       @              �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�p�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKkhnh4h7K ��h9��R�(KKk��hu�Bh         :                     @Fa}iۡ�?�	           ��@                          �2@w�~��O�?�           ��@                           @�r���?�           ��@                           �?�\;��?�            �r@                          �0@b���y��?x            �f@                            �?�h70�?             ?@������������������������       ��ˠT�?             &@������������������������       ��G�z��?             4@	       
                    �?�k-j�?f            �b@������������������������       �p�`��3�?)            �O@������������������������       ��K���?=            �U@                            �?Ng�fk�?I            @]@                          �0@��m���?A             Z@������������������������       ��1�^���?             A@������������������������       �|�ۨ�?,            �Q@������������������������       ��]�`��?             *@                          �0@@��wԘ�?'           @@                           @���/Z�??            @Z@������������������������       �      �?             (@                           @��y� �?8            @W@������������������������       �f�ft��?+            �Q@������������������������       ��nkK�?             7@                          �1@\�ʰj7�?�            �x@                           @8l#!���?r            �i@������������������������       ����a_�?U             c@������������������������       �#�o�h�?            �J@                           @�,����?v            �g@������������������������       �(��`���?S            �`@������������������������       �H���?#            �L@       +                    �?���Ǝ��?�           t�@       &                    �?��.�X�?�           ��@        #                    �?xu,����?�             p@!       "                   �:@�;�����?7            @T@������������������������       ���X��?'             L@������������������������       ���+e��?             9@$       %                    �?���o���?x             f@������������������������       �����K�?4             R@������������������������       �������?D            @Z@'       *                    @6hW���?"           �}@(       )                     �?���D���?           �|@������������������������       ��O�q��?�            �w@������������������������       �����|�?0            �S@������������������������       �g\�5�?             *@,       3                   �8@��7_�?           �@-       0                    @f{��<��?J           ȍ@.       /                    @�"j�!�?�            �l@������������������������       ��*S�`��?t            @i@������������������������       ��(ݾ�z�?             :@1       2                    �?Gl��?�           ��@������������������������       ��%����?�            �m@������������������������       �Sz�b��?4           �~@4       7                   �;@�Lw���?�            �t@5       6                    @��S�y8�?f            �e@������������������������       ���U &�?1            �U@������������������������       �7�A�0�?5             V@8       9                    �?��+��0�?^             c@������������������������       ��-��1��?$             O@������������������������       �E��l��?:            �V@;       P                    �?c����?�           8�@<       G                    �?��3TU�?�           H�@=       B                   �7@x��?r            �g@>       ?                   �1@*��-�?S            `a@������������������������       �lv�"��?             5@@       A                    �?�,�$�?D            �]@������������������������       ���WV��?             J@������������������������       ���+j�?'            �P@C       D                    �?�A`��"�?             I@������������������������       ��.k���?             1@E       F                    @���!pc�?            �@@������������������������       �ףp=
��?             4@������������������������       �����W�?             *@H       O                    @�f,�X�?;           �~@I       L                    �?�ͫ�gU�?3            ~@J       K                    @��I!k��?~            `j@������������������������       ������?w            �h@������������������������       �؂-؂-�?             .@M       N                   �5@-*W�`�?�            �p@������������������������       ��H��J��?X            �`@������������������������       ���}����?]            �`@������������������������       �      �?             (@Q       ^                    �?��bi�?           Pz@R       W                    �?�l����?�            @g@S       T                   �1@�m۶m��?(             L@������������������������       �      �?
             0@U       V                   �3@>
ףp=�?             D@������������������������       �r�q��?
             (@������������������������       �Y�Cc�?             <@X       [                    @��O_[�?X            @`@Y       Z                   �1@x¹�T��?             E@������������������������       ��.�?��?             .@������������������������       ��P���?             ;@\       ]                   �1@�|���?<             V@������������������������       ���>4և�?	             ,@������������������������       �������?3            �R@_       d                   �1@B)�®�?�            `m@`       a                   �0@�������?             H@������������������������       �     ��?	             0@b       c                    @     ��?             @@������������������������       �L�9���?             6@������������������������       �
ףp=
�?             $@e       h                    @/t��?            `g@f       g                    �?Z�S�O�?+            @P@������������������������       ��ѳ�w�?             1@������������������������       �     @�?             H@i       j                    @�յ?�?T            �^@������������������������       ��:�Ń��?              E@������������������������       �333333�?4             T@�t�bh�h4h7K ��h9��R�(KKkKK��h��B�?       �y@      X@     �s@     �D@     �V@      7@      T@     ؁@     ��@      M@     �T@     @h@     h�@     �z@      $@     �P@      L@     �\@      P@     �r@      N@      k@      5@     �J@      @     �H@     0~@     �~@      D@     �P@     �`@     �z@     q@      @      G@      @@      S@      D@     �U@      @      6@              �?               @     `o@     �h@      @      @      :@     @^@     �K@              @      @       @      @      D@              (@              �?              @      P@     �S@       @      @      1@      G@      5@                      �?      @      @      7@              @              �?              @     �A@     �D@               @      .@     �A@      (@                              @       @       @                                                      *@      $@                              @      �?                                              �?                                                      @      @                              @      �?                                              �?                                                      $@      @                               @                                                      5@              @              �?              @      6@      ?@               @      .@      >@      &@                              @       @      ,@               @                                      *@      &@              �?      @      ,@      @                                              @              @              �?              @      "@      4@              �?      &@      0@      @                              @       @      1@              @                                      =@      C@       @       @       @      &@      "@                      �?              �?      .@              �?                                      8@     �B@       @       @       @      &@       @                      �?              �?      �?                                                      @      4@                              @                                                      ,@              �?                                      2@      1@       @       @       @      @       @                      �?              �?       @              @                                      @      �?                                      �?                                              G@      @      $@                              @     `g@     @]@      �?              "@     �R@      A@              @       @      @              .@                                                      M@      .@                      �?      ,@      �?                              �?                                                                      @      @                                                                                      .@                                                      J@      "@                      �?      ,@      �?                              �?              @                                                      E@      @                      �?      &@      �?                              �?               @                                                      $@       @                              @                                                      ?@      @      $@                              @      `@     �Y@      �?               @     �N@     �@@              @       @       @              0@       @      @                               @     @Q@     @Q@                      @      :@      "@                              �?              @              @                               @     �L@      M@                      @      .@      @                                              "@       @      �?                                      (@      &@                      @      &@      @                              �?              .@      @      @                              @      N@     �@@      �?               @     �A@      8@              @       @      �?              @              @                              �?      J@      5@                      �?      >@      3@                                              "@      @       @                               @       @      (@      �?              �?      @      @              @       @      �?             @j@      K@     @h@      5@      J@      @     �D@      m@     pr@     �B@      O@     �Z@     @s@     @k@      @     �D@      =@      Q@     �B@      S@      7@      U@      @      7@      �?      :@     �H@     @R@      (@     �D@     �G@     �W@     �T@      �?      5@      ,@     �@@      <@     �C@      @      >@      �?      @              (@      <@      ;@      �?      *@       @     �F@      8@                      @      @      $@      0@      @      (@      �?      �?              �?      @      .@              @              ,@      @                              @               @              (@      �?      �?                      @       @              @              *@      �?                              @               @      @                                      �?              @               @              �?       @                                              7@       @      2@              @              &@      6@      (@      �?       @       @      ?@      5@                      @      @      $@      &@               @                              @      .@      @      �?      @       @      1@      @                              �?       @      (@       @      0@              @              @      @      @              @      @      ,@      .@                      @       @       @     �B@      1@      K@      @      2@      �?      ,@      5@      G@      &@      <@     �C@     �H@      M@      �?      5@      &@      ;@      2@      B@      1@     �J@      @      2@      �?      ,@      5@      F@      &@      ;@     �C@     �H@     �I@      �?      4@      &@      ;@      2@      >@      1@     �D@      @      0@      �?      ,@      1@     �B@       @      :@      9@     �D@      D@      �?      4@      @      7@      0@      @              (@               @                      @      @      @      �?      ,@       @      &@                      @      @       @      �?              �?                                               @              �?                      @              �?                             �`@      ?@     �[@      1@      =@       @      .@     �f@     �k@      9@      5@      N@     �j@      a@      @      4@      .@     �A@      "@     �Z@      5@     @R@      ,@      1@      �?      "@      b@     `h@      @      0@      F@     �c@      Y@      �?      .@      @      5@      @      3@      @      4@      @      @      �?      �?      6@      L@      �?      �?      "@     �G@      A@                              @              .@      @      0@      @      �?      �?      �?      6@     �K@      �?              "@      B@      A@                              @              @              @              @                              �?              �?              &@                                                      V@      1@     �J@      &@      &@               @     �^@     `a@      @      .@     �A@     �[@     �P@      �?      .@      @      1@      @      6@      @      &@                              �?      F@      Q@       @      @       @      C@      ;@              �?       @      �?       @     �P@      *@      E@      &@      &@              @     �S@     �Q@      @      "@      ;@      R@     �C@      �?      ,@      @      0@      @      ;@      $@     �B@      @      (@      �?      @     �C@      ;@      3@      @      0@     �L@      B@       @      @      $@      ,@       @      5@      @      4@              @      �?       @      ;@      ,@      @      @      "@      C@      *@              @              @              .@      �?      "@              �?      �?       @      2@      @      �?      �?      @      &@      @              @              @              @      @      &@              @                      "@      @      @      @      @      ;@      "@                              �?              @      @      1@      @      @              @      (@      *@      ,@              @      3@      7@       @              $@       @       @      @       @      @      �?      @              @      (@      @       @              @       @       @                                      �?       @      @      &@       @       @              �?               @      (@               @      &@      .@       @              $@       @      �?     �\@      B@     @Y@      4@      C@      4@      ?@      V@     �`@      2@      0@     �N@      d@     �b@      @      5@      8@      C@      8@     �Q@      :@     @Q@      ,@      ?@      2@      .@      A@     �P@      .@      *@     �E@      U@      Y@      @      *@      5@      6@      4@      4@      @      3@              @              @      .@      .@      "@      @      *@      8@      >@              �?      @      &@      @      ,@       @      ,@              @              @      ,@      *@       @      @      "@      4@      ,@              �?      @      $@      �?      @              @                                      @              �?              �?      �?                                      @               @       @      $@              @              @      $@      *@      @      @       @      3@      ,@              �?      @      @      �?      @              @                                      "@      @      @              @      &@       @                              @              @       @      @              @              @      �?      @      @      @      @       @      @              �?      @       @      �?      @      @      @                              �?      �?       @      �?      �?      @      @      0@                       @      �?      @      �?      �?       @                              �?               @              �?      �?      @      @                                       @      @       @      @                                      �?              �?              @      �?      *@                       @      �?      �?               @      @                                      �?              �?                      �?      "@                       @      �?              @                                                                                      @              @                                      �?     �I@      5@      I@      ,@      8@      2@      $@      3@      J@      @      @      >@      N@     �Q@      @      (@      0@      &@      0@      I@      4@      I@      *@      8@      1@      $@      3@      J@      @      @      :@      L@     �Q@      @      (@      0@      &@      0@      :@      @      0@       @      $@               @      &@      :@              @      &@     �B@      <@              @      &@      @      @      :@      @      $@       @      @               @      &@      8@              @      $@     �B@      <@               @      $@      @      @                      @              @                               @                      �?                               @      �?                      8@      ,@      A@      &@      ,@      1@       @       @      :@      @      @      .@      3@      E@      @       @      @      @      &@      7@      *@      .@      @      @      �?               @      ,@      @       @      @      (@      4@              �?      @      @              �?      �?      3@      @      "@      0@       @              (@       @       @       @      @      6@      @      @       @      �?      &@      �?      �?              �?              �?                                              @      @                                                      F@      $@      @@      @      @       @      0@      K@     �P@      @      @      2@      S@     �I@      �?       @      @      0@      @      3@       @      $@      �?      �?      �?      @      >@     �@@      @      @      @      A@      <@              @       @      @       @      @               @              �?      �?              @      ,@                      �?      *@      ,@              �?              �?                               @                                       @       @                              @                                                      @                              �?      �?               @      @                      �?      "@      ,@              �?              �?               @                                                      �?                                      @      @                                               @                              �?      �?              �?      @                      �?      @      $@              �?              �?              .@       @       @      �?                      @      :@      3@      @      @      @      5@      ,@               @       @       @       @      @               @      �?                              @      "@      �?      �?      @      ,@       @                                                                                                              @      �?                      "@                                                      @               @      �?                              @      @              �?      @      @       @                                              $@       @      @                              @      6@      $@       @       @      @      @      (@               @       @       @       @      @              @                                       @      �?                                      �?                                              @       @       @                              @      4@      "@       @       @      @      @      &@               @       @       @       @      9@       @      6@      @      @      �?      (@      8@      A@                      &@      E@      7@      �?      @      �?      *@       @      @              @                                      ,@      0@                      @      @                       @               @                              �?                                       @      @                                                                                      @               @                                      @      "@                      @      @                       @               @              @               @                                      @      @                      @       @                                       @                                                                       @      @                               @                       @                              6@       @      3@      @      @      �?      (@      $@      2@                      @      C@      7@      �?      @      �?      &@       @      @       @      @       @      �?              @      @      $@                       @      $@      (@               @              @              �?      �?      �?                                              @                      �?      �?      @                              @               @      �?      @       @      �?              @      @      @                      �?      "@      "@               @              @              3@      @      .@      @      @      �?      @      @       @                      @      <@      &@      �?      �?      �?      @       @      @       @      (@      @                      �?              @                       @      $@       @                              �?      �?      ,@      @      @              @      �?      @      @      @                      @      2@      "@      �?      �?      �?      @      �?�t�bub��	     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJYb)hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKqhnh4h7K ��h9��R�(KKq��hu�B�         6                    �?�#b���?�	           ��@                           �?���o0�?           �@                          �8@FN\y��?z           ��@                           @5�q�Y�?           `{@                           �?�+?��?�            �q@                          �6@[=;n,�?S            �`@������������������������       ���)x9��?H             \@������������������������       �333333�?             4@	       
                    �?"V��HD�?c             c@������������������������       �
ףp=
�?0             T@������������������������       �qm�UL�?3            @R@                            @Q}�֭h�?b             c@                            �?�{�~V�?:             U@������������������������       �     ��?             @@������������������������       ��h��9�?$             J@                          �2@��t{H�?(            @Q@������������������������       �8�Z$��?             :@������������������������       �#��,�?            �E@                          �?@��q�qj�?b            �c@                          �<@��6�?X            �a@                           @9��8���?;             X@������������������������       ��n�MJ��?             E@������������������������       ��c�_p��?"             K@                            �?3��'$��?            �F@������������������������       �j�V���?            �@@������������������������       ���8��8�?             (@������������������������       �ZZZZZZ�?
             1@       '                    �?��ls�D�?�           ��@                           �1@c��P2��?�            �q@                           �?Jf%�9��?            �B@������������������������       �$I�$I��?	             ,@������������������������       ����Q��?             7@!       $                   �3@���#���?�            �n@"       #                    �?L�9���?             F@������������������������       ���i��i�?             5@������������������������       ���JÝ�?             7@%       &                    �?��a��?�            @i@������������������������       �;N�F��?>            @W@������������������������       �	`��uW�?M            @[@(       /                   �5@�Q|�I�?�           ��@)       ,                   �3@���ӿ6�?�            Ps@*       +                     �?�6K@��?~             h@������������������������       �5���?%             J@������������������������       �;�Aξ��?Y            �a@-       .                    �?� B�~�?G             ]@������������������������       �j��i���?             E@������������������������       ��,b+���?,            �R@0       3                     @��P^Cy�?            z@1       2                    @�^�P�D�?�            �l@������������������������       ��j�Y�H�?"             N@������������������������       �O���3�?t            @e@4       5                   @A@��l�	j�?|            �g@������������������������       ���<4�?t            �e@������������������������       �n�����?             .@7       R                    @�"�3���?�           �@8       C                     �?&7�����?f           H�@9       <                   �0@��{��?}             j@:       ;                    @����<��?            �@@������������������������       �     ��?	             0@������������������������       �                     1@=       @                   �9@颋.�(�?m             f@>       ?                   �2@˱C;��?Z            �a@������������������������       ���؉���?             :@������������������������       ���p%]^�?F             ]@A       B                    �?�.k���?             A@������������������������       �hE#߼�?	             .@������������������������       �Ɓ�r�z�?
             3@D       K                   �6@r�yd}�?�            �w@E       H                   �3@��$� �?�             o@F       G                     @��f8K��?V            �`@������������������������       ��%���^�?,             R@������������������������       ��b�b�?*             O@I       J                   �4@}�3�)q�?C            �\@������������������������       ��q�1�?             H@������������������������       ���;���?)            �P@L       O                     �?{̭:���?P            �_@M       N                    �?�2�o�U�?&            �K@������������������������       �      �?             0@������������������������       �~T��@o�?            �C@P       Q                    �?����[��?*             R@������������������������       �-C��6�?             9@������������������������       �������?            �G@S       b                    �?�l;^t��?3           �@T       [                   �1@������?j           X�@U       X                    �?�z<�L�?`            `b@V       W                    @9��e���?;            �V@������������������������       �\���(\�?             D@������������������������       ���Ƽ���?             �I@Y       Z                    @����S��?%             L@������������������������       �*x9/��?             <@������������������������       �ܶm۶m�?             <@\       _                    @,mG8��?
           �{@]       ^                     @�c�_dE�?�            �q@������������������������       ��Kx��?�            �m@������������������������       �_|�!�?             G@`       a                    �?��d�)��?]            �c@������������������������       ��
�6�?/            �T@������������������������       ��
I���?.             S@c       j                    @{�&��?�           ��@d       g                    @D'K�҅�?�           �@e       f                    �?z�'���?'            }@������������������������       ���gג3�?�            `l@������������������������       �����G�?�            �m@h       i                    @ƫ�����?�            �p@������������������������       �JKA7���?�            �m@������������������������       �     ��?             @@k       n                   �5@*s9b��?�            �x@l       m                    @���Ƕ�?�             k@������������������������       ��E��Y��?$             O@������������������������       ��i+�v�?b            `c@o       p                    �?�������?s            �f@������������������������       �q�{%�?,            @P@������������������������       ��"sV�?G             ]@�t�bh�h4h7K ��h9��R�(KKqKK��h��BC        ~@      U@      t@     �D@     �T@      ;@     �U@     ��@     ��@     �Q@     �S@      e@     �@     �|@      .@      N@      G@     @`@      G@     @i@      F@     `d@      ,@     �K@      1@     �E@     �^@     �b@     �C@     �F@     �W@     @j@     �k@      $@      A@     �@@     �Q@      C@     �T@      *@     �E@              8@       @      &@      N@     �Q@      1@      .@     �A@     �W@     �Q@               @      (@      8@      *@     �Q@      @      <@              @      �?      @     �K@      N@      @      $@      ;@     �R@      J@              @       @      .@      $@      B@      @      .@              @              @      G@      E@       @      @      *@      L@      C@              @      @      @      @      3@              @                              �?      =@      4@               @      @      ;@      ,@               @      @              @      .@              @                              �?      :@      2@                      @      :@      ,@               @                      �?      @              �?                                      @       @               @              �?                              @              @      1@      @       @              @              @      1@      6@       @      @      $@      =@      8@              �?       @      @       @       @               @                               @      ,@      .@       @      @      @      ,@      @              �?       @      @      �?      "@      @      @              @               @      @      @                      @      .@      2@                                      �?      A@       @      *@              @      �?      �?      "@      2@      @      @      ,@      2@      ,@                      @      $@      @      3@      �?       @               @              �?       @      .@              @      "@      .@      @                               @              @      �?      �?                                      @       @              �?      @      $@      @                               @              .@              �?               @              �?      @      *@               @      @      @      @                                              .@      �?      &@               @      �?              �?      @      @      �?      @      @      @                      @       @      @      @              @                                              �?                                      @                              @      @      $@      �?      @               @      �?              �?       @      @      �?      @      @       @                      @      �?              (@       @      .@              1@      �?      @      @      &@      $@      @       @      5@      3@              @      @      "@      @      $@       @      ,@              *@      �?      @      @      &@      $@      �?      @      5@      3@               @      @      @      @      "@       @      @              "@      �?               @       @      "@      �?      �?      0@      0@               @      @      @      @      @                              @                              @      @                      $@      @              �?      @      @       @      @       @      @               @      �?               @      @      @      �?      �?      @      "@              �?              @      �?      �?      @      @              @              @      @      @      �?              @      @      @                      �?                              @      @              �?              @      @      @                      @       @       @                                              �?       @                      @                                      �?                      @      �?                      �?                       @              �?              @                                              @      �?                              @               @              ^@      ?@      ^@      ,@      ?@      .@      @@      O@      T@      6@      >@      N@     �\@     �b@      $@      :@      5@      G@      9@      G@      @      9@      @      .@       @      @      1@     �@@      @      @      *@      H@      ?@       @       @       @      ,@      @      @      �?                      @                       @      @                              &@      @                                      �?                                                              @      �?                              @       @                                              @      �?                      @                      �?       @                              @      @                                      �?     �E@      @      9@      @      (@       @      @      "@      >@      @      @      *@     �B@      8@       @       @       @      ,@      @      @      @      @                                       @      *@              @      �?      @       @                              @              �?      @      @                                      �?      @              �?              @                                       @               @              @                                      �?      @               @      �?      @       @                              �?              D@       @      2@      @      (@       @      @      @      1@      @              (@      >@      6@       @       @       @      &@      @      <@              @      �?       @               @      @      @                       @      4@      $@       @      �?              @              (@       @      *@      @      $@       @      �?      @      &@      @              @      $@      (@              �?       @      @      @     �R@      9@     �W@      $@      0@      *@      =@     �F@     �G@      0@      ;@     �G@     �P@     �]@       @      8@      *@      @@      4@     �J@      $@      D@      �?      �?              @      B@      ?@      �?      @      "@     �D@      I@              @      �?      $@       @      >@      @      .@      �?                       @      ?@      8@      �?      @      @      =@      =@              �?      �?       @      @      @       @       @                              �?      (@      @      �?      @               @      "@                              �?      @      ;@      @      *@      �?                      �?      3@      2@              �?      @      5@      4@              �?      �?      @       @      7@      @      9@              �?               @      @      @              @      @      (@      5@              @               @       @      *@              @                                      @      �?              �?       @      @      $@              �?                              $@      @      2@              �?               @       @      @               @      �?       @      &@              @               @       @      5@      .@     �K@      "@      .@      *@      9@      "@      0@      .@      4@      C@      :@     @Q@       @      2@      (@      6@      (@      .@      $@     �@@       @      @      @       @      @      @      &@      &@      4@      *@      C@              *@      "@      3@      @              @      @      �?      @              �?      @      �?      @      @      �?       @      .@              @      @      @              .@      @      ;@      �?      @      @      @      @      @       @      @      3@      &@      7@              @      @      ,@      @      @      @      6@      @      "@      $@      1@      @      $@      @      "@      2@      *@      ?@       @      @      @      @      @      @      @      6@      @      @      $@      ,@      @      $@      @       @      1@      *@      ?@              @      @      @      @                                       @              @                              �?      �?                       @                                     `q@      D@     �c@      ;@      <@      $@     �E@     �{@     Pz@      @@     �@@     �R@      w@     �m@      @      :@      *@      N@       @     @P@      .@     �C@      @      &@      @      &@      R@     �`@      "@      @      4@     �T@     �R@       @      @              6@      @      6@      @      $@      @      @      @      @      2@      Q@      @      @      $@      :@      *@              �?              &@      �?      �?                                                      @      8@                               @                                                      �?                                                      @      @                               @                                                                                                                      1@                                                                                      5@      @      $@      @      @      @      @      (@      F@      @      @      $@      8@      *@              �?              &@      �?      3@       @       @      @       @      @      @      &@     �E@      �?      @      @      7@       @              �?              @               @               @                                      @       @      �?              �?      @       @                                              &@       @      @      @       @      @      @      @     �D@              @       @      3@      @              �?              @               @      @       @              �?       @              �?      �?       @              @      �?      @                              @      �?       @      @                                              �?      �?                      @              @                               @                               @              �?       @                               @              @      �?       @                              @      �?     �E@      $@      =@      @       @      �?      @      K@     �P@      @      �?      $@     �L@      O@       @      @              &@       @      <@      @      .@              @              @      F@     �M@      �?      �?      @     �E@      B@                              @              2@      �?      @              @              @      =@      7@              �?       @      =@      2@                              @              @              �?              �?              @      :@      $@                              &@      &@                              @              (@      �?      @               @                      @      *@              �?       @      2@      @                                              $@       @      &@                               @      .@      B@      �?              @      ,@      2@                              �?              @                                              �?       @      2@                              @      &@                                              @       @      &@                              �?      @      2@      �?              @      $@      @                              �?              .@      @      ,@      @      @      �?       @      $@      @      @              @      ,@      :@       @      @              @       @      "@      �?      &@                      �?              @      @      @               @      @      *@              �?               @              @               @                                      �?      �?                              �?       @                                              @      �?      @                      �?              @       @      @               @       @      &@              �?               @              @      @      @      @      @               @      @      @      �?              �?      &@      *@       @      @              @       @      @      @              �?                                      �?                              @      @              �?               @              �?              @       @      @               @      @      @      �?              �?       @      @       @       @              @       @     �j@      9@      ^@      5@      1@      @      @@     @w@     �q@      7@      :@      K@     �q@     `d@      @      5@      *@      C@      @     �P@      @     �B@      @       @      @       @     �b@     @_@      @       @      $@     �T@      M@              @      @      @       @      (@      �?      @                                      S@     �@@                       @      *@      @                              �?              @      �?      @                                     �K@      2@                       @      @      �?                                              @      �?                                              3@      (@                      �?      @                                                      �?              @                                      B@      @                      �?       @      �?                                              @              �?                                      5@      .@                               @      @                              �?              @              �?                                      @      $@                              @      @                                              �?                                                      0@      @                              @                                      �?             �K@      @      @@      @       @      @       @      R@      W@      @       @       @     �Q@      K@              @      @      @       @      =@      @      6@      @      @      @      �?     �J@     @P@      @       @      @     �I@      9@                      @      �?      �?      7@      @      "@              �?      @              I@      P@      @       @      @     �C@      6@                      @      �?              @              *@      @       @              �?      @      �?                              (@      @                                      �?      :@      �?      $@              @              @      3@      ;@       @              @      3@      =@              @      @      @      �?      *@              @                                      (@      3@                              *@      2@                                              *@      �?      @              @              @      @       @       @              @      @      &@              @      @      @      �?     @b@      3@     �T@      1@      "@      �?      8@      l@     @d@      1@      2@      F@     @i@     @Z@      @      2@      @     �@@      @      W@      &@     �G@      $@      @              0@     �e@     �Z@      $@      *@      2@      a@     @P@      �?      @      @      4@      @     �Q@      @      <@      $@      @              ,@     @X@     �Q@      @      &@      *@     �R@     �C@              @       @      &@      @      B@              $@      �?                      &@     �J@      D@      @      @       @     �A@      6@                       @      @             �A@      @      2@      "@      @              @      F@      >@      @      @      &@      D@      1@              @              @      @      5@      @      3@                               @     �R@     �B@      @       @      @     �N@      :@      �?      �?       @      "@              5@      @      2@                                     �Q@      ?@      @       @      @      H@      5@      �?      �?       @      "@                              �?                               @      @      @                              *@      @                                              K@       @      B@      @      @      �?       @      J@     �K@      @      @      :@     �P@      D@       @      &@      @      *@             �A@      @      (@       @       @              @     �D@      D@      �?      �?      ,@      A@      *@              @              @              @      @      @               @                      @      ,@                      @      1@      @                              �?              ?@      �?      "@       @                      @      A@      :@      �?      �?      $@      1@      @              @              @              3@      @      8@      @       @      �?      @      &@      .@      @      @      (@      @@      ;@       @      @      @      @              @       @      @                                      @      (@      �?      @       @      &@      $@              @              @              (@       @      5@      @       @      �?      @      @      @      @              $@      5@      1@       @      �?      @      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ8)�LhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         @                    �?1gF�?�	           ��@       !                   �4@^��<�?
           d�@                           �?������?v           `�@                           �?��R�&�?�            Pp@                           @�j6��?P            �_@                           @xɃg\�?@             Z@������������������������       �t��O��?2            @T@������������������������       ���,d!�?             7@	       
                     �?�袋.��?             6@������������������������       ��z�G��?	             $@������������������������       �r�q��?             (@                            @�m���?R            �`@                           @     @�?(             P@������������������������       ��������?             8@������������������������       ��z�G��?             D@                           �?���T<�?*            �Q@������������������������       �      �?             8@������������������������       ��W+J���?            �G@                           @�`˛.4�?�            pt@                            @2$�?�            �n@                          �2@p��ю��?O            @^@������������������������       ��:8`�S�?+            @P@������������������������       �����>4�?$             L@                           �?
�2oD�?T            �_@������������������������       ��{��9��?            �A@������������������������       ��g��H��?<            �V@                           @�Q��k�?1             T@                           �?$�����?!            �J@������������������������       ��fG-B��?             5@������������������������       �     ��?             @@                            �?��F�� �?             ;@������������������������       �؂-؂-�?             .@������������������������       ��8��8��?	             (@"       1                    �?"�>�@��?�           4�@#       *                    @�Q0�?           �{@$       '                    �?�6��=�?�            �q@%       &                   �6@���߈�?X             c@������������������������       ���m(�9�?            �E@������������������������       �+1�o'��??            �[@(       )                   �6@�M�N��?R            �_@������������������������       ��LG�;6�?            �F@������������������������       �<�M��?5            �T@+       .                   �>@�,�V9��?h            �d@,       -                   �9@h/�����?[             b@������������������������       �튑DW�?A            @Z@������������������������       �ĒN0��?            �C@/       0                   �@@�7�A�?             6@������������������������       ��zv��?             &@������������������������       �b���i��?             &@2       9                    �?ġ���?�           x�@3       6                   �<@7���
�?�            �j@4       5                     @�弿���?s            �e@������������������������       �>
ףp=�?M             ^@������������������������       ����dIG�?&             K@7       8                     �?
ףp=
�?             D@������������������������       �P�|�@�?             1@������������������������       ��s-s��?             7@:       =                   �>@n�	ze}�?�            �w@;       <                     @�=q��N�?�            0u@������������������������       �o�}� �?v            �e@������������������������       �9N/o���?h            �d@>       ?                    @t��:��?             C@������������������������       �     @�?             0@������������������������       �J���#��?             6@A       `                     @����?�           �@B       Q                   �3@,��R��?�           ��@C       J                    @�T�����?�           X�@D       G                    @�]9V�?y           ��@E       F                    @J4��D�?%           p{@������������������������       ���XE���?�            `s@������������������������       ���q$�w�?R             `@H       I                    @������?T            �_@������������������������       ��KL���?.            �R@������������������������       ������?&            �J@K       N                   �0@����|6�?i            �f@L       M                    �?pƵHP�?             :@������������������������       ��>�>��?             .@������������������������       �Y�����?             &@O       P                    �?�����?[            `c@������������������������       ��y3�`�?            �I@������������������������       ��؉�؉�?<             Z@R       Y                    �?�m�B��?�           �@S       V                    @[��^�_�?E           �@T       U                   �6@���Q��?�             n@������������������������       ��}�g���?;            �X@������������������������       �*~*�sD�?Z            �a@W       X                    @gB� ݧ�?�            q@������������������������       ��`m:*G�?q            �e@������������������������       �ԝ�����??            @Y@Z       ]                    �?����?x            �@[       \                    �?Hy1���?|            `g@������������������������       �tz��y�?f            @b@������������������������       �
�c�"�?            �D@^       _                    @/"!�d��?�            �x@������������������������       ������?�            �s@������������������������       �ǁZ|� �?-            �R@a       d                   �0@}h��e�?"            |@b       c                    @��JY�8�?             9@������������������������       �؂-؂-�?	             .@������������������������       �p=
ףp�?	             $@e       l                   �7@�H���i�?           pz@f       i                    �?�X7�_ �?�            �s@g       h                    @^N��)8�?H             \@������������������������       ��E��\�?8            @V@������������������������       �@��Z��?             7@j       k                    @�q9'��?�            @i@������������������������       �����>�?S            �`@������������������������       �      �?.             Q@m       p                    @�����?G            @[@n       o                    @��v'���?3            �T@������������������������       ��H��;��?            �B@������������������������       �V_��0��?             G@q       r                    @ƵHPS!�?             :@������������������������       ���8��8�?	             (@������������������������       �
^N��)�?             ,@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       0{@     @V@     �u@      E@      S@      :@     �X@     P�@     ��@     �N@     �S@      d@     ��@     @{@      .@     @Q@      N@      c@     �J@      g@     �H@      e@      4@     �J@      4@      C@      ^@     �d@     �@@      K@      V@     �m@     �h@       @     �B@      E@      Q@      E@     �V@       @      H@      �?      "@                     �U@     @S@      $@      *@      :@     �\@     �M@              (@      @      9@      @      A@      @      0@              @                      O@     �D@      �?      @      @      K@      .@              @              $@       @      1@              @              �?                      @@      =@      �?      �?       @      >@      @              �?              @              .@              @                                      >@      4@                       @      :@      @              �?               @              "@              @                                      7@      0@                              7@      @              �?               @              @                                                      @      @                       @      @      �?                                               @              �?              �?                       @      "@      �?      �?              @                                      �?               @              �?              �?                       @              �?      �?               @                                                                                                                      "@                               @                                      �?              1@      @      (@              @                      >@      (@              @      @      8@      $@              @              @       @      *@       @      @                                      4@      @               @              "@       @              @                       @                      �?                                      &@       @              �?              @      �?                                       @      *@       @      @                                      "@      @              �?              @      �?              @                              @      @      @              @                      $@      @               @      @      .@       @                              @              �?      @                      @                               @                              @       @                              @              @              @                                      $@      @               @      @       @      @                               @             �L@      @      @@      �?      @                      9@      B@      "@       @      3@     �N@      F@               @      @      .@       @     �I@      @      3@      �?      @                      3@      :@      �?       @      &@     �H@     �B@               @       @       @              1@      �?      "@                                      $@      .@      �?       @      $@      >@      0@              @              @              "@               @                                       @      &@      �?       @      @      8@      �?                               @               @      �?      @                                       @      @                      @      @      .@              @              �?              A@       @      $@      �?      @                      "@      &@              @      �?      3@      5@              �?       @      @              (@      �?       @              �?                      �?      �?               @               @      @              �?      �?                      6@      �?       @      �?      @                       @      $@              @      �?      &@      0@                      �?      @              @              *@                                      @      $@       @               @      (@      @                      �?      @       @       @              @                                      @      $@       @              @      $@      @                      �?      @              �?              @                                               @       @              @              @                      �?      @              �?               @                                      @       @                      �?      $@       @                              @              @              @                                      �?              @              @       @       @                              �?       @       @              @                                                      @              @      �?                                                       @               @                                      �?              �?                      �?       @                              �?       @     �W@     �D@     @^@      3@      F@      4@      C@     �@@     �V@      7@     �D@      O@     @^@      a@       @      9@     �C@     �E@      C@     �H@      1@     �I@      @      *@       @      7@      3@     �G@       @      2@      1@      Q@      J@      @      &@      2@      2@      *@     �B@      $@      D@       @      @              (@      *@      <@       @      (@      "@      <@     �B@       @      &@      (@      0@      @      =@      $@      :@       @                       @       @      .@               @      @      .@      ,@       @      @      @      "@      �?      @              3@                                      �?      @                              @       @                                              7@      $@      @       @                       @      �?      (@               @      @      "@      @       @      @      @      "@      �?       @              ,@              @              @      &@      *@       @      @      @      *@      7@              @      "@      @      @      @              @                               @       @      @              �?              &@      @              �?      �?      �?              �?              &@              @               @      @      "@       @      @      @       @      1@              @       @      @      @      (@      @      &@      @      "@       @      &@      @      3@              @       @      D@      .@      �?              @       @       @      &@      @       @      @       @       @      @      @      2@              @       @      D@      ,@                      @       @       @      &@      @      @       @       @       @      @      @      2@              @      @      6@      (@                       @      �?      @              @       @      �?                      �?      @                              �?      2@       @                       @      �?      @      �?              @              @              @              �?                                      �?      �?               @                                      �?               @              @              �?                                      �?                       @                      �?               @              @               @                                                              �?                                     �F@      8@     �Q@      ,@      ?@      2@      .@      ,@     �E@      5@      7@     �F@     �J@     @U@      @      ,@      5@      9@      9@      .@      @      5@      �?      *@      @       @      @      1@       @      $@      0@      E@      8@              @      @      "@      &@      .@      @      0@      �?      @      @      @      @      *@       @       @      "@      E@      4@               @      @       @      $@      &@      �?      *@      �?       @      @      �?      @      (@              @      @      C@      &@              �?       @      @      @      @      @      @              @              @       @      �?       @       @      @      @      "@              �?       @      @      @               @      @               @              @              @               @      @              @              �?      �?      �?      �?              �?      �?              @              �?                              �?      @                              �?                                      �?      @              �?              @              @              �?       @              @                      �?      �?      �?      >@      1@     �H@      *@      2@      .@      @      @      :@      3@      *@      =@      &@     �N@      @      &@      0@      0@      ,@      >@      1@     �G@      $@      0@      ,@      @      @      8@      1@      (@      9@      &@      M@      �?      $@       @      0@      "@      7@      @      8@       @      @       @      @      @      $@      *@      @      "@      @      <@              @      @      (@      @      @      ,@      7@       @      &@      (@      @              ,@      @      @      0@      @      >@      �?      @      �?      @      @                       @      @       @      �?                       @       @      �?      @              @      @      �?       @              @                      �?       @       @                              �?      �?                              @      @      �?      �?                                      �?      �?              �?                      �?      �?      �?      @                                      @              @     @o@      D@      f@      6@      7@      @     �N@      y@     �z@      <@      8@      R@     �v@      n@      @      @@      2@      U@      &@     �i@     �A@     �a@      1@      3@      @      D@     �u@     �w@      ;@      .@      J@     q@     �e@      @      8@      0@     �O@      @     �T@      &@     �C@      �?                      @      l@     �f@      @      @      *@      Z@      H@              @      @      1@      �?     �J@      �?      <@                              @     �f@      b@      @      @      (@     �U@      @@              �?      �?      "@      �?      D@      �?      6@                              @      c@      X@      @      @      $@     �R@      5@              �?      �?       @      �?     �@@      �?      ,@                              @      ^@     �H@      @      @      @     �I@      1@              �?      �?      @      �?      @               @                                      @@     �G@      �?              @      7@      @                              @              *@              @                               @      ?@      H@                       @      *@      &@                              �?              @              @                               @      &@     �D@                              @      @                              �?              @               @                                      4@      @                       @       @       @                                              =@      $@      &@      �?                             �D@     �C@      �?              �?      1@      0@              @      @       @               @                                                      ,@       @                               @                                                      @                                                       @       @                              �?                                                      @                                                      @                                      �?                                                      5@      $@      &@      �?                              ;@     �B@      �?              �?      .@      0@              @      @       @              "@              @                                      @      (@                              @      (@                      �?       @              (@      $@       @      �?                              4@      9@      �?              �?      $@      @              @       @      @             �^@      8@     �Y@      0@      3@      @     �A@     �^@     `h@      6@      $@     �C@      e@     �_@      @      3@      (@      G@      @     �L@       @      B@      @      @              ,@      R@      `@      "@      @      $@      U@     @P@              @       @      &@             �A@      @      3@              @              ,@      2@      M@      "@      �?      @     �@@      ?@              @              @              (@      �?      $@              �?              @      @     �B@       @               @      "@      (@                              �?              7@       @      "@              @              @      *@      5@      @      �?      @      8@      3@              @              @              6@      @      1@      @                              K@     �Q@               @      @     �I@      A@              @       @      @              *@      @      *@                                      C@     �F@              �?       @      B@      (@              @       @      @              "@      �?      @      @                              0@      9@              �?      @      .@      6@                               @             �P@      0@     �P@      *@      .@      @      5@      I@     �P@      *@      @      =@     @U@      O@      @      (@      $@     �A@      @      2@      @      *@      @       @      @      @      @@      6@      @      �?      @      ;@      9@              "@      @      @       @      0@      @      $@       @       @      @      @      =@      2@      @      �?      @      3@      2@              @              @       @       @              @      @                              @      @       @                       @      @              @      @                      H@      &@     �J@      @      *@      �?      .@      2@     �F@       @      @      :@      M@     �B@      @      @      @      @@      @      E@      &@      C@       @       @      �?      "@      (@     �D@      @      @      9@      E@      A@      @      @      @      <@       @      @              .@      @      @              @      @      @      �?      �?      �?      0@      @                              @      �?     �F@      @      B@      @      @      �?      5@      L@     �J@      �?      "@      4@     �U@     @P@      @       @       @      5@      @      @              �?                                      (@      @                              �?       @                                              @                                                      @      @                              �?       @                                                              �?                                      @       @                                                                                     �D@      @     �A@      @      @      �?      5@      F@      H@      �?      "@      4@     �U@     �O@      @       @       @      5@      @      A@       @      9@      @      @              (@     �D@      C@              @      0@     �Q@     �D@              @              ,@      @      *@       @      $@       @       @              @      @      (@               @      @      <@      8@                              �?      �?      $@       @      $@       @       @                      @      $@               @      @      8@      1@                              �?      �?      @                                              @       @       @                              @      @                                              5@              .@       @      �?              @      A@      :@              @      *@     �E@      1@              @              *@       @      .@              *@                              @      ?@      1@              @      @      >@      @              @              @       @      @               @       @      �?               @      @      "@               @       @      *@      &@                              "@              @      @      $@      �?      �?      �?      "@      @      $@      �?       @      @      .@      6@      @      @       @      @       @      @      �?      @      �?              �?       @      @      $@      �?       @      @      ,@      .@      @      @       @      @       @      @              @      �?                              �?      @      �?       @      @              @      @      @               @       @       @      �?      @                      �?       @       @      @                      �?      ,@       @      �?               @       @              �?       @      @              �?              @                                              �?      @              �?              @              �?              �?              �?              �?                                                      @                               @                       @       @                              @                                              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�v�KhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmK]hnh4h7K ��h9��R�(KK]��hu�BX         ,                   �1@rx�����?�	           ��@                           �?�x��2��?t           ؁@                           @7'�s���?�            �r@                           @7�ٔ_�?�             m@                           �?��#���?�            �g@                           �?.�܃QN�?U             _@������������������������       �V}��b�?             9@������������������������       �b�A��?B            �X@	       
                    @I��7��?,            @P@������������������������       �������?             7@������������������������       ��t��*�?             E@                           @��-]W��?            �E@                             @     ��?             @@������������������������       �R���Q�?             4@������������������������       �      �?             (@������������������������       ���ˠ�?             &@                           @<*ǩ�?'            @P@                          �0@Y�Cc�?             <@������������������������       ������H�?             "@������������������������       ������?
             3@                           @=J�L���?            �B@������������������������       �����p9�?
             3@                           @e������?             2@������������������������       ��<ݚ�?             "@������������������������       ���"e���?             "@       !                    �?�A����?�             q@                            @������?>            @Y@                          �0@6�w���?)            �P@������������������������       ����N8�?             5@                           �?J� ��w�?             G@������������������������       ���"e���?             2@������������������������       �4և����?             <@������������������������       ���� =�?             A@"       '                    @�b [I��?r            �e@#       &                    @��y4F�?6             S@$       %                     @4��\Fs�?+            �L@������������������������       �Ҋ*� �?#            �H@������������������������       �      �?              @������������������������       �"P7��?             3@(       +                    @�#%k"�?<            @X@)       *                    @=���i�?5            @U@������������������������       �~������?            �B@������������������������       �     @�?             H@������������������������       ��q�q�?             (@-       >                    @PuR���?A           �@.       =                    !@B�2D�?�            �@/       6                    �?x�z:a�?�           ؞@0       3                     �?�4�A���?B           p@1       2                    �?�H���?_             b@������������������������       ��f��I��?+             O@������������������������       ��!_ �Z�?4            �T@4       5                   �4@v�G���?�            `v@������������������������       ��^a�M<�?K            �]@������������������������       �J��I���?�             n@7       :                    �?�A���?�           ��@8       9                    �?4���?z           h�@������������������������       �s�T:��?~            �l@������������������������       �G��.��?�            �x@;       <                    @�'9K�?           ��@������������������������       ��3ژ0�?<            �@������������������������       ���V �?�            �t@������������������������       ����(\��?             $@?       N                   �6@f���*�?m           8�@@       G                    @�	K�,��?,           ��@A       D                    �?���ma�?�            �w@B       C                   �5@�d�M#�?l            �d@������������������������       �T|}��(�?\             b@������������������������       ��ˠT�?             6@E       F                   �2@{�� ��?�            �j@������������������������       ��Y ���?             K@������������������������       �fffffF�?i             d@H       K                    @�KZ�gj�?8           ~@I       J                     @��Y�=��?{            �e@������������������������       ������9�?q             d@������������������������       �����X�?
             ,@L       M                   �5@� 檪��?�            0s@������������������������       �����?�            `p@������������������������       ��Tkט��?            �F@O       V                    �?S��/��?A            @P       S                    �?%�S�<%�?�            �k@Q       R                     �?1�*���?&             I@������������������������       ������H�?             "@������������������������       ��`D�?�?            �D@T       U                     �?�Ĭ�|d�?h            @e@������������������������       ���7��d�?              I@������������������������       �:m��:�?H             ^@W       Z                   �:@�GZ�<�?�            @q@X       Y                    @DC%��N�?u             g@������������������������       ��C�3�?6            �U@������������������������       � �p?��??            �X@[       \                   �>@h����?>             W@������������������������       ���� ��?)             O@������������������������       �B��S��?             >@�t�bh�h4h7K ��h9��R�(KK]KK��h��B87       �@     �T@     `u@     �B@     �U@      7@      S@     (�@     H�@      H@     �Q@     �c@     Ђ@     @z@      4@     �U@      N@      b@      I@     �Q@      @      7@              @              @     �e@     �_@       @      @      .@      Z@      =@              �?              "@      �?      A@       @      @                              @     �\@      S@       @              @     �G@      @                              �?              ;@       @      @                              @     �X@     �I@      �?               @     �C@       @                              �?              0@       @      @                               @      U@     �E@      �?               @      A@       @                                              &@       @       @                                      M@      >@      �?               @      0@       @                                              @                                                       @      @      �?               @      @       @                                              @       @       @                                      I@      ;@                              *@                                                      @              �?                               @      :@      *@                              2@                                                                      �?                                      @      @                              $@                                                      @                                               @      4@      @                               @                                                      &@               @                               @      ,@       @                              @                                      �?              @                                               @      *@      @                              @                                      �?              @                                               @      @      @                              �?                                      �?                                                                      @      @                              @                                                      @               @                                      �?      �?                              �?                                                      @               @                                      1@      9@      �?              �?       @      @                                                              �?                                      @      2@      �?                      @                                                                                                                       @                              �?                                                                      �?                                      @      $@      �?                      @                                                      @              �?                                      *@      @                      �?      @      @                                              @              �?                                       @      @                                      @                                              @                                                      @      @                      �?      @                                                      @                                                       @      �?                               @                                                                                                              @      @                      �?       @                                                      B@      �?      0@              @              �?     �M@     �I@              @      (@     �L@      7@              �?               @      �?      7@               @              �?                      0@      $@               @      @      8@      $@                              @      �?      3@               @              �?                      $@      @               @       @      6@      @                              �?              @                                                      @      �?                               @       @                                              *@               @              �?                      @      @               @       @      ,@      �?                              �?              @                                                      @                               @      @                                                      @               @              �?                              @               @              $@      �?                              �?              @              @                                      @      @                      �?       @      @                               @      �?      *@      �?       @               @              �?     �E@     �D@              @      "@     �@@      *@              �?              @              @      �?      @                              �?      8@      2@              @      @      @      @                              @              @      �?      @                              �?      3@      .@              @      @      @      @                                              @      �?       @                              �?      2@      (@               @       @      @      @                                                              �?                                      �?      @              �?       @                                                              @                                                      @      @                               @       @                              @              @              @               @                      3@      7@                      @      :@       @              �?               @              @              @               @                      1@      5@                      @      :@      @              �?              �?              �?               @               @                      @      (@                              *@      @                                               @              @                                      ,@      "@                      @      *@                      �?              �?              @                                                       @       @                                      @                              �?              {@      T@     �s@     �B@      U@      7@     �Q@     pu@     �|@      G@     �P@     �a@      @     px@      4@     @U@      N@      a@     �H@     �p@     �G@      i@      :@     �Q@      4@      K@     �]@     �m@      @@     �J@     @W@     �p@     @o@      ,@     �N@      F@     �V@     �B@     0p@     �G@      i@      :@     @Q@      4@      K@     �]@     �m@      @@      J@     @W@     �p@     @o@      ,@     �M@      F@     �V@     �B@     �Q@      .@     �D@       @      ,@              &@      A@      M@      @      2@      :@     @W@     �G@              1@      .@      6@      .@      4@      "@      $@       @       @               @      @      .@              @      @     �E@      @              @       @      @      @      $@      @      @                                       @      @              @      �?      7@      @               @       @      �?      �?      $@      @      @       @       @               @       @      "@               @      @      4@      @               @              @      @      I@      @      ?@              (@              "@      >@     �E@      @      (@      4@      I@      D@              *@      *@      .@      "@      *@      �?      @              �?              �?      ,@      :@      �?       @      $@      *@      *@              $@      �?      @      @     �B@      @      ;@              &@               @      0@      1@      @      $@      $@     �B@      ;@              @      (@      (@      @     �g@      @@      d@      8@     �K@      4@     �E@     @U@     `f@      ;@      A@     �P@      f@     `i@      ,@      E@      =@     @Q@      6@     �X@      2@     @Q@      �?      6@      @      .@     �G@     �T@      @      (@      6@     �V@     @R@      @      4@      .@      4@      @     �F@      "@      1@               @      �?      @      0@      <@      @      @      (@      ?@      8@      @      @              .@       @     �J@      "@      J@      �?      ,@       @      &@      ?@     �K@              @      $@     �M@     �H@      �?      ,@      .@      @      @     �V@      ,@     �V@      7@     �@@      1@      <@      C@      X@      8@      6@     �F@     �U@     @`@      $@      6@      ,@     �H@      0@     @R@      (@     �F@      3@      2@      (@      &@      ;@      M@      .@       @      ;@     �N@      R@      @      (@      @      9@       @      2@       @      G@      @      .@      @      1@      &@      C@      "@      ,@      2@      :@      M@      @      $@       @      8@       @      @                              �?                                              �?                                       @                              e@     �@@     �]@      &@      ,@      @      1@      l@     �k@      ,@      *@     �H@     �l@     �a@      @      8@      0@     �F@      (@     �\@      (@      K@      @       @              *@     `e@      b@      @       @      :@     @d@     �V@              .@      @      :@      @     �F@      @      B@      @                      @     �P@      I@       @      @      ,@     �W@     �B@              @      @       @      @      2@      �?      (@      �?                      �?      A@      9@      �?      @      @      J@      &@                      @       @              2@      �?      (@      �?                      �?      <@      3@      �?      @      @      G@      "@                      �?       @                                                                      @      @                              @       @                       @                      ;@       @      8@       @                      @      @@      9@      �?       @      &@     �E@      :@              @              @      @       @              &@                               @       @      �?      �?                      1@      @                                              3@       @      *@       @                      �?      8@      8@               @      &@      :@      4@              @              @      @     �Q@      "@      2@      @       @              "@     @Z@     �W@       @      @      (@     �P@     �J@              "@      @      2@      @      3@      @      @      �?                              L@      D@       @      �?              8@      0@               @              @      �?      0@      @      @                                      K@      D@       @      �?              4@      ,@               @              @              @              �?      �?                               @                                      @       @                                      �?     �I@      @      ,@      @       @              "@     �H@      K@               @      (@     �E@     �B@              @      @      .@       @     �H@      @       @               @              @     �G@      G@               @      &@      B@      <@              @      @      &@       @       @              @      @                      @       @       @                      �?      @      "@                              @              K@      5@      P@      @      (@      @      @     �J@     @S@      $@      @      7@     �P@     �I@      @      "@      $@      3@      @      :@      "@      :@       @      @              �?      B@      E@              @      (@      7@      8@              @              @      �?      @      @      @              �?              �?      @      2@                      �?      @      @                                              �?              @                              �?      �?       @                                      �?                                              @      @      �?              �?                      @      0@                      �?      @      @                                              3@      @      6@       @      @                      =@      8@              @      &@      3@      4@              @              @      �?      &@              @                                      @      @                      �?      @      ,@              �?               @               @      @      .@       @      @                      9@      3@              @      $@      ,@      @              @              @      �?      <@      (@      C@       @      @      @      @      1@     �A@      $@      �?      &@     �E@      ;@      @      @      $@      ,@      @      0@      @      :@      �?      @               @      1@      9@      @              @      D@      .@      @      @      @      @              @      �?      0@      �?       @               @       @      1@      @              �?      *@      @               @      �?      @              &@      @      $@              @                      "@       @      �?              @      ;@       @      @       @      @      �?              (@       @      (@      �?      �?      @      �?              $@      @      �?      @      @      (@      �?      �?      @       @      @      $@      @      @      �?                                      @      @      �?      @       @      &@      �?      �?      @      @      @       @       @      @              �?      @      �?              @                      @      �?      �?                              @        �t�bub��      hhubh)��}�(hhhhhKhKhKhG        hh.hNhJXC)hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         @                     @ݪ�M���?�	           ��@       !                    �?׮i�?�           B�@                          �2@N�K3��?#           $�@                            �?��_���?�            �u@                           @�6�+��?F            �\@                           @��9k��?1            @T@������������������������       ��U���H�?            �J@������������������������       �����S��?             <@	       
                   �1@� =[y�?             A@������������������������       ��0�*�?             9@������������������������       ��2�tk~�?             "@                           @%�V�?�            �l@                           @     T�?(             P@������������������������       ��^����?            �A@������������������������       �d����?             =@                           @��-�?n            �d@������������������������       �LXdp|��?9            @U@������������������������       �XntX�?5            @T@                          �5@�� �JH�?G           ��@                            �?��f�>�?�             x@                            �?���x�?�            �r@������������������������       �c����?X            `a@������������������������       �g����?`            �c@                           @Q������?7            @V@������������������������       �{	�%���?,             R@������������������������       �|�l�]�?             1@                          �:@yo�ñ�?X           p�@                           @Ԯ�(!�?�            �x@������������������������       �HQU"�?}            �i@������������������������       �QH�Cf�?y            �g@                           �>@D��sS�?b            �d@������������������������       �9��8���?@             [@������������������������       ����L���?"            �L@"       1                   �5@gч����?�           `�@#       *                    @��?�           x�@$       '                    �?��Ƕ�?�            0t@%       &                   �2@tJV�B�?�            �k@������������������������       ���J;�?@            �X@������������������������       ������?P            �^@(       )                   �0@/lu�(�?C            @Y@������������������������       �      �?             0@������������������������       ��D��8��?7            @U@+       .                   �2@@(�t|R�?           �z@,       -                    @jվI��?{            `i@������������������������       �<҂�@�?Y            �a@������������������������       ����c���?"            �O@/       0                    @j���ґ�?�             l@������������������������       ��G��?`            @b@������������������������       �Li��X�?1            �S@2       9                    @y�7�vf�?�           H�@3       6                     �?:8�w_�?�           ��@4       5                   �9@�重+H�?�            �o@������������������������       ���T�?T            @`@������������������������       �
�:$x}�?N             _@7       8                     �?��J��?�?�            `u@������������������������       �2G����?�             j@������������������������       ��CQ7;�?[            �`@:       =                   �:@7(
���?6            @U@;       <                     �?캮뺮�?             E@������������������������       �{�G�z�?             4@������������������������       �,�Ra���?             6@>       ?                    @b@��MP�?            �E@������������������������       �6�h$��?             >@������������������������       �؉�؉��?             *@A       X                    @�>q;E��?�           ��@B       Q                    @N�x&�?           �@C       J                    �?j�)/'��?�           ��@D       G                    �?|y�����?�            @p@E       F                    �?     ��?)             P@������������������������       �KKKKKK�?             A@������������������������       �6�h$��?             >@H       I                    �?��I���?�            �h@������������������������       ��q�a�?:             X@������������������������       �!�rh���?G             Y@K       N                    �?��p����?�            �w@L       M                   �2@�.�s�?X             c@������������������������       �p�u=q��?             G@������������������������       �2��M��?>            �Z@O       P                    @:(g����?�            `l@������������������������       �o_Y�K�?!             J@������������������������       �Eoax_��?l            �e@R       W                    @]��<�"�?�            @l@S       V                   �=@�����?�             j@T       U                    �?��2w��?u            �g@������������������������       ��.�6�G�?             G@������������������������       ��n����?X            �a@������������������������       �(������?             3@������������������������       ����Hx�?
             2@Y       h                   �5@:ފ,CF�?�            pt@Z       a                    �?�,-j��?�            �l@[       ^                    �?�F1-C�??            @X@\       ]                    @���d;�?            �D@������������������������       �v��`��?             =@������������������������       �r�q��?	             (@_       `                    @N��)x9�?$             L@������������������������       ��@�Y��?             =@������������������������       ��&y��?             ;@b       e                    �?��P�4 �?F            �`@c       d                    @��&�l��?$            �P@������������������������       �������?            �F@������������������������       �ŕ�(�?             5@f       g                   �3@Ӏ����?"            �P@������������������������       �!XA�H�?            �J@������������������������       �����W�?             *@i       n                    �?c`x�OR�?A            �X@j       k                    @,�2���?             ?@������������������������       �      �?              @l       m                   �9@K����?             7@������������������������       ��1G����?             *@������������������������       �>
ףp=�?             $@o       r                    �?�%o��?.            �P@p       q                   �8@��ɒ�z�?             ;@������������������������       ��T�x?r�?
             &@������������������������       �     @�?
             0@������������������������       ��p=
ף�?             D@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       �|@     @U@     �t@      =@      U@      7@      T@     �@     �@     �R@     @U@     `f@     ��@     �y@      *@      P@     �P@     �^@     �N@     0t@     �K@     �l@      (@      G@      @      O@      |@     P}@     �M@      N@     �]@     0x@     `n@      @     �E@      C@     �S@      C@      c@      4@     �V@       @      ,@              6@     �p@     Pq@      &@     �@@      E@      f@     �\@              ,@      "@      <@      ,@      =@      @      "@                              @     ``@     �Z@      �?       @      @      C@      ,@                              �?              "@       @       @                              �?     �A@     �F@              �?      @      (@      @                              �?               @               @                              �?      6@      B@              �?      @      @      �?                              �?               @               @                                      2@      3@              �?      �?      @      �?                                                                                              �?      @      1@                      @       @                                      �?              �?       @                                              *@      "@                              @       @                                                                                                      $@       @                              @                                                      �?       @                                              @      �?                                       @                                              4@      �?      @                              @      X@      O@      �?      �?       @      :@      &@                                              *@              @                                      1@      6@              �?       @      @      �?                                               @              �?                                      ,@      .@                               @      �?                                              &@               @                                      @      @              �?       @      @                                                      @      �?      @                              @     �S@      D@      �?                      5@      $@                                               @      �?      �?                              @     �G@      ,@                              (@      @                                              @              @                                      @@      :@      �?                      "@      @                                             �^@      1@     @T@       @      ,@              2@     @a@     @e@      $@      ?@      B@     `a@     @Y@              ,@      "@      ;@      ,@     �H@       @      9@               @              @      U@     �S@      @      @      0@     �P@      @@              @              @       @     �E@       @      5@              �?              @      H@      O@      @      @      (@      L@      9@              @              @       @      9@              @              �?                      5@      8@      @      @      (@      9@      *@              @              �?              2@       @      ,@                              @      ;@      C@       @       @              ?@      (@               @               @       @      @              @              �?                      B@      1@              �?      @      $@      @                              @              @              @                                      <@      1@                      @      @      @                              @              �?                              �?                       @                      �?              @       @                                             �R@      .@      L@       @      (@              (@      K@     �V@      @      8@      4@     @R@     @Q@              "@      "@      5@      (@     �I@       @      J@              @              @      E@     �R@              ,@      $@     �I@      K@              @      @      $@      @      :@      @      C@              @               @      (@      :@               @      @      >@      @@              @      @      @      @      9@      @      ,@                              @      >@      H@              @      @      5@      6@               @      �?      @              7@      @      @       @       @              @      (@      1@      @      $@      $@      6@      .@               @       @      &@      "@      .@      @       @       @       @              @      $@      ,@      �?      @       @      2@      @                      �?      @      @       @      �?       @                              @       @      @      @      @       @      @      &@               @      �?      @      @     `e@     �A@     �a@      $@      @@      @      D@     �f@      h@      H@      ;@      S@     @j@      `@      @      =@      =@      I@      8@     �[@      "@     �K@      �?      @      �?      1@     �a@     �a@      @      &@     �A@     �Z@     @P@              "@      @      4@      ,@      J@      �?      C@              @      �?      &@     �D@     �N@       @      @      $@     �C@      B@               @              &@      "@     �B@      �?      :@               @              "@      :@     �B@       @      @      $@      ?@      3@               @              $@      @      ,@              @               @               @      2@      2@       @       @       @      8@      @                              @       @      7@      �?      6@                              @       @      3@               @       @      @      *@               @              @      @      .@              (@               @      �?       @      .@      8@              �?               @      1@                              �?      @                                                              @      &@                              �?      �?                                              .@              (@               @      �?       @      (@      *@              �?              @      0@                              �?      @      M@       @      1@      �?      @              @      Y@     �T@      �?      @      9@      Q@      =@              @      @      "@      @      <@      @      @                               @      O@      ?@      �?      @      @     �@@      *@              @              @              $@      @      @                              �?     �J@      6@      �?      @      @      7@      &@                              �?              2@       @      �?                              �?      "@      "@                              $@       @              @              @              >@       @      $@      �?      @              @      C@     �I@              @      4@     �A@      0@              �?      @      @      @      4@      �?      @                                      ?@     �B@               @      &@      5@      $@              �?              @       @      $@      �?      @      �?      @              @      @      ,@              �?      "@      ,@      @                      @              @     �N@      :@     �U@      "@      9@      @      7@      D@     �H@     �F@      0@     �D@     �Y@     �O@      @      4@      :@      >@      $@      J@      :@     �Q@      @      6@      @      0@      @@     �D@     �E@      ,@     �C@      X@      K@      @      1@      8@      ;@       @      *@      *@      C@       @      &@      @      "@      "@      $@      1@       @      1@      D@      8@      �?       @      1@      &@      @      &@      "@      @@      �?       @      �?      @      @      @      @      @      @      8@      "@               @      @      @               @      @      @      �?      "@       @      @      @      @      $@      @      ,@      0@      .@      �?      @      &@      @      @     �C@      *@      @@      @      &@      �?      @      7@      ?@      :@      @      6@      L@      >@      @      "@      @      0@      @      8@      @      3@       @      @              @      5@      6@      0@      @      *@      @@      3@              @      �?      &@      @      .@       @      *@      @      @      �?      @       @      "@      $@       @      "@      8@      &@      @       @      @      @       @      "@              0@       @      @              @       @       @       @       @       @      @      "@              @       @      @       @       @              &@       @       @                       @      @               @      �?      @      @               @               @      �?      �?              @       @                              @      �?               @      �?      �?      @               @                      �?      �?               @               @                      @       @                               @                                       @              @              @              �?              @              @       @              �?      @      @              �?       @      �?      �?      @               @              �?              @              @       @              �?      �?      @              �?       @              �?                      @                              @                                              @       @                              �?              a@      >@      Y@      1@      C@      2@      2@     @X@      e@      .@      9@     �N@     �e@     �d@      "@      5@      <@     �F@      7@     �Y@      5@     �Q@      .@      @@      0@      1@     �G@     �]@      ,@      4@      G@      ^@      _@      @      1@      7@      B@      5@     �S@      0@     �E@       @      9@      ,@       @      @@     �Y@      *@      1@     �A@     �W@      V@      @      0@      .@      2@      *@      @@      &@      3@              1@      @              &@      G@       @      @      $@      =@     �B@              $@      @      $@      @      "@      @      @              �?                      @      *@      @      @      @      @      @              @      �?              �?      "@      @      @                                      @      @       @      �?       @      �?                      @                                      �?                      �?                      �?      @      @       @       @      @      @               @      �?              �?      7@      @      0@              0@      @              @     �@@       @      @      @      7@      A@              @      @      $@      @      (@              @              @       @              @      .@              �?              0@      8@              @              @       @      &@      @      $@              &@       @               @      2@       @       @      @      @      $@              �?      @      @      @      G@      @      8@       @       @      $@       @      5@     �L@      @      &@      9@     @P@     �I@      @      @      &@       @      @      6@              (@      �?      @      @      @      $@      :@              @      *@      ;@      &@                      @       @      @       @               @                                      @      @                       @      4@                                       @              ,@              $@      �?      @      @      @      @      4@              @      &@      @      &@                      @              @      8@      @      (@      @      @      @      @      &@      ?@      @      @      (@      C@      D@      @      @      @      @       @      @                      �?      �?      �?      �?      @      @                      @      (@      @      @       @              @              4@      @      (@      @       @      @      @      @      8@      @      @      @      :@     �A@              @      @               @      9@      @      ;@      @      @       @      "@      .@      .@      �?      @      &@      :@      B@       @      �?       @      2@       @      4@      @      ;@      @      @      �?      "@      .@      .@      �?      @      "@      7@     �@@       @      �?       @      2@       @      3@      @      :@      @       @              "@      .@      .@      �?      @      "@      6@     �@@              �?      @      0@       @       @               @                               @       @      �?      �?       @      �?      @      @                      @       @      @      &@      @      2@      @       @              @      *@      ,@              �?       @      1@      :@              �?              ,@      @      �?              �?       @      @      �?                                                      �?               @              @       @              @       @               @              �?                                               @      @      @                                              A@      "@      >@       @      @       @      �?      I@      I@      �?      @      .@     �K@     �E@      @      @      @      "@       @      :@              9@       @      @                      G@      C@              @      ,@     �C@      6@              �?              @       @      .@              *@       @                              1@      "@              @      �?      1@      2@                              �?      �?       @               @                                       @      @                               @      "@                              �?              �?              @                                      @      @                              @      @                              �?              �?              �?                                       @                                       @      @                                              *@              @       @                              "@      @              @      �?      "@      "@                                      �?       @                      �?                              �?      @              @      �?      @      @                                      �?      @              @      �?                               @                                      @      @                                              &@              (@              @                      =@      =@               @      *@      6@      @              �?              @      �?      "@              @                                      7@      "@               @              &@      @              �?              @               @              @                                      *@      @               @              "@       @              �?                              �?              �?                                      $@       @                               @       @                              @               @               @              @                      @      4@                      *@      &@                                      �?      �?      �?              @              @                      @      4@                      $@      @                                      �?      �?      �?              @                                                                      @      @                                                       @      "@      @               @       @      �?      @      (@      �?              �?      0@      5@      @      @      @      @              �?      @                      �?              �?               @                      �?      @      @                      @       @              �?      @                                                      �?                                      @                                                       @                      �?              �?              @                      �?      @                              @       @                                                              �?              @                               @                              @                               @                      �?                               @                      �?       @                                       @              @      @      @              �?       @              @      @      �?                      (@      2@      @      @               @               @      @      �?                                       @      @      �?                      @      @              @              �?                              �?                                       @       @      �?                      �?      @                              �?               @      @                                                       @                              @                      @                              @      �?      @              �?       @               @                                      @      .@      @                      �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         :                   �2@ 8����?�	           ��@                           �?(�d�n�?�           T�@                           �?&1w�Ǐ�?B           �@       	                    �?P�W
���?P            �`@                          �1@�q�q\�?             H@                            �?�Cc}h��?             <@������������������������       �؉�؉��?             *@������������������������       �{�G�z�?	             .@������������������������       ��(\����?             4@
                           �?�3_<�?5             U@                           @4և����?            �A@������������������������       ��E]t��?             6@������������������������       �pƵHP�?             *@                           @!i���t�?"            �H@������������������������       ���!pc�?             6@������������������������       ��.sxQ��?             ;@                            @2���?�            �w@                           @�4�V͝�?�            �s@                            �?k�y�ʍ�?n             g@������������������������       ��c�B�?(            @Q@������������������������       �x������?F            �\@                            �?D!ޮ��?U            @`@������������������������       �     ��?             @@������������������������       ��d�(��?>            �X@                           @'T����?/             Q@                           @�� wKn�?             5@������������������������       �h/�����?             "@������������������������       ��q�q�?             (@                            @^1��d��?!            �G@������������������������       �0�w¹��?             5@������������������������       ���1G���?             :@        /                     @�`�6���?O           ��@!       (                    @�QG>�)�?�            �u@"       %                    @�sPR�?{            @g@#       $                   �1@Q��)���?V            �^@������������������������       ��EƐ�K�?2            @S@������������������������       ��)F�?$            �F@&       '                   �0@     ��?%             P@������������������������       ��m۶m��?             ,@������������������������       ��$��C�?             I@)       ,                    @
ףp=��?b             d@*       +                    @$���U�?>            @Y@������������������������       �`��� ��?            �J@������������������������       �r�qG�?             H@-       .                   �0@���~��?$            �M@������������������������       ����k���?             &@������������������������       �r�q��?             H@0       3                   �0@f�1�?r             g@1       2                    @�Cc}�?             <@������������������������       �n�����?             2@������������������������       ����Q��?             $@4       7                    @�7f	�?`            �c@5       6                   �1@1�qfg��?E            �]@������������������������       �b*
/�?             �L@������������������������       ���Gӹ�?%            �N@8       9                    �?��n=���?            �C@������������������������       �     ��?	             0@������������������������       ��_�����?             7@;       X                    �?m��}��?            h�@<       K                     @1M�3`�?            ��@=       D                   �7@�:��?.           ��@>       A                   �5@���4c�?a           p�@?       @                    @��� � �?�            �w@������������������������       ���>91�?�            �n@������������������������       �J�{���?Z            �`@B       C                     �?VDu����?w             f@������������������������       ��'2�ޟ�?\            �a@������������������������       ����
�?            �B@E       H                    @�����?�            s@F       G                    �?6��t{�?�            @q@������������������������       �;'u�?D            �X@������������������������       �������?r             f@I       J                    @���Rp�?             =@������������������������       ����c���?             5@������������������������       �      �?              @L       S                    @���(Ɣ�?�            Px@M       P                    �?u9	h���?�            �q@N       O                    @�:G��?)            �L@������������������������       ��{~���?!            �G@������������������������       �
ףp=
�?             $@Q       R                    �?�c��?�            �l@������������������������       �M�a���?(            �P@������������������������       �ylւͷ�?\            `d@T       W                   �:@d��'�T�?E            �Y@U       V                    @�x�����?=            �V@������������������������       �T�r
^N�?             <@������������������������       �T�
�	�?-             O@������������������������       ��q�q�?             (@Y       h                    �?�����K�?            @�@Z       a                    �?�Q譂|�?�           0�@[       ^                     �?���A�)�?�            �q@\       ]                    �?V����?b            `d@������������������������       �<<<<<<�?             A@������������������������       �����m�?L             `@_       `                     @�xPy���?K            @]@������������������������       �S�f��?             C@������������������������       ��)J����?3            �S@b       e                    @Xw�T��?C           �~@c       d                    @��v�|�?�            r@������������������������       �*%�fox�?�            �k@������������������������       �S��a`��?.            �P@f       g                   �=@ą�+.�?�            �i@������������������������       �촜�ׇ�?p            �d@������������������������       ����#E��?            �D@i       p                    @Ԏah��?           P�@j       m                   �8@<�l=t�?v           ��@k       l                    @Q6���?           �z@������������������������       ����!�?�            p@������������������������       �W�v����?b            �d@n       o                    @�Q1t4�?k            �e@������������������������       �d�%
�?^            @c@������������������������       �lv�"��?             5@q       t                     �?>�6H�/�?�            `n@r       s                    �?t{����?\            �b@������������������������       �������?             K@������������������������       �\L|bp�?=            �W@u       v                     @��_Drf�?>            �W@������������������������       �,\&�Y�?            �G@������������������������       �i�����?            �G@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       �|@     �R@     �t@      C@      R@      <@     @T@     X�@     �@      P@     @W@      e@     Ђ@     �y@      (@     �Q@     �N@     @`@      I@      ^@      @      Q@      �?      @              $@     s@      j@       @      &@      9@      e@     �P@              (@      @      7@      @     �L@      �?      :@                              �?     `h@     �\@              �?      (@     �R@      4@              @              @              7@      �?      @                                     �D@      0@                      @      :@      @              @              @              ,@              @                                      &@      @                      @      @      �?              @              @              "@              @                                      $@       @                      @              �?                                              @              @                                      @       @                                      �?                                              @                                                      @                              @                                                              @                                                      �?      �?                              @                      @              @              "@      �?      @                                      >@      *@                              7@      @                                              @              �?                                      $@      @                              $@      @                                              @                                                      $@                                      @      @                                              �?              �?                                              @                              @                                                      @      �?      @                                      4@      @                              *@      �?                                              �?      �?                                              (@      @                              @                                                      @              @                                       @      @                               @      �?                                              A@              3@                              �?     @c@     �X@              �?      "@     �H@      .@                              �?              9@              @                              �?     @a@     @V@              �?      "@     �@@      $@                              �?              ,@              @                              �?     �V@      I@              �?      @      ,@      @                              �?              @              @                                      8@      :@              �?      @      @                                      �?              "@              �?                              �?     �P@      8@                              $@      @                                              &@              @                                      H@     �C@                      @      3@      @                                               @                                                      &@      .@                      �?      �?       @                                              "@              @                                     �B@      8@                      @      2@      @                                              "@              (@                                      0@      $@                              0@      @                                               @                                                      �?      @                              *@       @                                               @                                                                                              @       @                                                                                                      �?      @                               @                                                      @              (@                                      .@      @                              @      @                                                              &@                                      @      @                              @                                                      @              �?                                      (@      @                                      @                                             �O@      @      E@      �?      @              "@     �[@     �W@       @      $@      *@     @W@      G@               @      @      0@      @      D@      @      1@                              "@     �T@     �Q@       @      @      $@     �M@      ;@              @      �?      @       @      3@       @      .@                              @      ;@      D@       @      @      @      E@      .@                              �?       @      .@       @       @                               @      4@      1@      @      @      @     �A@      @                              �?       @      &@       @      @                              �?      *@      (@              @       @      8@      @                                       @      @              @                              �?      @      @      @               @      &@      @                              �?              @              @                              @      @      7@       @               @      @       @                                               @                                                      �?      &@                                                                                       @              @                              @      @      (@       @               @      @       @                                              5@       @       @                              @     �K@      >@                      @      1@      (@              @      �?      @              &@                                                      H@      6@                      �?      &@      @                              �?               @                                                      >@      ,@                                      �?                                              @                                                      2@       @                      �?      &@      @                              �?              $@       @       @                              @      @       @                      @      @      @              @      �?      @              @                                                       @       @                                                                                      @       @       @                              @      @      @                      @      @      @              @      �?      @              7@      �?      9@      �?      @                      <@      8@              @      @      A@      3@              �?       @      "@      @      @                               @                      "@       @                              �?      @                                              @                               @                       @      @                                       @                                                                                                      @      �?                              �?      �?                                              2@      �?      9@      �?      @                      3@      0@              @      @     �@@      0@              �?       @      "@      @      .@      �?      ,@      �?      @                      0@      "@              @      �?      ;@      .@                       @       @      �?      $@              @              @                      $@       @                      �?      ,@      @                       @      @              @      �?      "@      �?                              @      @              @              *@      $@                              @      �?      @              &@                                      @      @               @       @      @      �?              �?              �?       @      �?              $@                                      �?       @                      �?      �?                                                       @              �?                                       @      @               @      �?      @      �?              �?              �?       @     0u@     @Q@     �p@     �B@     �P@      <@     �Q@     �q@      w@      L@     �T@     �a@      {@     �u@      (@      M@      M@     �Z@     �F@      c@      ;@     @[@      @      1@      @      :@     �d@     �i@      (@      C@      I@     �j@     �a@       @      ,@      :@     �@@      (@      [@      4@     �R@       @      @              1@     ``@      d@       @      :@      =@      `@     �Y@               @      "@      :@      @     �R@       @      F@      �?      @              "@     @Z@     �]@      @      "@      2@     �X@      F@              @       @      &@      @      L@      @      7@      �?      @              @     @T@     �T@      @      @      $@     @Q@      6@              @              "@      �?      C@       @      ,@      �?                      @      C@     �J@       @      @      @     �J@      *@              @              "@      �?      2@      �?      "@              @                     �E@      >@       @      �?      @      0@      "@                                              2@      @      5@              �?               @      8@      B@              @       @      =@      6@              �?       @       @       @      .@      @      ,@              �?               @      7@      @@              @      @      1@      3@              �?       @      �?       @      @      �?      @                                      �?      @                      @      (@      @                              �?              A@      (@      >@      �?       @               @      :@      E@      @      1@      &@      >@     �M@              @      @      .@      @      >@      (@      9@      �?      �?              @      4@      E@      @      1@      &@      8@     �L@              @      @      ,@      @      .@      @      @                              @      ,@      1@      �?      @      @       @      (@              �?      �?      @              .@      @      2@      �?      �?                      @      9@      @      *@       @      0@     �F@               @      @      $@      @      @              @              �?              @      @                                      @       @                              �?      �?       @              @              �?              @      @                                      @       @                              �?               @               @                                                                              @                                              �?      F@      @     �A@       @      &@      @      "@      B@     �E@      @      (@      5@      U@     �C@       @      @      1@      @      @      A@      @      @@       @      "@      @      @      7@     �B@       @       @      3@     �J@      ;@       @      @      1@      �?      @      @      �?      "@                      �?      �?      @      *@       @      �?      @      @      @              �?       @              �?      @      �?      "@                      �?              @      (@       @      �?      @       @      @              �?       @              �?                                                      �?      �?      �?                              @      @                                              >@       @      7@       @      "@      @      @      1@      8@              @      0@     �G@      5@       @       @      .@      �?      @      0@      �?      @              @                       @      &@                              ,@       @      �?                      �?      �?      ,@      �?      4@       @      @      @      @      "@      *@              @      0@     �@@      *@      �?       @      .@               @      $@      @      @               @              @      *@      @       @      @       @      ?@      (@              @              @      �?      $@       @      @               @              @      *@      @       @      @       @      7@      (@               @              @      �?       @       @                       @                      @       @                              &@      �?                              @      �?       @              @                              @      "@      @       @      @       @      (@      &@               @               @                       @                                                                                       @                      �?              �?             `g@      E@     �c@     �@@      I@      7@     �F@     �\@     �d@      F@      F@     @W@     �k@     `i@      $@      F@      @@     �R@     �@@     @R@      :@     �V@      &@      A@      3@      5@      5@     �K@      8@      @@      K@     @W@      Z@      @      :@      6@     �C@      7@      C@      @      @@       @      .@      @      $@      "@      2@      $@      @      3@      E@     �@@              @       @      &@      &@      7@      @      3@       @      &@      @      @      @       @      @       @       @      A@      &@              @       @      @      "@      @               @               @              @              @                      �?      @      @              �?       @       @              3@      @      1@       @      "@      @      @      @      @      @       @      @      =@      @              @              @      "@      .@              *@              @              @      @      $@      @      @      &@       @      6@              @      @      @       @       @              @               @                              @       @      �?      @      @       @                      �?      �?              *@              @               @              @      @      @      @      @      @      @      ,@              @      @      @       @     �A@      4@     �M@      "@      3@      0@      &@      (@     �B@      ,@      :@     �A@     �I@     �Q@      @      3@      ,@      <@      (@      :@      &@      B@      @      .@      "@      @      "@     �@@      "@       @      ,@      ?@      A@      @      "@      @      1@      @      0@      @      9@      @      ,@      @      @       @      ;@      @      @      $@      8@      <@      @      @      @      1@      @      $@      @      &@       @      �?       @              �?      @      @      @      @      @      @               @                      @      "@      "@      7@      @      @      @      @      @      @      @      2@      5@      4@     �B@      �?      $@       @      &@      @      "@      "@      4@      @      @      �?      @      @       @      @      &@      ,@      4@     �B@              $@               @       @                      @      �?              @                       @              @      @                      �?               @      @      @     �\@      0@     @P@      6@      0@      @      8@     �W@     �[@      4@      (@     �C@      `@     �X@      @      2@      $@     �A@      $@      W@       @      B@      ,@      "@      @      (@     �R@     �W@      ,@      (@      6@     @X@     �O@      @      "@      @      6@      @     �R@      @      8@      "@      @              @     @Q@     @S@      @      @      *@      Q@      D@      �?      @       @      &@      @      ?@      @      2@      @      @              @      F@     �E@       @      @      $@     �C@     �@@              �?              @      @     �E@      �?      @       @                              9@      A@      @       @      @      =@      @      �?      @       @      @      �?      2@      @      (@      @      @      @      @      @      2@      "@      @      "@      =@      7@       @      @      @      &@              (@      @      (@      @       @      @      @      @      0@       @      @      "@      =@      5@       @      @      @      @              @                               @              �?               @      �?                               @              �?              @              6@       @      =@       @      @              (@      3@      0@      @              1@      @@      B@      �?      "@      @      *@      @      $@      @      6@      @      @              @      .@      (@      @              0@      4@      ,@              @      @      @      �?       @              @              �?              @      @      @      @               @      *@      @               @              �?               @      @      0@      @      @              @       @      @      �?              ,@      @       @              �?      @      @      �?      (@      @      @      @       @              @      @      @       @              �?      (@      6@      �?      @              @      @      $@      @      @      @                              �?      �?       @                      �?      (@              @              @      @       @      �?       @               @              @      @      @                      �?      &@      $@      �?      @              @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��zhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         8                    �?YfB>x�?�	           ��@                           �?v8ߌ���?�           8�@                          �3@*���h�?�           ��@                          �1@�q�q��?q             h@                           @��N�p��?/            �U@                           �?"-@/w��?             �P@������������������������       ����2j��?            �I@������������������������       �l�l��?
             .@	       
                   �0@4և����?             5@������������������������       �      �?              @������������������������       ��(ݾ�z�?	             *@                           �?���H��?B            @Z@                           �?��;�\`�?             E@������������������������       �����>4�?             ,@������������������������       �$I�$I��?             <@                          �2@���nJ~�?&            �O@������������������������       ����+	�?            �@@������������������������       ��?�P�a�?             >@                          �?@�z�f��?"           0}@                           �?�Fy@n�?           �{@                           @�*+�j!�?b            �c@������������������������       �OX~�L�?G            �\@������������������������       �Y�����?             F@                           �?b�2�t[�?�             r@������������������������       ��u�B��?D            �\@������������������������       �x7�_��?p            �e@                           @      �?             4@������������������������       �*L�9��?             &@������������������������       ������H�?             "@       +                    �?+��\�?[           ؍@       &                   �<@R�绹�?�            w@        #                   �7@8��;a�?�             u@!       "                    @N�QD�T�?�            `m@������������������������       �|z3���?g             e@������������������������       ��z�� �?)            �P@$       %                    @./�<���?=            @Y@������������������������       ��5�h�?6            @U@������������������������       �      �?             0@'       *                   �?@vK�B#��?            �@@(       )                   �=@�&%�ݒ�?             5@������������������������       ��zv��?             &@������������������������       �
ףp=
�?             $@������������������������       �r�q��?             (@,       1                     @��$�?y           P�@-       0                    @b�؞�0�?�            �r@.       /                     �?F�V15�?�            0r@������������������������       ��T����?m            @e@������������������������       ����s�@�?U            @^@������������������������       �      �?              @2       5                   �5@�qӸ��?�            �q@3       4                   �0@<ݚ��?X             b@������������������������       �ffffff�?             $@������������������������       �(�?=���?R            �`@6       7                    �?']����?Y            �a@������������������������       ���F�� �?             ;@������������������������       ��Ϧ���?G             ]@9       X                     @0�ܫ���?�           ��@:       I                   �4@1��Չ�?q           �@;       B                    �?�3Dz��?E           ،@<       ?                    @�MK<��?8           p~@=       >                   �2@�!7p��?�            p@������������������������       �x�>�M��?`            �b@������������������������       ���P6�?@            �Z@@       A                   �0@tQ-���?�            �l@������������������������       ��:y�z��?             �H@������������������������       �+7̺W��?x            �f@C       F                     �?������?           @{@D       E                     �?�f��Z�?�            `s@������������������������       �ر�4���?a            @d@������������������������       ��%G$n�?a            �b@G       H                    @�����?K            �_@������������������������       ��趱��?=            �Z@������������������������       ��p=
ף�?             4@J       Q                    �?ח��+k�?,           X�@K       N                   �;@�8���?�            �q@L       M                    @����<�?�             o@������������������������       ��n1��?q            @g@������������������������       �����?)            �O@O       P                   �=@8�q_��?            �@@������������������������       ��"w����?             3@������������������������       �^N��)x�?             ,@R       U                    @�Y�ܓ�?}           ��@S       T                    @@��]#�?G            �\@������������������������       �_Y�K�?#             J@������������������������       �8։'�?$            �O@V       W                    @z�u�?6           �}@������������������������       ��.n�<�?            y@������������������������       �!�����?0            �S@Y       f                    �?���=�q�?0           P@Z       a                    @�`���?s            �g@[       ^                   �5@m_!'1�?>            �X@\       ]                    �?e	wX�r�?.            �Q@������������������������       �6YE�?            �@@������������������������       ����}��?             C@_       `                   �9@[\!	V��?             ;@������������������������       �     @�?	             0@������������������������       �F]t�E�?             &@b       c                    �?x�|&�?5            �V@������������������������       �x�(�?            �F@d       e                    �?���U_�?             G@������������������������       �     p�?             @@������������������������       ���>4և�?             ,@g       l                    @	�kā�?�            �s@h       k                    @E����\�?_            �c@i       j                    @���m���?T            �`@������������������������       ��}�l^�?4            �T@������������������������       �������?              J@������������������������       ������?             7@m       p                   �2@*��-��?^            @c@n       o                    �?���#�F�?             E@������������������������       �<+	���?             .@������������������������       �L�t��>�?             ;@q       r                    �?
^N��i�?A             \@������������������������       �]�I���?            �K@������������������������       �/�s��?#            �L@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       �}@     �U@     Pv@      <@      Q@      4@     @S@     ��@     ؃@      Q@     �Q@     �c@     ��@     Py@      @      P@      ?@     �_@     �P@     �k@      G@     �d@      @     �E@      .@     �@@     �W@     `j@     �B@     �F@     @U@     �o@     �f@       @      E@      6@     �P@      F@     @V@      ,@     �M@       @      $@      @      *@      N@      Y@      @      3@     �@@     �`@      M@      �?      1@      "@      5@      (@      9@      @       @                                     �E@      F@      �?       @      @      C@      $@              @              @      @      1@              @                                      9@      1@                      @      .@      @                                              0@              �?                                      5@      $@                      @      *@      �?                                              (@              �?                                      2@       @                      @      @      �?                                              @                                                      @       @                              @                                                      �?              @                                      @      @                               @       @                                                               @                                      �?       @                              �?       @                                              �?              @                                      @      @                              �?                                                       @      @       @                                      2@      ;@      �?       @      �?      7@      @              @              @      @      @                                                      "@      @      �?      �?      �?      (@      @               @               @                                                                      @      @                                       @               @                              @                                                      @      @      �?      �?      �?      (@       @                               @              @      @       @                                      "@      4@              �?              &@      @              �?              @      @      @      @                                              @      *@                              @      �?              �?              @              �?               @                                      @      @              �?               @       @                              �?      @      P@      $@     �I@       @      $@      @      *@      1@      L@      @      1@      <@     �W@      H@      �?      ,@      "@      .@      "@      O@      $@      I@       @       @      @      $@      1@     �K@      @      0@      <@     �W@      F@              (@      "@      .@      "@      1@      @      "@                       @       @      "@      ;@      @       @      (@     �B@      ,@              @      �?      @      @      (@       @      "@                       @      �?      @      6@      @       @      (@      6@      @               @      �?       @      @      @      �?                                      �?      @      @                              .@      @               @              @             �F@      @     �D@       @       @      �?       @       @      <@               @      0@     �L@      >@               @       @      $@      @      >@      @      $@      �?      @               @      @      *@              �?      @      <@      &@               @               @              .@      @      ?@      �?      @      �?      @      @      .@              @      *@      =@      3@              @       @       @      @       @              �?               @              @              �?      @      �?                      @      �?       @                              �?                                                                      @      �?                      @               @                              �?              �?               @              @              �?                                              �?                                     �`@      @@     �Z@      @     �@@      (@      4@     �A@     �[@      >@      :@      J@     �^@      _@      �?      9@      *@      G@      @@     @Q@      .@      @@              *@       @      @      (@      E@      *@       @      3@     �M@      ?@              @      @      6@      .@      Q@      &@      ;@              $@       @       @      (@     �D@      *@      @      0@     �M@      >@              @      @      2@      *@      H@       @      5@              @               @      &@      C@      $@       @      *@      A@      1@               @      @      $@      "@     �B@       @       @              @              �?      $@      ?@      @       @      @      :@      *@               @      @      @       @      &@              *@                              �?      �?      @      @              @       @      @                       @      @      �?      4@      @      @              @       @              �?      @      @      @      @      9@      *@               @               @      @      (@      @      @              @       @              �?      @      @      @      @      5@      *@               @              @      @       @               @                                                                              @                                       @              �?      @      @              @              @              �?              @      @              �?               @      �?      @       @              @      @                              @              �?                      @              �?                      �?       @       @                      @                                              �?                      @                                               @       @              @      �?                              @                                                      �?                      �?                      �?              �?              @                                              @                                       @               @             �O@      1@     �R@      @      4@      $@      .@      7@     @Q@      1@      2@     �@@     �O@     @W@      �?      3@      @      8@      1@     �A@      @      B@       @      @      �?      &@      2@      D@      ,@      @      2@      <@     �B@      �?      *@      @      0@       @     �A@      @      B@       @      @      �?      &@      2@     �C@      *@      @      2@      <@      @@      �?      *@      @      0@       @      2@      @      7@              @      �?      @      @      8@      @       @      "@      3@      7@      �?      @      �?      &@      @      1@              *@       @      @              @      (@      .@       @       @      "@      "@      "@              @      @      @       @                                                                      �?      �?      �?                      @                                              <@      *@      C@      �?      *@      "@      @      @      =@      @      *@      .@     �A@      L@              @       @       @      "@      7@      @      1@      �?      @       @      @      @      1@       @      @      �?      <@      :@               @              @              @       @                                              �?                                              @                                              3@      @      1@      �?      @       @      @      @      1@       @      @      �?      <@      7@               @              @              @      @      5@              "@      @      �?              (@      �?      $@      ,@      @      >@              @       @      @      "@      �?      �?      @              @      @                       @                              �?      �?                      �?              @      @      @      0@              @      @      �?              $@      �?      $@      ,@      @      =@              @      �?      @      @     `o@     �D@      h@      7@      9@      @      F@     p{@     �z@      ?@      9@     @R@      x@     �k@      @      6@      "@      N@      7@     �i@      >@     `b@      1@      2@      @      =@     @w@     �v@      6@      4@      G@     r@     �b@       @      0@       @     �D@      .@     �Z@      @     �F@      @       @              @     @q@     `j@      @      @      0@     @b@      O@              @      @      1@      @      I@       @      0@      �?                      @     �d@     �_@      @      @       @      T@      :@              �?              @              =@       @      @      �?                      @     �Q@     �Q@      @       @      @     �C@      2@                              @              .@       @       @                               @      J@      I@              �?      @      0@      @                                              ,@              @      �?                       @      3@      5@      @      �?      @      7@      &@                              @              5@              "@                                     @W@     �K@              �?      �?     �D@       @              �?                               @              �?                                      @@      "@                              @                                                      3@               @                                     �N@      G@              �?      �?      B@       @              �?                             �L@      @      =@      @       @              @      \@     @U@       @      �?       @     �P@      B@               @      @      ,@      @      E@      @      .@      @      �?               @      O@     �P@      �?      �?       @      I@      =@               @      @      &@      @      5@       @      @      @      �?              �?     �D@     �@@      �?      �?      @      :@      $@              �?      �?      @       @      5@       @      "@                              �?      5@      A@                      @      8@      3@              �?      @      @      @      .@              ,@              �?              �?      I@      2@      �?                      0@      @                              @              $@              *@              �?              �?      H@      0@      �?                      "@      @                              @              @              �?                                       @       @                              @      @                                             �X@      8@     �Y@      &@      0@      @      6@      X@     �c@      1@      0@      >@     �a@      V@       @      *@      @      8@      "@      :@      ,@      >@      �?               @       @      8@     @R@      @       @      @      F@      @@              @      �?       @      @      9@      $@      =@                               @      8@     @Q@      @      @      @      B@      >@              @              �?      �?      0@      @      4@                              @      2@      M@      �?      @      @      >@      4@               @                              "@      @      "@                               @      @      &@       @                      @      $@              @              �?      �?      �?      @      �?      �?               @                      @              @      �?       @       @                      �?      �?       @      �?       @      �?                                              @              @      �?      @                                               @               @              �?               @                                                      @       @                      �?      �?             @R@      $@      R@      $@      0@      �?      ,@      R@     �T@      ,@       @      8@     �X@      L@       @       @      @      6@      @      2@      @      2@      @                       @      7@      "@      �?      �?      @       @      ,@              �?       @      @              *@      @      @      �?                      �?      @      @      �?      �?      @      @      @                      �?       @              @      �?      (@       @                      �?      1@      @                       @      @      "@              �?      �?       @             �K@      @      K@      @      0@      �?      (@     �H@     �R@      *@      @      1@     �V@      E@       @      @      �?      2@      @     �F@      @     �A@      @      *@      �?      @     �C@     @Q@      (@      @      1@     �T@      D@       @      @              ,@      @      $@              3@       @      @              @      $@      @      �?       @              "@       @              @      �?      @      �?     �F@      &@     �F@      @      @       @      .@     �P@     �L@      "@      @      ;@     �W@     @R@      @      @      �?      3@       @      :@      @      1@      @      @      �?      �?      ,@      <@               @      (@     �C@      >@              �?              @       @      1@       @      @      @       @      �?              @      *@               @      $@      4@      $@                              @       @      $@      �?      @      @              �?              @      &@               @      @      3@      @                              �?       @      @               @                      �?              @      @                              &@       @                                              @      �?      @      @                                      @               @      @       @       @                              �?       @      @      �?      �?               @                               @                      @      �?      @                               @              @      �?                       @                              �?                                      @                                              �?              �?                                              �?                      @      �?                                       @              "@       @      &@               @              �?      @      .@                       @      3@      4@              �?               @              @      �?      @                                      @      ,@                               @      (@                                              @      �?       @               @              �?      @      �?                       @      &@       @              �?               @               @      �?      @               @              �?      @      �?                       @      "@       @              �?               @              @              @                                                                               @      @                                              3@      @      <@      @      @      �?      ,@     �J@      =@      "@      @      .@      L@     �E@      @      @      �?      ,@      @       @      �?      0@      @       @              @      1@      1@       @      �?      &@      B@      3@       @      �?      �?      @      @      @      �?      *@      @                      @      1@      1@      @               @      A@      1@       @      �?      �?      @      @      @      �?      @       @                       @      *@      *@      @              �?      5@      (@       @      �?                      @      �?               @      �?                      @      @      @                      @      *@      @                      �?      @      �?      @              @               @              �?                      @      �?      @       @       @                                              &@      @      (@              �?      �?       @      B@      (@      �?       @      @      4@      8@      �?      @              $@      �?      @              @                                      5@      @                              @      �?                              �?      �?      @               @                                      @      �?                                      �?                                              �?              �?                                      ,@      @                              @                                      �?      �?      @      @      "@              �?      �?       @      .@      @      �?       @      @      1@      7@      �?      @              "@               @              @                              @      ,@      �?      �?       @       @      @      $@              @              @              @      @      @              �?      �?      @      �?      @                       @      &@      *@      �?                      @        �t�bub��(     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�-�yhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         @                     @&9��Ƀ�?�	           ��@       !                    �?���/�?�           �@                          �2@�,���4�?*           �@                            �?Nd���?�            Pw@                           �?
鬶]�?X            `a@                           �?*L�9��?            �@@������������������������       ��)O�?             2@������������������������       ��h$���?             .@	       
                    @������??            �Z@������������������������       �8cU�3�?+            @Q@������������������������       �9g�9���?            �B@                          �1@�������?�            @m@                           @%W��e��?b            �a@������������������������       �^�4�,�?H            @X@������������������������       ��a%����?            �E@                            �?��e���?9            �W@������������������������       �paRC4%�?            �I@������������������������       �RB)��.�?            �E@                           @E�����?7           8�@                          �6@�k�X��?           �y@                           @������?}            �g@������������������������       ��c�ZB�?@             Y@������������������������       ������?=             V@                           �?v�X,�Z�?�            @l@������������������������       �����<��?*            �P@������������������������       ����Q�?j             d@                           @�-*z"��?&           �~@                           >@��~j��?�             u@������������������������       ��7�/�t�?�            @t@������������������������       �X�Cc�?             ,@                             �?��X��?_            �b@������������������������       �"�D�g��?A            �Y@������������������������       �m%A����?            �H@"       1                    �?�����?�           <�@#       *                    �?ig.�+�?W           x�@$       '                     �?ML	��H�?`            `d@%       &                    �?p�j���?.            �S@������������������������       ���<,��?             9@������������������������       �F�ǧ�?            �J@(       )                    �?�b��L�?2            @U@������������������������       �D��2(�?             F@������������������������       �ĭ[F�?            �D@+       .                    @eę�L�?�            �x@,       -                    �?l<�1�'�?@            �Z@������������������������       ��Z=;n�?             F@������������������������       �|m�SF��?"             O@/       0                    �?��oh�?�             r@������������������������       ���1+��?E             [@������������������������       ���/Y3;�?r            �f@2       9                    @=�R4S�?:            �@3       6                   �3@������?�           (�@4       5                   �0@�/����?�            p@������������������������       ���j;�?            �F@������������������������       ����ƥ�?�            �j@7       8                    @��׎�t�?            @x@������������������������       ���QS�?�             l@������������������������       ��7����?j            `d@:       =                    @�H�m�?�            `k@;       <                   �1@\�tӸ�?q            �c@������������������������       �d���+��?             :@������������������������       �q��s0��?a            ``@>       ?                    @��f��I�?$             O@������������������������       ���ˠ�?             F@������������������������       ��E��ӭ�?             2@A       Z                    �?�`�A �?�           ��@B       K                    �?4�/�r�?A           �@C       D                   �2@�S�v��?{            �i@������������������������       �а�����?%            �N@E       H                   �6@M��;�?V            �a@F       G                    @��S����?-             S@������������������������       �ndG�+�?%             O@������������������������       ��m۶m��?             ,@I       J                   �;@c����?)            �P@������������������������       ����V�/�?             I@������������������������       �躍`3�?
             1@L       S                    @Vڵ��?�            ps@M       P                    �?*0����?�            �k@N       O                   �6@�������?            �E@������������������������       �F]t�E�?            �@@������������������������       �
ףp=
�?             $@Q       R                   �;@>���]��?p            `f@������������������������       �?�ƨBR�?_             c@������������������������       ��P���?             ;@T       W                    @]��bC��?:            @V@U       V                   �1@UUUUU��?             H@������������������������       �~h����?             ,@������������������������       ����.L�?             A@X       Y                   �3@V?B���?            �D@������������������������       �*L�9��?	             &@������������������������       �1u��A��?             >@[       h                   �4@���K�+�?�           ؅@\       c                    @�Ʊ��S�?�            �t@]       `                   �1@��7x,�?�            �q@^       _                   �0@U��`�?9            �W@������������������������       �p�u=q��?             7@������������������������       ��&7bv�?(            �Q@a       b                   �2@�0�J���?x             h@������������������������       �m��
I��?&             K@������������������������       ��+�W��?R            `a@d       e                    @A�@���?             �E@������������������������       �      �?
             0@f       g                    �?���d�?             ;@������������������������       �ƵHPS!�?
             *@������������������������       �������?             ,@i       n                    @���)�i�?�            w@j       m                   �@@�`so�y�?�            �r@k       l                   �>@��v��b�?�            �q@������������������������       �d�N&�T�?�            0p@������������������������       �2G�����?             :@������������������������       �b���i��?             &@o       r                   �;@R�U��U�?0            @R@p       q                    @n�T�~`�?'             M@������������������������       ��"��Q�?             E@������������������������       �     ��?             0@������������������������       ��h$���?	             .@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       @{@     �S@     �v@      E@      P@      ?@      T@     ��@     �@     �H@     �V@     `e@     (�@     �|@      $@     �L@     �F@      _@     �B@     �r@      E@     `n@      8@      C@       @     �I@     �{@     `}@      ?@      L@     @Y@     �z@     0r@       @      A@      >@      U@      1@      a@      0@     �W@      @      "@              4@      q@     �p@      @      1@      =@     �k@      a@              &@      @      8@      @     �C@      @      @                              �?     @c@     �R@               @      "@     �N@      3@                              @              2@      @      @                              �?      F@     �A@              �?      @      5@      @                              @              $@      �?       @                                      &@       @                              @                                                      @               @                                      @      �?                              @                                                      @      �?                                              @      �?                              @                                                       @       @      �?                              �?     �@@     �@@              �?      @      ,@      @                              @              @       @      �?                                      >@      0@              �?      �?      &@      @                                              @                                              �?      @      1@                       @      @      @                              @              5@              @                                     �[@     �C@              �?      @      D@      *@                                              .@              �?                                      O@      9@                      @      >@       @                                              @              �?                                      I@      4@                       @      .@       @                                               @                                                      (@      @                      @      .@                                                      @              @                                      H@      ,@              �?      �?      $@      &@                                              @                                                      9@      @              �?              @      "@                                              @              @                                      7@       @                      �?      @       @                                             �X@      *@     �U@      @      "@              3@      ^@      h@      @      .@      4@      d@     @]@              &@      @      4@      @      J@       @     �L@      �?      @              @      =@      Q@      �?      "@      *@     @S@     �L@              $@       @      ,@      @      4@       @      3@              @              @      2@      D@               @      @      H@      6@               @              @      �?      @      �?      &@                              �?      $@      7@              �?      @      ;@      1@                               @      �?      1@      �?       @              @              @       @      1@              �?      �?      5@      @               @              �?              @@      @      C@      �?      @               @      &@      <@      �?      @      "@      =@     �A@               @       @      &@      @      @      @      @              �?                       @      &@      �?      @              0@       @              @      �?       @              :@      @      ?@      �?       @               @      "@      1@               @      "@      *@      ;@              @      �?      "@      @      G@      @      >@      @      @              *@     �V@      _@      @      @      @      U@      N@              �?      @      @      �?      4@      @      2@              @              *@     �O@     @W@      @      @      @      O@      D@                      @      @              4@      @      0@              @              *@     �O@     @W@      @      @      @     �N@      >@                      @      @                               @                                                      �?                      �?      $@                                              :@       @      (@      @                              <@      ?@               @      @      6@      4@              �?                      �?      .@              $@      @                              2@      8@              �?      @       @      2@              �?                      �?      &@       @       @                                      $@      @              �?              ,@       @                                             �d@      :@     �b@      4@      =@       @      ?@     �e@     �i@      8@     �C@      R@     �i@     `c@       @      7@      9@      N@      (@     @P@      &@     �Q@      "@      4@      @      ,@      E@      I@      (@      6@     �@@      R@     @R@      �?      &@      &@      =@      $@      @@              ,@              @              @      0@      6@       @       @       @      5@      6@      �?               @       @      @      $@              @              @                      @      (@       @       @      @      (@      "@      �?               @       @              �?              �?                                      @      @               @      @      �?      @                               @              "@              @              @                      �?      @       @               @      &@      @      �?               @      @              6@               @               @              @      &@      $@                       @      "@      *@                                      @      .@               @               @              @      �?      @                      �?      @      @                                       @      @              @                               @      $@      @                      �?      @      @                                      �?     �@@      &@      L@      "@      .@      @      "@      :@      <@      $@      4@      9@     �I@     �I@              &@      "@      5@      @      @      @      1@               @              @      @      @      �?      @      �?      8@      .@              @       @      @      �?      @      �?      $@                                      �?                              �?      1@      @               @                      �?              @      @               @              @      @      @      �?      @              @      "@              @       @      @              <@      @     �C@      "@      *@      @      @      4@      5@      "@      0@      8@      ;@      B@              @      @      2@      @      $@      @      *@              @      �?      @      @      $@      @      @      (@      1@      "@                      @       @      @      2@      �?      :@      "@      $@      @       @      0@      &@      @      *@      (@      $@      ;@              @      @      $@       @     @Y@      .@     �S@      &@      "@      @      1@     @`@     @c@      (@      1@     �C@     �`@     �T@      �?      (@      ,@      ?@       @     �P@      @     �K@      @      @      @      &@      [@      a@      $@      .@      7@     �Z@      P@      �?       @      @      .@       @      ?@              (@                              �?     @P@     @R@      @      @      @     �C@      .@              �?              @      �?      @                                                      &@      "@                      @      $@      @                              @              <@              (@                              �?      K@      P@      @      @      @      =@      "@              �?                      �?      B@      @     �E@      @      @      @      $@     �E@     �O@      @      &@      0@     �P@     �H@      �?      @      @      (@      �?      9@      @     �B@      @              @      @      7@      :@      @      @      "@      A@     �A@              @      @      @              &@      @      @      �?      @      �?      @      4@     �B@      �?      @      @     �@@      ,@      �?      @       @      @      �?      A@      "@      8@      @      @              @      6@      2@       @       @      0@      <@      2@              @      "@      0@              7@       @      7@      @       @              @      0@      .@       @              @      8@      (@              �?      @      @              "@      @                                              �?      @                              @                                                      ,@      @      7@      @       @              @      .@       @       @              @      2@      (@              �?      @      @              &@      �?      �?               @                      @      @               @      $@      @      @              @      @      $@              @      �?      �?               @                      @       @               @      @       @      @              @      @      @              @                                                              �?                      @       @      @                              @             �`@     �B@     �]@      2@      :@      7@      =@     �\@     �`@      2@      A@     �Q@      g@     �d@       @      7@      .@      D@      4@      M@      @      E@      @      (@      @      ,@     �Q@     �Q@      @      *@      .@      X@     �N@              $@      @      0@      @      ?@      @      4@              @                      :@      =@       @       @      @      >@     �E@              @              @      �?      .@       @       @                                      *@      @       @                       @      @                              @              0@      @      (@              @                      *@      7@               @      @      6@     �C@              @               @      �?       @              @               @                      (@      *@                              (@      <@                               @      �?       @              @               @                      &@      *@                              $@      1@                               @      �?                                                              �?                                       @      &@                                              ,@      @       @               @                      �?      $@               @      @      $@      &@              @                               @       @       @               @                      �?      $@                      @      @      "@                                              @      �?                                                                       @              @       @              @                              ;@      �?      6@      @       @      @      ,@     �F@      E@      @      &@      (@     �P@      2@              @      @      &@      @      1@              .@      @       @      @      *@      7@      @@      �?      @      &@      I@      .@              @      @      @      @      �?                                      �?      @      $@      @                      �?      *@       @              �?              @              �?                                                      $@      @                              *@      �?              �?              @                                                      �?      @              @                      �?              �?                                              0@              .@      @       @      @      "@      *@      9@      �?      @      $@     �B@      *@              @      @              @      *@              (@      @      �?      @      @      *@      6@      �?      @      $@      B@      $@              �?      @              @      @              @              @               @              @                              �?      @              @      �?              �?      $@      �?      @                              �?      6@      $@      @      @      �?      0@      @               @               @               @      �?      @                                      1@      @              @              @      �?                              �?              @              �?                                      @                                                                                               @      �?      @                                      $@      @              @              @      �?                              �?               @              @                              �?      @      @      @      �?      �?      "@       @               @              @                                                                      �?      @              �?      �?      �?      �?              �?                               @              @                              �?      @              @                       @      �?              �?              @             �R@      ?@     @S@      (@      ,@      3@      .@     �E@      P@      (@      5@     �K@     @V@     �Z@       @      *@       @      8@      *@      K@      @      F@      @      @              @      @@      =@      �?      @      ,@      K@      H@              @      @      &@      @     �I@      @      E@      @      @              @      5@      5@      �?      @      *@      G@     �F@               @      @      $@      @      0@      �?       @               @                      .@       @              @      @      @      8@               @              @              "@      �?      �?              �?                      @      �?                                      @                                              @              @              �?                      "@      @              @      @      @      4@               @              @             �A@      @      A@      @       @              @      @      *@      �?      @       @     �D@      5@                      @      @      @      @      @      0@                                      @      @              �?              $@      @                              �?       @      =@      @      2@      @       @              @       @      @      �?       @       @      ?@      0@                      @      @       @      @               @                              �?      &@       @                      �?       @      @              @              �?      �?      �?                                                       @       @                      �?      @                                              �?       @               @                              �?      @      @                              @      @              @              �?               @                                              �?       @                                       @      @              @                                               @                                      �?      @                              @                      �?              �?              5@      8@     �@@       @      $@      3@      "@      &@     �A@      &@      ,@     �D@     �A@      M@       @      @      @      *@       @      .@      &@      ?@       @      "@      3@      @      @      8@      &@      ,@      B@      3@      G@       @      @      @      (@       @      .@      &@      ?@       @       @      3@      @      @      8@      &@      (@      A@      3@      G@      @      @      @      (@      @      .@      &@      >@      @       @      ,@      @      @      7@       @      &@      >@      3@      E@      @      @      @      (@      @                      �?      �?              @              @      �?      @      �?      @              @              @                                                              �?                                               @       @                      @                              �?      @      *@       @              �?               @      @      &@                      @      0@      (@                              �?              @      "@      �?              �?              �?      @      $@                      @      $@      (@                              �?              @      @      �?              �?                      @       @                      @      "@      @                                                      @                                      �?      �?       @                              �?      @                              �?               @      @      �?                              �?              �?                              @                                                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���8hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         :                    �?"������?�	           ��@                           �?*�M�!�?�           ��@                            @k�iژ�?�           �@                            �?y?r��5�?�             v@                          �5@����_R�?�            �s@                           @�"����?]            �a@������������������������       ��"�Ȳy�?V            �`@������������������������       ������H�?             "@	       
                    �?�o�5��?q            @e@������������������������       �������?,            �O@������������������������       ���SNY��?E            �Z@                          �3@���\��?            �C@������������������������       ���ˠ�?             &@                          �8@�)x9/�?             <@������������������������       ��E��ӭ�?             2@������������������������       ��G�z��?             $@                          �;@I�b���?�             r@                           �?�BE���?�             o@                           �?�5$``�?4            @T@������������������������       �X�<ݚ�?             B@������������������������       �~X�<��?            �F@                          �5@sBI:P�?o            �d@������������������������       �r�q��?@             X@������������������������       ����Ր�?/            �Q@                           �?�r
^N��?             E@������������������������       ��������?             (@������������������������       ��z�G��?             >@       +                     �?���ҟS�?N           ��@       $                   �2@\ж�N�?           �|@       !                    �?�G�zT�?2             T@                           �1@     ��?             @@������������������������       ��ˠT�?             &@������������������������       �Z�eY�e�?             5@"       #                     �?UUUUU��?             H@������������������������       �� ˔xG�?            �A@������������������������       ��T�6|��?             *@%       (                   �:@����@�?�            �w@&       '                     �?׷�s���?�            @q@������������������������       �8"��Wf�?_            �d@������������������������       ��h�EE��?D            �[@)       *                     �?�� 8o��?B            �Y@������������������������       �Dc}h��?-            �Q@������������������������       �     P�?             @@,       3                     @
]�e�?�?7            @-       0                    �?��U"t.�?-            �S@.       /                   �6@v��`��?             =@������������������������       �      �?
             0@������������������������       ��(ݾ�z�?             *@1       2                   �6@���YՏ�?            �H@������������������������       �J���#��?             6@������������������������       ��:���?             ;@4       7                   �9@N���8a�?
           @z@5       6                    �?� �M��?�            t@������������������������       ����pk��?9            �U@������������������������       �ް�Q���?�            `m@8       9                    �?�00s���?9            �X@������������������������       �L�9���?             6@������������������������       ��:� �z�?-            @S@;       Z                   �5@�� ���?�           �@<       K                    �?��$����?y           |�@=       D                   �1@�rl�P�?�           (�@>       A                    @z������?�            �o@?       @                     @�F�����?r             g@������������������������       �������?`            �c@������������������������       �/�����?             <@B       C                     �?`��q�?+            �P@������������������������       �2(&ޏ�?             6@������������������������       ��ks����?            �F@E       H                   �4@�P���?+           �~@F       G                     �?��\�d��?�            �v@������������������������       �O
�|�s�?6            @V@������������������������       ��oB���?�             q@I       J                    @     ��?E             `@������������������������       ��D�����?             5@������������������������       �������?:            �Z@L       S                     @�tnښ�?�           Ѕ@M       P                   �4@�؃�7l�?K           @�@N       O                   �1@�B�5�?            {@������������������������       ��اh�I�?_            `b@������������������������       �	�Şxy�?�            �q@Q       R                     �?;n,�R�?2             V@������������������������       �θ	�?             :@������������������������       ��y��A�?!             O@T       W                    �?�G�v�?f            @f@U       V                   �3@F�&�;�?(            �Q@������������������������       �UUUUUU�?             H@������������������������       ��7�A�?             6@X       Y                    @k絊��?>             [@������������������������       ��?1            @U@������������������������       �'�%����?             7@[       j                    �?o�J	k��?            `�@\       c                     �?L	���#�?�            �x@]       `                    @`����x�?�             m@^       _                    @ɉa���?l            `d@������������������������       �i��A���?<            @U@������������������������       �8��,�?0            �S@a       b                    @4�	~���?-            @Q@������������������������       �F�{0X��?            �A@������������������������       �r������?             A@d       g                     @�2t5�?e            �d@e       f                    @���>�?8            @W@������������������������       �DU(Ǐ��?,            �Q@������������������������       ��Ҍ���?             7@h       i                   �8@F������?-            �Q@������������������������       �|>�+78�?            �A@������������������������       �������?             B@k       r                    @��Q���?"            ~@l       o                     @괨���?�             u@m       n                    @Ю���?�            �q@������������������������       ���$�W�?z            `i@������������������������       �:"�*���?/            �T@p       q                    @	j*D�?             J@������������������������       �G���H�?             5@������������������������       �[�>��?             ?@s       v                   �>@�������?^            �a@t       u                    @��3L?l�?U            �_@������������������������       �����~�?J             \@������������������������       ��K~���?             .@������������������������       ��o^M<+�?	             .@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       `~@      T@     Pu@      ?@     @S@      ?@     �Q@     �@     �@     �M@      U@      g@     x�@     }@      1@     @Q@      B@     �\@      M@     �i@     �B@     �e@      5@      J@      6@      =@     �[@      d@      B@     �J@     �W@     `k@     @j@      $@     �C@      6@      M@      F@      X@      2@     �O@              $@              0@      O@      V@      $@      .@      >@     �Y@     �S@      @      *@      &@      ,@      *@     �P@      .@      B@              @              $@      C@      J@      @      $@      "@     �K@     �A@              @      @      @      @      L@      .@     �@@              @              $@      ?@      G@      @      "@      @      H@     �@@              @      @      @      @     �A@      �?      $@                              @      <@      4@       @       @       @      =@      @              �?              �?      �?      @@      �?      "@                              @      ;@      3@       @               @      =@      @              �?              �?      �?      @              �?                                      �?      �?               @                      �?                                              5@      ,@      7@              @              @      @      :@       @      @      @      3@      :@               @      @      @      @      (@       @      @                                       @      0@       @      @              $@      "@              �?      �?                      "@      (@      4@              @              @      �?      $@               @      @      "@      1@              �?      @      @      @      $@              @                                      @      @      �?      �?       @      @       @                                              @                                                      �?      �?                      �?       @                                                      @              @                                      @      @      �?      �?      �?      @       @                                               @              �?                                      @      @              �?      �?      �?       @                                               @               @                                              �?      �?                      @                                                      >@      @      ;@              @              @      8@      B@      @      @      5@     �G@     �E@      @      $@      @       @       @      5@      @      8@              @              @      8@      B@      @       @      4@      F@      A@       @      @      @       @      @       @               @                                      *@      ,@      @              "@      "@      (@              @              @      �?       @              �?                                      @      @      @              @      �?      @              @              �?                              �?                                      "@       @                      @       @      "@               @               @      �?      *@      @      6@              @              @      &@      6@               @      &@     �A@      6@       @       @      @      @      @      @       @      .@               @              �?      @      &@              �?      "@      9@      (@              �?              @       @      "@      �?      @              �?              @      @      &@              �?       @      $@      $@       @      �?      @              �?      "@              @              @              �?                              @      �?      @      "@      �?      @      �?              @      @               @                                                              @               @                                                      @              �?              @              �?                                      �?      �?      "@      �?      @      �?              @     �[@      3@     @[@      5@      E@      6@      *@     �H@     @R@      :@      C@     @P@     @]@     �`@      @      :@      &@      F@      ?@     @P@       @      I@      @      1@       @      (@      ;@     �C@      *@      4@      >@     �J@     �K@      @      0@      @      1@      ,@      @               @                              �?      (@      2@      �?      �?      @      1@      @                               @      @      @              @                                      @      "@                      @      @                                       @              @                                                      @      @                      �?      �?                                                      �?              @                                              @                      @      @                                       @              �?              @                              �?      "@      "@      �?      �?      �?      *@      @                                      @      �?              �?                              �?      @      @      �?      �?      �?      &@      @                                      @                       @                                      @       @                               @                                              @      N@       @      E@      @      1@       @      &@      .@      5@      (@      3@      8@      B@      J@      @      0@      @      .@       @      J@      @     �B@      @      "@              @      *@      0@      @      &@      &@     �@@     �F@      @      @      �?      *@      @      7@      @      ?@      @      @              @      "@      (@      @      @      @      9@      7@      @      �?      �?      "@       @      =@       @      @              @              @      @      @       @      @      @       @      6@              @              @      @       @       @      @       @       @       @      @       @      @      @       @      *@      @      @              &@      @       @       @      @       @       @      �?       @       @      @              @      �?       @       @       @      @              &@      �?       @       @      @              @      �?                       @       @       @      @              @      �?      @                      @                      G@      &@     �M@      .@      9@      ,@      �?      6@      A@      *@      2@     �A@      P@     @S@      @      $@      @      ;@      1@      $@              $@              @                      @      @      �?      �?      @      ,@      ,@                      �?      @      @      @                              @                      @      @                              @      @                                              @                                                      @      @                              @       @                                              @                              @                                                              @       @                                              @              $@                                      �?      �?      �?      �?      @      @      $@                      �?      @      @      @              @                                      �?      �?                      @      @                                       @                              @                                                      �?      �?       @      @      $@                      �?      @      @      B@      &@     �H@      .@      6@      ,@      �?      0@      >@      (@      1@      =@      I@     �O@      @      $@      @      6@      ,@      B@      "@      C@      @      *@      @      �?      .@      ;@       @      (@      5@      E@     �K@              @      @      5@      @      (@      �?      @               @                      @      $@      @      @      @      ,@      (@                       @      @      @      8@       @     �@@      @      &@      @      �?      "@      1@      @      @      2@      <@     �E@              @       @      .@      �?               @      &@      "@      "@      "@              �?      @      @      @       @       @       @      @      @      �?      �?      $@                      @               @                      �?              �?              �?      �?      @               @                      @               @      @      "@      @      "@                      @      @      @      @      @      @      @      @      �?      �?      @     pq@     �E@      e@      $@      9@      "@     �D@     �x@      |@      7@      ?@     �V@     @w@     �o@      @      >@      ,@      L@      ,@      h@      .@     �X@       @      @      �?      6@     �t@     Ps@       @      0@     �I@      n@      \@              $@      @      0@      @     �W@      @     �B@               @               @     �j@      e@      @      $@      5@     @]@     �G@              @      �?      @             �@@              @                              �?      X@      Q@              �?      @     �C@      @                              �?              5@              @                              �?     �T@      C@              �?      @     �@@      �?                                              0@              �?                              �?     @S@      ?@              �?      @      9@      �?                                              @               @                                      @      @                               @                                                      (@              �?                                      *@      >@                       @      @       @                              �?              �?                                                      @      0@                              �?                                      �?              &@              �?                                      $@      ,@                       @      @       @                                              O@      @     �@@               @              @     �]@      Y@      @      "@      .@     �S@      F@              @      �?      @             �H@      @      5@                               @     @V@     @S@      @      @      *@      H@     �D@              @              @              &@      @      @                                      5@      >@                      @      @      @                                              C@      �?      1@                               @      Q@     �G@      @      @      @      E@      A@              @              @              *@      �?      (@               @              @      >@      7@      @      @       @      >@      @                      �?                       @              @                                               @                              *@                                                      &@      �?       @               @              @      >@      5@      @      @       @      1@      @                      �?                     �X@      $@      O@       @      @      �?      ,@     @\@     �a@       @      @      >@     �^@     @P@              @      @      $@      @     �S@      @      ?@              @      �?      "@     �W@     @\@       @      @      4@      U@     �G@              @      @      $@      @     �O@      @      3@              @              @     �V@     �V@       @      @      1@     �Q@     �E@              @      @      "@      @      1@      @      @                              �?     �A@     �D@              @      @      4@      (@                              �?              G@       @      (@              @              @     �K@      I@       @      �?      $@      I@      ?@              @      @       @      @      .@       @      (@                      �?      @      @      6@               @      @      ,@      @                              �?      @       @              "@                      �?      @      @      @                               @      �?                              �?              *@       @      @                              �?      �?      2@               @      @      (@      @                                      @      4@      @      ?@       @      �?              @      3@      <@                      $@     �C@      2@               @                              *@      @      .@                              @      @      @                      @      ,@      @                                              @              .@                              @      @      @                       @       @      @                                              @      @                                               @                              @      @      �?                                              @              0@       @      �?               @      *@      7@                      @      9@      *@               @                              @              *@       @      �?               @      &@      (@                      @      5@      *@                                              �?              @                                       @      &@                              @                       @                             �U@      <@     �Q@       @      3@       @      3@     @Q@     �a@      .@      .@     �C@     �`@     �a@      @      4@      $@      D@      @      C@      &@      A@      �?      &@              @     �H@      U@       @      $@      1@      J@     �L@              $@       @      (@       @      <@      @      &@      �?      @              @      9@     �M@      �?      "@       @      4@      F@              @       @      @              *@      @       @              @              �?      3@     �H@      �?      @      @      *@      ?@              @      �?      @              @      @      @              @              �?       @      6@      �?               @      @      6@              @               @              @              @                                      &@      ;@              @      @       @      "@                      �?       @              .@       @      @      �?                      @      @      $@              @      �?      @      *@               @      �?      �?              &@       @                                      @      @      @               @              @      @                              �?              @              @      �?                               @      @               @      �?      @      @               @      �?                      $@      @      7@              @                      8@      9@      �?      �?      "@      @@      *@              @              @       @      @      @      2@              @                      *@      2@                      @      3@      @              �?               @               @       @      @              @                      "@      1@                      @      1@      @              �?                               @      �?      &@                                      @      �?                               @                                       @              @      @      @               @                      &@      @      �?      �?      @      *@      @              @              @       @       @      �?      �?               @                      $@      @      �?              @      @      @                              @              @       @      @                                      �?      @              �?       @      $@      �?              @               @       @      H@      1@      B@      @       @       @      .@      4@     �L@      *@      @      6@      T@     �U@      @      $@       @      <@      @      =@      (@      6@      @      @      @      $@      .@      I@      (@      @      0@     �N@      M@      @      @      @      .@       @      9@      (@      6@      @      @      @      "@      &@     �F@      (@      @      *@      L@     �C@       @       @      @      $@       @      (@      (@      3@       @       @      @      @      @      ?@      &@      @       @     �B@     �B@       @              @      @              *@              @      @      @              @      @      ,@      �?              @      3@       @               @              @       @      @                                              �?      @      @                      @      @      3@      @       @              @              @                                                               @                      @              @      @                      �?                                                              �?      @      @                              @      (@               @              @              3@      @      ,@       @       @      �?      @      @      @      �?              @      3@      <@      �?      @      @      *@      @      1@      @      $@       @       @              @      @      @      �?              @      3@      ;@      �?      @      @      (@      @      1@      @      @       @       @              @      @      @      �?              @      1@      6@      �?      @      @      &@       @                      @                              �?                                               @      @                              �?      �?       @              @                      �?                      @                      @              �?                              �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�xyhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmK}hnh4h7K ��h9��R�(KK}��hu�BX         >                    �?l�D���?�	           ��@                          �3@�n�X���?p           <�@                          �1@8�QR���?�           H�@                            @�7�<3��?�            �r@                           �?���J�?�             k@                           �?�q�q��?             H@������������������������       �T#G�h�?             7@������������������������       �+�����?             9@	       
                    @�y��y��?u             e@������������������������       �N��T>;�?L            @\@������������������������       ��cU��#�?)            �K@                           �?R���Q�?2             T@������������������������       �}��7�?             &@                           @��.����?+            @Q@������������������������       ��ˠT��?             F@������������������������       �a��+e�?             9@                            @�*9�b��?�            x@                            �?<�<�?�            �q@                           @vq��u�?}            �i@������������������������       ��Q2�?X            �b@������������������������       ��>u0i�?%            �L@                           �?c�����?2            �S@������������������������       �^p�F�?            �@@������������������������       �{�m<��?            �F@                           �?]19A~�?=            @Y@                           �?��V��?%            �O@������������������������       ���,d!�?             7@������������������������       �>
ףp=�?             D@                           �?Lt�<��?             C@������������������������       ���1G���?
             *@������������������������       ��������?             9@        /                    @�Π'f�?�           ��@!       (                   �7@����A��?�           ؄@"       %                    �?��H�T�?�            �t@#       $                   �6@\
t�?U            �a@������������������������       �P-����?<            �W@������������������������       ������j�?             H@&       '                   �4@$�&�k$�?y            �g@������������������������       ��K2���?            �G@������������������������       ��K�}
��?Z            �a@)       ,                    �?ð�E���?�            �t@*       +                     �?�-�)8D�?:            �W@������������������������       ��UbQ[F�?%            �J@������������������������       ��ܤ�?             E@-       .                   �9@yV4���?�             n@������������������������       ����&�?<             Y@������������������������       � 6�����?W            �a@0       7                   �6@li�c�z�?&           �|@1       4                   �5@����v�?�             n@2       3                     @_��4���?s            �f@������������������������       ��Zr_�?]            �b@������������������������       �����?             ?@5       6                    @�A�I��?%            �M@������������������������       �\���(\�?             D@������������������������       ����	"�?
             3@8       ;                    @*�o� �?�            @k@9       :                    @S�i�M�?P            @^@������������������������       ��������?             D@������������������������       �F��d&(�?5            @T@<       =                    @{�
;�?>            @X@������������������������       ��9����?             F@������������������������       ���1�P�?             �J@?       ^                    �?��H�	�?4           t�@@       O                    @�Ukt3m�?N           8�@A       H                    �?7�=��J�?s            �@B       E                     �?;�l�/�?�            �n@C       D                    �?���.{=�?+            �M@������������������������       ��9����?             6@������������������������       ���0\K5�?            �B@F       G                   �9@�(��?t            @g@������������������������       �mJ�Y ��?]            �b@������������������������       �'a����?             C@I       L                   �8@�\t�'<�?�            �t@J       K                    �?��{o�?�            �i@������������������������       �j�V���?            �@@������������������������       �#�,��.�?v            �e@M       N                    @     ^�?J             `@������������������������       ��paRC4�?'             Q@������������������������       �����2�?#             N@P       W                   �4@tfKS�?�            0v@Q       T                   �3@������?C             \@R       S                    @������?-             R@������������������������       �=�U����?             9@������������������������       ��{~���?            �G@U       V                    �?�Q����?             D@������������������������       �������?
             .@������������������������       �Ǻ����?             9@X       [                   �>@,I¢ʌ�?�            `n@Y       Z                   �;@D;���U�?�            `j@������������������������       ��
A(0�?q            @g@������������������������       �)\���(�?             9@\       ]                    @     ��?             @@������������������������       ��(\����?             $@������������������������       �1�~�4_�?             6@_       n                   �3@'�q���?�           L�@`       g                     �?��q�?�?           p|@a       d                     �?"ĕ�wF�?�            @o@b       c                    @��2�i]�?S            �`@������������������������       �x�R���?$            �M@������������������������       �į�JƓ�?/            �R@e       f                    @o�����?I             ]@������������������������       �c}h���?"             L@������������������������       �hE#߼�?'             N@h       k                   �0@/�b����?            �i@i       j                     @PR�5�`�?             ?@������������������������       ��n_Y�K�?             *@������������������������       ��^B{	��?             2@l       m                     @�8���?l            �e@������������������������       ��ܤ�[�?1             U@������������������������       ��N'�T�?;            �V@o       v                   �9@��2Z��?�           `�@p       s                    �?���6��?N           p�@q       r                   �6@�|�6��?`            `c@������������������������       ��S�v��?A            �Y@������������������������       �f|�We��?            �J@t       u                     �?4�5��?�            0w@������������������������       �>��;�T�?C            �Z@������������������������       ��Y}�l�?�            �p@w       z                     �?Q'37��?}            �g@x       y                    @��9"�?A            �X@������������������������       ���@^���?5            �S@������������������������       �q=
ףp�?             4@{       |                     @r��/���?<             W@������������������������       ��*�C��?             �I@������������������������       �tĖ��?            �D@�t�bh�h4h7K ��h9��R�(KK}KK��h��B8J        |@     �U@     �t@     �E@     �Q@      9@      T@     8�@     ��@      K@     @R@     �f@     P�@     �z@      0@     �S@      L@      \@     �O@     �k@     �B@     �\@       @      :@      @      <@     �t@     �t@      2@      =@     �J@     �r@     �h@      @      :@      4@     �B@      2@     �S@       @     �B@      �?                       @     �j@     �a@      @      @      0@     �Z@     �J@              @              "@      @      ?@              (@                              @     �[@     �P@      @               @      G@      .@                                              4@              @                              @     �W@     �H@                      @      :@      &@                                               @              @                                      5@      @                       @      @      @                                              @              @                                      @      @                       @      �?      �?                                               @              �?                                      ,@                                      @      @                                              (@               @                              @     �R@      G@                      @      6@      @                                              "@                                              @     �L@      =@                      �?      $@      @                                              @               @                                      1@      1@                       @      (@       @                                              &@              @                                      0@      1@      @              @      4@      @                                                                                                      @      �?      �?              @      �?                                                      &@              @                                      &@      0@       @                      3@      @                                               @              @                                      $@      @                              .@      �?                                              @              @                                      �?      "@       @                      @      @                                              H@       @      9@      �?                      @     �Y@     �R@      �?      @       @      N@      C@              @              "@      @      D@       @      2@      �?                              U@      M@      �?      @      @      D@      6@                              @       @     �@@       @      &@      �?                              K@      E@              @      @     �@@      2@                              @       @      1@       @      @      �?                              C@      C@               @      @      8@      .@                               @       @      0@              @                                      0@      @              �?              "@      @                              �?              @              @                                      >@      0@      �?               @      @      @                              @              @              @                                      ,@      $@                                                                      �?               @              @                                      0@      @      �?               @      @      @                              @               @              @                              @      3@      0@              �?       @      4@      0@              @               @      �?      �?                                              @      $@      *@                       @      ,@      (@              @               @      �?                                                              @      @                              @      @              @                              �?                                              @      @      @                       @       @      @              �?               @      �?      @              @                                      "@      @              �?              @      @              �?                              �?              @                                      �?                                      @      �?                                              @               @                                       @      @              �?              �?      @              �?                             �a@     �A@     @S@      @      :@      @      4@      ]@     @h@      ,@      9@     �B@     `h@     @b@      @      5@      4@      <@      .@      W@      9@     �L@      @      1@      @      *@     �A@     @W@       @      3@      :@     �]@     @U@      @      0@      0@      3@      *@     �L@      @      >@               @      @      @      7@     �H@      @      "@      1@     �O@      =@       @      @      �?      &@      @      :@      @      @              @      �?       @      @      =@      @      @      &@      8@      $@       @                      @      @      ,@       @      @              @      �?      �?      @      <@                      @      1@      @                              @      @      (@      @       @                              �?              �?      @      @       @      @      @       @                                      ?@       @      7@              @      @      �?      3@      4@              @      @     �C@      3@              @      �?       @              "@               @                                      @       @              �?      �?      @       @               @              @              6@       @      .@              @      @      �?      (@      (@              @      @      A@      1@              @      �?      @             �A@      2@      ;@      @      "@              $@      (@      F@       @      $@      "@     �K@      L@       @      $@      .@       @      @      @      @      @              �?                      @      7@       @      @              7@      &@              @      @      @      @       @      @      @              �?                       @      (@      �?      @              @       @              @       @      @      �?      �?               @                                      �?      &@      �?      �?              1@      @                      @               @      @@      .@      5@      @       @              $@      "@      5@              @      "@      @@     �F@       @      @      $@      @      @      @      �?      $@      @      �?               @      @      *@              �?      @      (@      ?@              @      @       @              9@      ,@      &@      @      @               @      @       @              @      @      4@      ,@       @      @      @      @      @     �H@      $@      4@      �?      "@              @     @T@     @Y@      @      @      &@     @S@     �N@              @      @      "@       @      ;@       @      @               @              @      F@     �Q@              @      @      D@      ;@                      @      @              8@       @      @               @              @      C@     �F@              @      @      ?@      0@                      �?       @              5@       @       @               @              @     �@@     �F@              @      @      5@      &@                                              @              @                                      @                                      $@      @                      �?       @              @                                                      @      9@                              "@      &@                      @       @              @                                                      @      (@                               @      "@                      @                                                                              �?      *@                              �?       @                               @              6@       @      *@      �?      @               @     �B@      ?@      @      @      @     �B@      A@              @              @       @      *@      @      $@              @               @      5@      7@      @      �?      @      ,@      (@              @              �?       @      @      �?      @              @               @      �?      @      �?               @      &@      @               @                      �?      "@      @      @              @                      4@      3@      @      �?      �?      @       @               @              �?      �?      "@      @      @      �?      �?                      0@       @       @       @       @      7@      6@              �?              @              @      �?       @              �?                      ,@      @                      �?      @      "@                              �?              @       @      �?      �?                               @      @       @       @      �?      0@      *@              �?              @             �l@      I@     �j@     �A@     �F@      4@      J@     �k@     �p@      B@      F@      `@     �s@     `l@      (@     �J@      B@     �R@     �F@     �X@     �@@     �Z@      2@      @@      .@      9@      I@      X@      *@      A@      R@     �]@     @Y@      @     �@@      5@      B@      ;@     @P@      5@     �I@      $@      9@      @      *@      C@     �S@       @      2@      C@     �S@      N@       @      4@      0@      5@      &@      B@       @      0@      @      *@      �?      @      4@      B@      @       @      *@      <@      6@              @      "@       @      @      "@              �?              @              �?      $@      @      �?       @      @       @      @                      �?       @              �?                               @              �?       @      @               @       @                                      �?       @               @              �?              �?                       @      @      �?              @       @      @                              @              ;@       @      .@      @      $@      �?      @      $@      =@      @      @       @      4@      3@              @       @              @      ;@       @      *@      �?      @      �?       @      $@      :@              @       @      *@      1@              @      @              @                       @      @      @               @              @      @       @              @       @              �?      @               @      =@      *@     �A@      @      (@      @       @      2@      E@      @      $@      9@      I@      C@       @      *@      @      *@      @      8@      "@      1@      @      @      �?      @      (@      A@       @       @      @      A@     �@@              @              "@              �?      �?      @              @               @               @              @       @      @      "@                              �?              7@       @      *@      @      @      �?      �?      (@      @@       @      @      @      ?@      8@              @               @              @      @      2@       @      @      @      @      @       @      �?       @      2@      0@      @       @      $@      @      @      @      �?      @       @      �?      @       @      @      @      @                      @      &@      @       @       @      @      @      �?      @      �?      $@      �?       @      @       @       @      @      �?       @      .@      @       @               @              �?      @     �@@      (@     �K@       @      @       @      (@      (@      2@      @      0@      A@     �D@     �D@      @      *@      @      .@      0@      *@              2@                                      @      (@       @      �?      .@      7@      (@                      �?      @      @      @              @                                      @      &@      �?      �?      "@      0@      $@                      �?      @      @      �?                                                               @      �?      �?       @       @       @                               @              @              @                                      @      "@                      �?       @       @                      �?       @      @       @              (@                                       @      �?      �?              @      @       @                                      �?       @               @                                              �?      �?              @      �?      �?                                      �?      @              $@                                       @                                      @      �?                                              4@      (@     �B@       @      @       @      (@      @      @      @      .@      3@      2@      =@      @      *@      @      &@      (@      4@      (@      @@      @      @      @      &@      @      @       @      .@      ,@      2@      =@      @      (@      �?      "@       @      0@      (@      @@      @      @      @      "@      @      @       @      (@      ,@      .@      :@      @       @      �?       @       @      @                      @      �?      �?       @                              @              @      @              @              �?                              @       @      @      @      �?                      �?              @                      �?      �?      @       @      @                                      @       @                                                                              �?       @               @                      @       @               @      �?                      �?              @                      �?              �?       @       @     @`@      1@     @[@      1@      *@      @      ;@     `e@     @e@      7@      $@     �L@     �h@     �_@      @      4@      .@     �C@      2@      H@      @      B@      @      �?              @     �Z@     �V@      @      �?      *@     �R@      F@              @      @       @      @     �A@      @       @       @                      @     �M@     �G@       @      �?       @      D@      5@              @      @      @      @      3@      �?      @       @                             �@@      ?@       @      �?      @      9@      "@                              @      �?      "@               @                                      .@      @              �?      �?      .@       @                                      �?      $@      �?      �?       @                              2@      8@       @              @      $@      �?                              @              0@      @      @                              @      :@      0@                      @      .@      (@              @      @      @      @      @      @      @                                      &@      *@                      �?      �?      @                      @      @      @      $@              �?                              @      .@      @                      @      ,@      @              @      @                      *@      �?      <@       @      �?               @     �G@     �E@      �?              @      A@      7@              @              �?      �?                                                              0@      @                               @       @                                                                                                       @                                              @                                                                                                       @      @                               @      @                                              *@      �?      <@       @      �?               @      ?@      C@      �?              @      @@      .@              @              �?      �?      @              1@              �?                      *@      5@      �?                      ,@      &@                              �?               @      �?      &@       @                       @      2@      1@                      @      2@      @              @                      �?     �T@      (@     @R@      *@      (@      @      6@     @P@      T@      4@      "@      F@      _@     �T@      @      ,@      "@      ?@      *@      R@      @      P@      &@      @      �?      .@     �K@      Q@      @      @      @@     �W@      F@      @      $@      @      2@      (@      6@              &@       @      �?      �?      @      8@      >@               @      @      ;@      0@              @               @      @       @              @       @      �?      �?      �?      4@      3@              �?      @      3@      (@              @                      @      ,@              @                              @      @      &@              �?               @      @               @               @              I@      @     �J@      "@      @              &@      ?@      C@      @      @      =@      Q@      <@      @      @      @      0@      @      "@              8@      @                      @      "@      "@       @      @      @      0@      @              @              @             �D@      @      =@      @      @              @      6@      =@       @       @      8@      J@      5@      @              @      "@      @      $@      @      "@       @       @      @      @      $@      (@      0@       @      (@      =@      C@       @      @      @      *@      �?       @      �?      @              @      �?       @      @              $@              @      5@      3@              @      @      @      �?       @      �?      @               @      �?              @              "@              @      4@      (@               @      @      @      �?                      �?              @               @      @              �?                      �?      @              �?                               @      @       @       @       @      @      @      @      (@      @       @      @       @      3@       @      �?              @              @      @       @       @              �?       @      �?      "@      @       @      @      @       @       @                       @               @      �?                       @       @      @       @      @      �?              @      @      &@              �?              @        �t�bub��     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�cwhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKqhnh4h7K ��h9��R�(KKq��hu�B�         <                     @u�`��?�	           ��@                            �?�ϕ�U�?�           ��@                          �5@ey��aj�?�           �@       	                   �0@piq�.�?�           ��@                           @(�B'�?-            �P@                           �?      �?!             H@������������������������       ���3L��?             ;@������������������������       ��3_<�?             5@������������������������       ��)O�?             2@
                           �?@��a!r�?T           ��@                           �?;Ocw���?|            �i@������������������������       ����\uR�?5            �U@������������������������       �y�*3��?G            @]@                           @	ڬre��?�            @t@������������������������       �
�:�1��?�            @r@������������������������       �     ��?             @@                           �?TVZ���?@           p~@                          �6@��Z`�E�?�            �g@                           @     ��?             @@������������������������       �ܶm۶m�?             ,@������������������������       ��n����?
             2@                           @�q�q�?k            �c@������������������������       �po���?O             ]@������������������������       �X�EQ]N�?            �E@                           @�n0E>��?�            �r@                           �?�W%�v��?�            Pp@������������������������       �ÞGi���?-            �R@������������������������       ��<+�?y            `g@                          �:@�j U��?            �A@������������������������       ��&%�ݒ�?             5@������������������������       ����S�r�?
             ,@        /                    �?��E��'�?           D�@!       (                    @�+69x�?�           ȉ@"       %                   �4@�Y}9p�?�            �t@#       $                     �?<��|L�?N            �`@������������������������       �t�Qe6�?7            �X@������������������������       ��E����?             B@&       '                    �?�x�_��?w            �h@������������������������       �c�_����?V            @b@������������������������       �F%u��?!             I@)       ,                    �?�[C�]�?2           �~@*       +                    �?��k��&�?�             j@������������������������       �7����?r             f@������������������������       ��~$7q�?             ?@-       .                     �?��N.-��?�            �q@������������������������       �>A�F<�?\             c@������������������������       �X��`k�?V            �`@0       7                    @NrHҬ�?           ��@1       4                    @���I���?�           h�@2       3                   �;@����Bu�?�            �@������������������������       �]�����?j           0�@������������������������       �D�95��?9            �V@5       6                     �?���,3��?K            @[@������������������������       �.��d��?.            @P@������������������������       ��9����?             F@8       ;                    @[h#&
i�?0            �R@9       :                    @��6�/�?(             O@������������������������       ��s-s��?             G@������������������������       �      �?	             0@������������������������       �������?             *@=       Z                   �7@۞���?�           ��@>       K                    �?ܕp(U��?�           H�@?       F                   �4@�m3 H��?�            �l@@       C                    �?h�����?e            `d@A       B                    @�G�z.�?2             T@������������������������       �'�z.���?"            �J@������������������������       ���h�C�?             ;@D       E                    @�3l��?3            �T@������������������������       �b�n`��?%             O@������������������������       �Z�eY�e�?             5@G       J                    �? \��M�?-             Q@H       I                   �5@     ��?             @@������������������������       �9��8���?             2@������������������������       �d}h���?	             ,@������������������������       ��Kh/���?             B@L       S                    @��Փ�M�?j           �@M       P                    �?�I�{VP�?$           �}@N       O                   �6@UUUUU5�?w             h@������������������������       �D�����?j             e@������������������������       ��������?             8@Q       R                    @���JMn�?�            �q@������������������������       ���/5��?P            �_@������������������������       �\37U[v�?]            �c@T       W                    �?��� =�?F            �Y@U       V                    @p��G��?             �E@������������������������       �r�q��?             B@������������������������       �����>4�?             @X       Y                   �1@��x�5�?&            �M@������������������������       �j�V���?             &@������������������������       ���8��x�?             H@[       d                    �?'첃%[�?�            `u@\       c                   �>@�\�dD\�?Q            �\@]       `                    @�����?G            @X@^       _                    @������?,            �L@������������������������       ���(\���?              D@������������������������       �4%���?             1@a       b                    @�(\����?             D@������������������������       �������?             ;@������������������������       �3�E��?             *@������������������������       ��ѳ�w�?
             1@e       l                   �=@�!����?�            �l@f       i                   �8@ Ս����?f            @d@g       h                    @�M7�o��?#            �M@������������������������       ��ۚ�R�?             G@������������������������       ��θ�?             *@j       k                   �9@�d�M��?C            �Y@������������������������       ��?�߾�?             9@������������������������       �\��[���?2            �S@m       p                    @�;�JBf�?"            �P@n       o                    �?�q�MU�?            �J@������������������������       ��j">���?            �D@������������������������       �9��8���?             (@������������������������       ��s�n_�?             *@�t�bh�h4h7K ��h9��R�(KKqKK��h��BC       ~@     �S@     �u@     �B@     �U@      9@     @W@     �@     �@      N@     @V@     `d@     Ђ@     {@      .@     �O@     �K@     �]@      H@     `v@     �F@     �m@      0@     �G@      @     �M@     @{@     |@      F@      O@      Z@     �z@     pq@      @     �K@     �@@     �R@      9@     �^@      &@      Y@      "@      *@      @     �@@     @]@      g@      .@      7@      I@     �g@     �^@      �?      A@      &@      @@      "@     �R@      @     �C@      @      �?      �?      $@      Z@     �`@      @      "@      :@     @^@      D@              $@              "@      @      @              �?                                      8@      =@                              @      �?                                              @              �?                                      5@      .@                              @      �?                                              �?              �?                                      ,@      &@                                                                                      @                                                      @      @                              @      �?                                              �?                                                      @      ,@                                                                                     �P@      @      C@      @      �?      �?      $@      T@     @Z@      @      "@      :@     @]@     �C@              $@              "@      @      A@       @      7@      @                      @      2@      9@       @      @      0@      I@      .@              �?              @      @      0@       @      @                                      ,@       @              @      @      ;@      @              �?                      �?      2@              4@      @                      @      @      1@       @      �?      "@      7@      $@                              @       @     �@@      @      .@       @      �?      �?      @      O@      T@      �?      @      $@     �P@      8@              "@              @              7@      @      &@       @      �?      �?      @      L@      S@      �?      @       @      O@      8@              "@              @              $@              @                                      @      @                       @      @                                      �?              H@      @     �N@      @      (@      @      7@      *@     �I@      (@      ,@      8@     @Q@     �T@      �?      8@      &@      7@      @      ;@      @      3@      �?      @               @      @     �A@      @      @      @      :@      ?@              @       @      "@      @      @      �?       @              @                              *@                      �?      @       @                                               @      �?       @              @                               @                      �?      �?       @                                              @                                                              &@                              @                                                      6@      @      1@      �?                       @      @      6@      @      @      @      5@      =@              @       @      "@      @      0@      @      .@      �?                       @      �?      2@              @       @      ,@      .@              @       @       @      @      @               @                                      @      @      @              @      @      ,@                              �?              5@       @      E@      @      "@      @      .@      "@      0@      "@      $@      2@     �E@     �I@      �?      2@      "@      ,@      @      5@       @     �D@              "@      @      (@      @      *@      "@      $@      0@      D@      G@      �?      0@      @      "@      @      @              .@               @              �?      �?      @      @      �?       @      4@      ,@      �?      @              @              1@       @      :@              @      @      &@      @      "@      @      "@      ,@      4@      @@              *@      @      @      @                      �?      @                      @      @      @                       @      @      @               @      @      @                                      @                      �?      @      @                      �?       @       @               @               @                              �?                               @                                      �?      �?      @                      @      @             �m@      A@      a@      @      A@       @      :@     �s@     �p@      =@     �C@      K@      n@     �c@       @      5@      6@      E@      0@     @^@      0@      P@       @      *@               @     @g@     �b@      @      5@      2@     �\@     �S@              @      @      (@      @      J@      &@     �C@              "@              @      F@      H@       @      "@      (@     �E@      B@              @      @       @      @      7@              @              @              @     �@@     �@@                       @      2@      *@                              @              3@                              @              @      6@      8@                      �?      .@      $@                              �?              @              @                                      &@      "@                      �?      @      @                               @              =@      &@      B@              @               @      &@      .@       @      "@      $@      9@      7@              @      @      @      @      2@       @      8@              @               @       @       @      �?      "@      $@      4@      2@              @      @      @      @      &@      @      (@               @                      @      @      �?                      @      @              �?                             @Q@      @      9@       @      @              @     �a@     @Y@      @      (@      @      R@      E@                       @      @      �?      B@       @      "@                               @      S@      A@              @      @      5@      6@                                              :@       @      "@                               @     @Q@      @@              @      @      3@      (@                                              $@                                                      @       @                               @      $@                                             �@@      @      0@       @      @              �?     �P@     �P@      @      "@      @     �I@      4@                       @      @      �?      6@              @       @                      �?      8@      G@      @      @       @      =@      @                       @      �?      �?      &@      @      "@              @                      E@      5@      �?      @      �?      6@      ,@                              @             �\@      2@     @R@      @      5@       @      2@     �`@     �\@      7@      2@      B@     @_@     �S@       @      ,@      1@      >@      (@     �[@      2@     �N@      @      3@       @      $@     @`@     �Z@      5@      2@     �@@     @]@     @P@       @      *@      .@      9@      (@     @T@      1@     �J@      @      ,@       @       @     �^@     �V@      2@      1@      >@     @[@      J@       @      &@      *@      2@      $@     �S@      ,@     �G@       @      @              @     �^@     �T@      "@      (@      5@      Z@     �H@               @       @      (@      @       @      @      @       @      "@       @       @              @      "@      @      "@      @      @       @      @      &@      @      @      =@      �?       @              @               @      @      0@      @      �?      @       @      *@               @       @      @       @      *@              �?              @               @      @      .@       @      �?      @      @       @              �?       @      @              0@      �?      @              �?                       @      �?      �?                      @      @              �?              @       @      @              (@      �?       @               @      @      "@       @              @       @      ,@              �?       @      @              @               @      �?       @               @      @      @       @              @      @      ,@              �?       @      �?              @              @              �?              @      @      @                      @      @      &@              �?       @      �?              �?               @      �?      �?              @                       @                       @      @                                              �?              @                                              @                              �?                                      @             �^@      A@      [@      5@      D@      3@      A@     @Z@     @`@      0@      ;@     �M@     �e@     @c@      (@       @      6@      F@      7@     �Y@      0@      T@       @      4@      "@      *@     @Z@     @Y@      &@      2@     �C@     �a@     �V@       @      @      @     �@@      @      G@      @      5@      @      @      @      @      =@      =@      @      @      @      7@      4@      �?      @      @      *@      @     �C@      @      2@      @      @       @      @      ;@      5@      �?      @      @      ,@      &@              �?      �?       @              1@              @               @       @              2@      $@      �?                      @      &@                              @              0@                               @       @              @      @      �?                      @      @                              @              �?              @                                      &@      @                                      @                                              6@      @      (@      @       @              @      "@      &@              @      @      @                      �?      �?       @              4@      @      @               @                      @      &@              @      @      @                      �?      �?       @               @              @      @                      @      @                                       @                                                      @      @      @              @      @               @       @      @              @      "@      "@      �?       @       @      @      @      @              �?               @                       @      �?                              @       @      �?      �?               @      �?                                                               @      �?                              @      @              �?               @      �?      @              �?               @                                                                      @      �?                                              @       @              �?      @                      @      @              @      @      �?              �?       @      @       @     �L@      "@     �M@      @      *@      @      $@      S@      R@      @      .@     �@@     @]@     �Q@      �?      @      @      4@      @     �F@       @     �I@      @      $@      @       @     �H@     @P@      @      &@     �@@     �X@     �M@              @      @      .@      @      .@              ,@              �?      �?      �?      A@      D@               @      3@      E@      *@               @      �?      @      �?      (@              *@                      �?      �?      ;@      A@               @      *@      E@      *@               @      �?      @      �?      @              �?              �?                      @      @                      @                                                              >@       @     �B@      @      "@       @      @      .@      9@      @      "@      ,@      L@      G@              �?      @      "@      @      (@      @      .@      @       @      �?              "@      1@       @      @      @      ?@      0@              �?              @              2@      @      6@       @      @      �?      @      @       @      @      @      &@      9@      >@                      @      @      @      (@      �?       @              @               @      ;@      @      �?      @              3@      (@      �?                      @              @              @                               @      *@      @      �?      @              @      @                              �?              @               @                                      *@       @      �?      @              @      @                              �?                              �?                               @              �?                              @                                                       @      �?      @              @                      ,@      @                              (@      @      �?                      @                                                                       @       @                              �?                                                       @      �?      @              @                      @       @                              &@      @      �?                      @              4@      2@      <@      *@      4@      $@      5@              =@      @      "@      4@      @@     �O@      $@       @      .@      &@      0@      @      @      $@      @      "@              "@              *@       @      @      @      0@      (@      �?       @       @       @      @      @      @      $@      @      @              @              *@       @      @      @      0@      $@               @      @       @      @       @       @       @      �?      @                              "@       @      @      @      @      @               @       @       @      @       @       @      @      �?      @                              @       @      �?      @      @      @               @               @                              @                                              @               @                       @                       @              @      �?      @       @       @                      @              @                      @      "@      @                      @               @               @      �?       @                      @              @                       @      @      �?                       @               @      �?      �?      �?                              �?                                      �?      @       @                       @                      @                              @               @                                                       @      �?               @              �?      ,@      *@      2@      $@      &@      $@      (@              0@      @      @      *@      0@     �I@      "@              @      "@      $@      ,@      @      (@      @      @      �?      (@              (@               @       @      0@     �H@      @              @      @      @       @      @      @              �?              @              @               @       @      @      :@      @                      �?               @      �?      @              �?               @              @                       @      �?      :@      @                      �?              @       @                                      �?                               @               @                                                      @      @       @      @      @      �?      "@              "@                      @      *@      7@      �?              @      @      @       @       @       @       @       @              �?              @                       @      @      �?                      �?                      @       @      @       @      @      �?       @              @                      @       @      6@      �?               @      @      @              @      @      @      @      "@                      @      @      @      @               @      @              @       @      @              @      @       @      @       @                      @      @      @       @               @      @              @              @               @      @       @      @      @                      @       @      @                      �?      @              @              @              @                              @                      �?      �?               @              �?                                                                      @       @      �?                                              @                      �?                       @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJn�i0hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKmhnh4h7K ��h9��R�(KKm��hu�B�         :                    �?9�HB��?�	           ��@                           �?�!���?           �@                           �?�ũ���?p           @�@                          �4@    �	�?�             p@                          �1@�]�"�?T            �_@                            �?�]�"R�?            �C@������������������������       ���!pc�?             &@������������������������       ��Cc}h�?             <@	       
                   �3@ˠT�x?�?:             V@������������������������       � ��9�?'             M@������������������������       �N<+	��?             >@                           @��e Ʊ�?M             `@                          �6@������?D            �[@������������������������       �<ݚ)�?             B@������������������������       ��H
����?.            �R@������������������������       �窷uJ��?	             3@                          �<@���D|��?�            �t@                            �?��au�?�            Pr@                          �2@^HT`!��?b            @c@������������������������       �����>4�?             <@������������������������       �Y�'��+�?O            �_@                            @��H���?W            `a@������������������������       ���QN�?             ?@������������������������       ��Ju�?F             [@                          �?@�0J5y�?            �A@                            �?��6��?             9@������������������������       �     ��?
             0@������������������������       �0�����?             "@������������������������       ��(\����?             $@       +                    �?hT���?�           ��@       $                    �?�Ϯ�_�?�            �q@        !                   �1@����"�?S            �`@������������������������       ��q-�?             *@"       #                     �?#Jp
���?M            @^@������������������������       �*Yp����?)            �N@������������������������       ��Y�H�7�?$             N@%       (                     @?�:��D�?g            �b@&       '                     �?���@^��?7            �S@������������������������       �j���� �?0             Q@������������������������       ��G�z��?             $@)       *                   �:@;�1����?0            @R@������������������������       �8��1��?)            �N@������������������������       �VUUUUU�?             (@,       3                   �6@6�z':�?�           �@-       0                   �4@VN�x�?�            pw@.       /                    �?Ƶ逕�?�            �m@������������������������       ��h$���?
             .@������������������������       �^t�D.��?�            �k@1       2                    @�k��]�?S             a@������������������������       �4'���a�?J            @^@������������������������       �      �?	             0@4       7                    �?���e�?�            �v@5       6                   �;@�1H1�?P             _@������������������������       ��p=
�#�?5             T@������������������������       ��A�0�~�?             F@8       9                     �?$����=�?�            �m@������������������������       ���1�>�?M            �]@������������������������       �	���ĳ�?L             ^@;       N                    �?�������?�           �@<       E                     @�q����?�           ܑ@=       D                    @x><]��?J           `�@>       A                     �?�s�G��?A           ��@?       @                    @n�2�?�           ��@������������������������       ��t����?A           p@������������������������       ���ݷl�?_             c@B       C                    �?�k����?�            �p@������������������������       ���o��?G            �]@������������������������       �,"���?Z            �b@������������������������       �      �?	             0@F       M                    @Vzk��l�?            `i@G       J                    @�Z�/?�?w             h@H       I                   �1@R�i\�:�?             �K@������������������������       �REQE�?
             5@������������������������       ��������?             A@K       L                    @�&^Ň�?W            @a@������������������������       ��k�n�?4            @U@������������������������       � �T`��?#            �J@������������������������       ��������?             $@O       ^                    @v���_L�?�           ,�@P       W                     @67,�?"           ��@Q       T                   �4@��S����?�           ��@R       S                     �?C%��NM�?�             w@������������������������       �-րR��?�            �p@������������������������       ��
�J�u�?>            �Y@U       V                   �:@dK.[C��?�            Pt@������������������������       ������?�             n@������������������������       �M�4M�4�?4             U@X       [                   �4@UUUUUa�?w             h@Y       Z                    @�<"H��?D            @[@������������������������       �R����?            �@@������������������������       �90\�Uo�?/             S@\       ]                   �=@�����?3            �T@������������������������       �B��Q,�?-            �R@������������������������       �B{	�%��?             "@_       f                     @3pLo��?�            `q@`       c                    �?K8�_��?|             i@a       b                   �2@�z��R�?*            �Q@������������������������       �B{	�%��?             2@������������������������       �������?"             J@d       e                     �?M���_��?R            ``@������������������������       �AM�h���?@             Z@������������������������       �v�Ë���?             ;@g       j                   �8@]��{�W�?.            @S@h       i                    @IPS!���?             J@������������������������       �z�}wi��?            �B@������������������������       �hE#߼�?             .@k       l                   �:@�
F%u�?             9@������������������������       �      �?              @������������������������       �{�/��>�?	             1@�t�bh�h4h7K ��h9��R�(KKmKK��h��B�@       �}@     �U@     �s@      9@      Q@      ;@      V@     ��@     H�@     @R@     �V@     �c@     H�@     }@      *@     �H@     �E@      ]@      K@     �j@     �D@     �a@      .@      F@      5@      F@     �V@     �i@     �C@     �I@      U@      l@     @k@      $@      8@      @@     �P@      D@      W@      (@     �E@              1@      �?      ,@     �F@      W@      3@      2@      4@      X@     �K@               @      $@      8@      2@     �B@      @      2@              @      �?      @      >@     �K@      @      "@      @     �D@      6@              @      �?      @      "@      5@              @              �?                      :@     �@@      @      �?      @      :@      @              �?               @              $@               @                                      "@      *@      �?              �?      @                                                      @                                                      @       @                                                                                      @               @                                      @      &@      �?              �?      @                                                      &@              �?              �?                      1@      4@      @      �?       @      7@      @              �?               @              "@              �?                                      "@      (@      @      �?       @      (@      @              �?               @               @                              �?                       @       @                              &@                                                      0@      @      .@               @      �?      @      @      6@       @       @       @      .@      1@              @      �?       @      "@      $@      @      .@               @      �?      @      @      6@       @       @       @      $@      .@              @      �?       @      @                      @                              @      @      @              �?      �?      @      "@               @              �?              $@      @       @               @      �?                      3@       @      @      �?      @      @              �?      �?      �?      @      @                                               @      �?                                      @       @                                      @     �K@       @      9@              ,@               @      .@     �B@      (@      "@      .@     �K@     �@@              @      "@      4@      "@     �J@      @      7@              $@               @      ,@     �A@      (@      @      "@     �J@     �@@              @       @      1@      "@      <@       @      $@              @               @      @      7@      @      �?      @      B@      6@              @      �?      @      @      @              @                                       @      "@       @              @      @                                      �?              9@       @      @              @               @       @      ,@      @      �?      �?      ?@      6@              @      �?      @      @      9@       @      *@              @                      $@      (@      @      @      @      1@      &@              �?      @      (@      @      @              @                                      @      @              �?       @       @      @                               @              3@       @      @              @                      @      "@      @      @      @      .@       @              �?      @      $@      @       @      @       @              @              @      �?       @               @      @       @                              �?      @                      @       @               @              @      �?       @                      @       @                              �?       @                       @                      �?              @               @                      @                                               @                       @       @              �?                      �?                                       @                              �?                       @                               @                                               @      @                                              �?             @^@      =@      Y@      .@      ;@      4@      >@     �F@     �\@      4@     �@@      P@      `@     `d@      $@      0@      6@     �E@      6@     �L@      @      =@      @      $@       @      @      1@     �@@      @      @      "@      C@      E@      @      �?       @      ,@      @      ;@       @      *@       @      @              @       @      (@              @      �?      8@      1@      @      �?              &@              �?                                                      @                                      �?      @                                              :@       @      *@       @      @              @       @      (@              @      �?      7@      (@      @      �?              &@              $@      �?       @       @      @              @       @      @               @      �?      0@       @                              @              0@      �?      @               @                              @               @              @      $@      @      �?               @              >@       @      0@       @      @       @       @      "@      5@      @      �?       @      ,@      9@                       @      @      @      5@              @                               @      @      "@      @              @      @      2@                      �?       @              2@              @                               @      @      @      @              @      @      .@                      �?       @              @                                                               @                       @              @                                              "@       @      "@       @      @       @              @      (@      �?      �?      @      "@      @                      �?      �?      @      "@       @      "@       @      @       @              @      &@      �?      �?      @      @      @                              �?      �?                                      �?                              �?                              @                              �?              @      P@      9@     �Q@      &@      1@      2@      8@      <@     �T@      .@      <@     �K@     �V@     @^@      @      .@      4@      =@      2@     �H@      $@      >@      @       @       @      @      9@      J@       @      ,@      *@      O@     �O@              @      @      4@      @      =@       @      7@      �?                      �?      6@     �C@      @      "@      "@     �G@      ?@              @              ,@      @                                                      �?               @              @      �?      �?      @                                              =@       @      7@      �?                              6@     �B@      @      @       @      G@      ;@              @              ,@      @      4@       @      @       @       @       @       @      @      *@      @      @      @      .@      @@                      @      @       @      4@       @      @       @       @      @       @      @      @      @      @      @      .@      ;@                      @      @       @                      �?                       @                      @                      �?              @                                              .@      .@     �D@       @      .@      $@      5@      @      >@      @      ,@      E@      <@      M@      @      $@      1@      "@      *@      @      @      2@              "@              (@      �?      (@              @      &@      0@      *@      �?       @      $@       @      @      �?      @      &@              �?              "@      �?      (@              �?      "@      *@      "@              �?      "@                      @              @               @              @                               @       @      @      @      �?      �?      �?       @      @      "@      (@      7@       @      @      $@      "@       @      2@      @      &@      ?@      (@     �F@      @       @      @      @       @      @      @      .@      @      @       @      @       @      @      @      @      1@      $@      2@              @      @      @      @      @      @       @      @      @       @      @              .@       @      @      ,@       @      ;@      @      �?      @      @      @     Pp@      G@     �e@      $@      8@      @      F@     �{@     �{@      A@      D@     @R@     �v@     �n@      @      9@      &@     �H@      ,@      b@      1@     �Q@       @       @              *@     �q@     `l@      0@      4@      <@     �f@     @Y@              @      @      4@      @     �]@      (@     �J@      �?       @              &@     `n@      i@      ,@      0@      :@     �`@     �T@              @       @      *@       @     �]@      (@     �I@      �?       @              &@      n@     �h@       @      0@      :@     �`@     �T@              @              *@       @      W@      @     �B@      �?      @              &@      c@     �a@      @      .@      5@     @W@      P@              @              (@       @     �O@      @     �@@      �?      @              &@     @^@      ]@      �?      @      *@      R@     �F@               @              $@      �?      =@              @                                      ?@      8@      @       @       @      5@      3@               @               @      �?      :@      "@      ,@              @                      V@     �M@      @      �?      @      D@      2@                              �?              (@       @       @               @                     �C@      A@              �?      @      &@      @                                              ,@      �?      (@               @                     �H@      9@      @                      =@      *@                              �?                               @                                      @      �?      @                      �?                      �?       @                      ;@      @      1@      �?                       @     �B@      ;@       @      @       @      H@      3@               @      �?      @       @      ;@      @      0@      �?                             �B@      ;@       @      @      �?      H@      0@               @      �?      @       @      &@      �?       @      �?                              @      @                              9@      @                                              @                                                              @                              *@                                                       @      �?       @      �?                              @      �?                              (@      @                                              0@       @      ,@                                      @@      5@       @      @      �?      7@      (@               @      �?      @       @      *@              "@                                      :@      ,@               @              $@      @              �?      �?      @       @      @       @      @                                      @      @       @       @      �?      *@      "@              �?               @                       @      �?                               @                                      �?              @                              �?              ]@      =@     �Y@       @      0@      @      ?@     `d@     �j@      2@      4@     �F@     `f@     @b@      @      2@       @      =@      $@      W@      5@     �Q@      @      &@      @      3@      b@     @f@      ,@      2@      @@     �`@     @Y@       @      @      @      6@      @     @R@      *@      L@      @       @      @      &@     �_@      b@      *@      ,@      3@     @Y@     �R@      �?      @      @      0@      @      E@              8@      �?      �?              @     �Y@     @V@      @      @      @     �H@      >@              �?      �?      @      @     �C@              1@      �?                       @     �N@     �M@       @      @      @      B@      :@              �?      �?       @      @      @              @              �?              �?     �D@      >@       @                      *@      @                              �?              ?@      *@      @@       @      @      @       @      8@      L@      "@       @      (@      J@     �F@      �?      @       @      *@              ;@      "@      8@      �?       @       @      @      8@     �I@      �?      @      @     �D@      @@      �?      �?              "@              @      @       @      �?      @       @      �?              @       @      @      @      &@      *@              @       @      @              3@       @      ,@       @      @               @      2@     �@@      �?      @      *@      A@      :@      �?                      @       @      @      @      *@               @              @      ,@      0@              @      (@      ;@      @                                              �?       @      �?              �?               @      @       @               @              ,@      @                                              @       @      (@              �?              �?      &@      ,@               @      (@      *@       @                                              (@      @      �?       @      �?              @      @      1@      �?              �?      @      3@      �?                      @       @      (@      @      �?       @                      @      �?      1@                      �?      @      0@                              @       @                                      �?                      @              �?                              @      �?                                      8@       @     �@@      @      @       @      (@      3@     �B@      @       @      *@      F@     �F@      �?      &@      @      @      @      3@      @      =@      @       @              @      0@      2@      @       @      (@      =@      @@              $@      @      @      @      $@       @      @      �?                      @      @      @       @               @      $@      4@              @      �?      �?              @      �?                                      �?                                              @      @                              �?              @      �?      @      �?                       @      @      @       @               @      @      ,@              @      �?                      "@      @      6@       @       @              @      *@      .@       @       @      $@      3@      (@              @      @      @      @      @      @      .@       @      �?              @      &@      $@       @       @       @      3@      @              @      @      @      @      @      �?      @              �?                       @      @                       @              @                              �?              @       @      @              @       @      @      @      3@                      �?      .@      *@      �?      �?      �?      �?              @      �?      @               @                      @      2@                              "@      @      �?      �?              �?              @              @                                      @      2@                              @      @                                               @      �?                       @                                                              @      @      �?      �?              �?                      �?                      �?       @      @              �?                      �?      @      @                      �?                                                      �?              @                                              �?      �?                      �?                              �?                               @       @              �?                      �?      @      @                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ*�aEhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKshnh4h7K ��h9��R�(KKs��hu�B(         :                    @,����?�	           ��@                          �4@m����?�           \�@                          �0@m/����?6           ��@       	                    @���X�??             \@                            �?�~_�{��?(            @Q@                           �?\")�i��?             G@������������������������       �����X�?             <@������������������������       �x�5?,R�?             2@������������������������       ���x�(��?             7@
                           �?l��i�?            �E@������������������������       ��������?
             1@                            �?��Q�}e�?             :@������������������������       �                     .@������������������������       ���!pc�?             &@                            @A��G��?�           8�@                            �?b�	�O��?           �z@                          �1@��vH��?�            `k@������������������������       ���c����?"             J@������������������������       � �gXq�?o            �d@                           �?H�et��?�            `j@������������������������       �܋;�J�?E            �Y@������������������������       �z��$9�?E            @[@                           �?"��w	��?�            �u@                           �?�h^���?I            @\@������������������������       �)栤�?%             O@������������������������       �仓kC�?$            �I@                           �?�;\�?�             m@������������������������       ��tP���?}            �h@������������������������       ��]1�[��?            �@@       -                    �?D�u�u�?P           ܔ@       &                    �?�����7�?!           P|@        #                    �?����?d�?�            �j@!       "                   �7@�Y]�S�?c            @c@������������������������       �����.�?,            �Q@������������������������       ��py�[��?7            �T@$       %                     @�L�@��?%             M@������������������������       ���w�AV�?            �E@������������������������       �������?	             .@'       *                     �?x���?�             n@(       )                    �?�$�4��?P            �]@������������������������       ���8����?@             X@������������������������       �&ޏ���?             6@+       ,                    �?�c��M�?I            �^@������������������������       ��A͈\w�?:            @X@������������������������       �ƵHPS!�?             :@.       5                   �?@R0\}x�?/           ��@/       2                    �?EB�-�H�?�           ��@0       1                   �5@    ���?�             p@������������������������       ��q�q�?             8@������������������������       ������?�             m@3       4                    �?j3�a�Z�?d           ��@������������������������       ����n�?�            �i@������������������������       ����7�R�?�            �t@6       9                     @0�w¹��?0             U@7       8                    �?����S�?             L@������������������������       �3�E��?             *@������������������������       ��s���?            �E@������������������������       �����S�?             <@;       T                    �?�Ns�H��?<           l�@<       E                   �0@������?           ��@=       >                     �?BR�8	�?.             S@������������������������       ��q�q�?	             2@?       B                    �?�CE5��?%             M@@       A                    @�����?             7@������������������������       ��z�G��?             $@������������������������       ��T�6|��?	             *@C       D                    @F����?            �A@������������������������       ��������?	             (@������������������������       �'�%����?             7@F       M                    @}T����?�           P�@G       J                    @�+Fi��?v             g@H       I                   �1@�������?J            @]@������������������������       �ffffff�?             4@������������������������       ��^�X�?=            @X@K       L                    @�ӫ����?,            �P@������������������������       �      �?             8@������������������������       �.T�J��?            �E@N       Q                     �?�����?t           ��@O       P                    @���ko�?_            �c@������������������������       �~X�<��?-             R@������������������������       �~VC�1��?2             U@R       S                    @��6��P�?           `{@������������������������       ��Uu�3�?�            �o@������������������������       ���<C�l�?t             g@U       d                    @-��� .�?$           (�@V       ]                    @����?V           x�@W       Z                   �2@Gb�4���?�            �k@X       Y                    @���c��?'            �P@������������������������       �h�����?             L@������������������������       ��9����?             &@[       \                     �?�.�U��?`            `c@������������������������       �     ��?2             T@������������������������       �R���ȿ�?.            �R@^       a                    �?_��^��?�            s@_       `                     @"1gE<�?P             ]@������������������������       �3=G�4��?J            �Z@������������������������       ��n���?             "@b       c                     @�i��X�?            �g@������������������������       �I��-X�?p            �d@������������������������       ���ճC��?             6@e       l                   �5@=�(���?�            `s@f       i                     �?�ڀ���?j             d@g       h                   �4@�(�Tw��?            �C@������������������������       ��j��p�?             ?@������������������������       �      �?              @j       k                    @N��IP��?N            �^@������������������������       �ݚ)�?0             R@������������������������       ���n���?             I@m       p                     �?d��R��?d            �b@n       o                    @������?             C@������������������������       �     ��?             0@������������������������       �.�袋.�?             6@q       r                    �?�[�	O��?J            �[@������������������������       �`�;��K�?             C@������������������������       �߉��`w�?3            @R@�t�bh�h4h7K ��h9��R�(KKsKK��h��BHD       �z@      T@     0t@     �C@      U@      ?@     @V@     ��@     0�@     �N@      U@      e@     ��@     �z@      &@      R@     �F@     �`@      M@     �p@     �G@     �i@      =@     �P@      :@     �N@     �g@     0r@      C@     �O@     @\@     �t@     �o@      @      J@      B@     @Y@     �G@      a@      $@     �J@      @      @              @     @`@      d@      "@      .@      A@     �d@     �U@              &@      @     �C@      (@      ,@      @      @                                      =@     �E@                              (@      @                                              *@      @       @                                      7@      .@                              $@       @                                              @               @                                      1@      *@                              @       @                                              @               @                                      "@      &@                                                                                      �?                                                       @       @                              @       @                                              @      @                                              @       @                              @                                                      �?              @                                      @      <@                               @      @                                              �?              @                                      @      @                                      �?                                                                                                      �?      5@                               @       @                                                                                                              .@                                                                                                                                              �?      @                               @       @                                             �^@      @      H@      @      @              @     @Y@     �]@      "@      .@      A@     `c@     @T@              &@      @     �C@      (@     �R@       @      =@      @      @              @     �R@     �Q@      @      @      ;@      R@      ?@              @       @      (@      $@     �C@       @      $@      @                       @     �C@      9@      @      @      1@     �F@      ,@               @              @      @      @                                                      5@      @                      @      *@      @                                       @      A@       @      $@      @                       @      2@      6@      @      @      (@      @@      &@               @              @      @     �A@              3@              @               @     �A@      G@       @      �?      $@      ;@      1@              @       @      @      @      .@              @                                      8@      9@              �?      @      3@      @                              @      @      4@              .@              @               @      &@      5@       @              @       @      (@              @       @       @      �?     �H@      @      3@       @      @              @      ;@     �G@      @      $@      @     �T@      I@              @      �?      ;@       @      8@              @              @                      $@      &@              @       @      5@      .@              @              &@              (@                              �?                       @      @                              &@      "@              @              &@              (@              @              @                       @      @              @       @      $@      @                                              9@      @      *@       @                      @      1@      B@      @      @      @      O@     �A@              @      �?      0@       @      4@      @      *@       @                      @      .@      =@      @      @      @     �H@      >@              @      �?      0@       @      @                                                       @      @              �?              *@      @                                              `@     �B@     @c@      7@      N@      :@      K@      M@     @`@      =@      H@     �S@     �d@     �d@      @     �D@     �@@      O@     �A@      K@      2@      F@      @      2@      "@      &@      ,@     �P@      1@      &@      3@     �L@      J@      @      $@      $@      6@      (@     �A@      &@      :@      @      @              @       @      D@       @      @       @      8@      8@      @      @      �?      @      �?      ?@      @      7@      @      @              @      @      6@      �?      @       @      0@      1@      @      @      �?      @      �?      .@              0@              @              �?      @      (@              �?       @       @      @      @                      �?              0@      @      @      @                      @              $@      �?      @               @      &@              @      �?      @      �?      @      @      @                                      @      2@      �?              @       @      @               @                               @      @      @                                      @      1@      �?              @      @       @              �?                               @      �?                                              �?      �?                              @      @              �?                              3@      @      2@       @      .@      "@      @      @      :@      .@      @      &@     �@@      <@      �?      @      "@      0@      &@      (@       @      ,@               @      @      @      @       @      @      @       @      5@      *@      �?      @      @      "@      @      "@      �?      (@               @      @      @      @      @      @      @       @      1@      (@      �?      �?              "@      @      @      �?       @                              �?              �?      @                      @      �?               @      @                      @      @      @       @      *@      @              @      2@       @      �?      "@      (@      .@              �?      @      @       @      @      @      @       @      $@      @              @      *@      @      �?      "@      &@      @              �?      @      @      @       @                              @                              @       @                      �?       @                              @      �?     �R@      3@     �[@      2@      E@      1@     �E@      F@      P@      (@     �B@      N@     �Z@     �\@      @      ?@      7@      D@      7@     �Q@      3@     �Y@      .@      B@      *@      E@      F@     �O@       @      A@     �D@     @Z@      \@              :@      *@      A@      4@      =@      @      ;@              *@      �?      "@      6@      9@      �?      @      "@     �H@      >@              $@      �?      $@      "@      @                                              @      �?      @              �?       @       @      �?              @              @              9@      @      ;@              *@      �?      @      5@      6@      �?      @      @     �G@      =@              @      �?      @      "@      E@      .@     �R@      .@      7@      (@     �@@      6@      C@      @      ;@      @@      L@     �T@              0@      (@      8@      &@      3@      @      B@      @      (@       @      $@      .@      0@              @      &@      9@      9@               @       @      @       @      7@      "@     �C@      &@      &@      $@      7@      @      6@      @      7@      5@      ?@     �L@              ,@      @      4@      @      @               @      @      @      @      �?              �?      @      @      3@       @       @      @      @      $@      @      @       @              @       @      @       @      �?              �?      @      @      2@       @                      �?      @      @       @       @               @              �?              �?              �?              @                                              @                                       @       @       @       @                              @              2@       @                      �?       @      @       @       @              @      �?      @       @                                              �?               @      @      @      @              �?      d@     �@@      ]@      $@      1@      @      <@     0x@     0r@      7@      5@     �K@     �r@     �e@      @      4@      "@      @@      &@     @T@      @     �J@      @      @              (@      n@      e@      &@       @      1@     �`@      V@              @      @      (@      @      "@              �?                                     �F@      *@                               @                                                                                                              (@      @                                                                                      "@              �?                                     �@@      @                               @                                                      �?              �?                                      1@      �?                              @                                                                                                              @                                      @                                                      �?              �?                                      $@      �?                                                                                       @                                                      0@      @                              @                                                      �?                                                      @      @                              �?                                                      @                                                      "@      @                              @                                                      R@      @      J@      @      @              (@     `h@     �c@      &@       @      1@     �_@      V@              @      @      (@      @      <@      @      @      �?       @              (@     �@@      B@      @              @      ;@      1@                       @      �?      @      6@      �?      �?      �?                      @      ;@      3@       @              @      2@      ,@                                      @       @                                                      ,@      �?                              @                                                      4@      �?      �?      �?                      @      *@      2@       @              @      .@      ,@                                      @      @      @      @               @               @      @      1@      @               @      "@      @                       @      �?               @                                              @              $@                       @      @       @                                              @      @      @               @              @      @      @      @                      @      �?                       @      �?              F@      @      G@       @       @                     @d@      ^@      @       @      &@      Y@     �Q@              @      �?      &@       @      4@              $@                                      <@     �E@      �?      �?      @      :@      4@              �?               @              @              @                                      9@      3@              �?      �?      "@      @                               @              .@              @                                      @      8@      �?              @      1@      *@              �?                              8@      @      B@       @       @                     �`@     @S@      @      @      @     �R@     �I@              @      �?      "@       @      @              9@              �?                     �W@     �F@      �?      @       @     �D@      9@              �?      �?      @      �?      1@      @      &@       @      �?                      D@      @@      @       @      @     �@@      :@              @              @      �?     �S@      :@     �O@      @      *@      @      0@     `b@     �^@      (@      *@      C@     @d@      U@      @      .@      @      4@      @      G@      0@      B@       @      "@      @      @      [@      U@      @      &@      4@     �]@      E@       @      @       @      "@       @      ?@      "@      0@      �?      @               @      C@      ,@      @      @      &@      K@      4@              �?              @       @      @      @      @              @               @       @      @      �?      @      �?      <@      @                                              @      @      @                                       @       @      �?      @      �?      :@      �?                                              �?                              @               @              �?                               @       @                                              9@      @      (@      �?      @                      >@      &@      @      @      $@      :@      1@              �?              @       @      $@       @       @               @                      "@       @      @      @      @      0@      @                              @      �?      .@      @      @      �?       @                      5@      @                      @      $@      $@              �?                      �?      .@      @      4@      �?       @      @      @     �Q@     �Q@      �?      @      "@      P@      6@       @       @       @      @              @      @      @      �?              @      �?      :@     �A@               @              (@      0@              �?      �?                      @      @      @      �?              @      �?      :@     �A@               @              "@      ,@              �?      �?                                      @                                                                              @       @                                              $@       @      *@               @              @      F@     �A@      �?       @      "@      J@      @       @      �?      �?      @               @       @      (@               @               @      A@      >@      �?       @      "@      I@      @       @      �?      �?      @               @              �?                               @      $@      @                               @                                                     �@@      $@      ;@      @      @      �?      "@     �C@      C@      @       @      2@      F@      E@       @      (@      @      &@      @      7@       @      @              �?              @      >@      A@               @      @      9@      ,@              $@      �?      @      �?      @       @      �?                              @       @       @                              &@      �?                                              @       @      �?                                      @       @                              $@                                                       @                                              @      �?                                      �?      �?                                              2@              @              �?              �?      6@      :@               @      @      ,@      *@              $@      �?      @      �?      (@              @                              �?      3@      $@                      �?      @      $@              @      �?              �?      @              �?              �?                      @      0@               @       @      @      @              @              @              $@       @      4@      @      @      �?      @      "@      @      @              .@      3@      <@       @       @      @      @       @                       @       @                      �?      @              �?              @      @      @                       @      @      �?                      �?      �?                               @              �?                       @      @                      �?      @                              �?      �?                      �?      @                              @      @      @                      �?              �?      $@       @      2@      @      @      �?      @      @      @      @               @      ,@      5@       @       @      �?      @      �?      @       @      @              @              @       @       @      @              @      �?      @               @      �?      �?      �?      @      @      .@      @              �?      �?      �?       @       @              @      *@      0@       @                       @        �t�bub��%     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ@��ThG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmK}hnh4h7K ��h9��R�(KK}��hu�BX         >                    �?�CD���?{	           ��@       !                    �?��R���?           �@                           �?�T�t<f�?-           @@                           �?������?�            �l@                            �?�m��1�?<             Z@                           3@      �?             D@������������������������       ��(ݾ�z�?             *@������������������������       �g�WH��?             ;@	       
                   �2@     ��?'             P@������������������������       �\���(\�?             4@������������������������       ���Z=;�?             F@                          �:@�W�\T�?M            @_@                            @P�_>L��?=            �X@������������������������       �=J�5��?$            �O@������������������������       ��q�q�?             B@                            @�Q�}e�?             :@������������������������       ���1G���?             *@������������������������       �*D>��?             *@                           �?Rk<��?�            �p@                          �9@c��@{��?8            @X@                            �?9��8���?,             R@������������������������       �<ݚ�?             2@������������������������       ��F&K:�?              K@                            �?a��+e�?             9@������������������������       �t�E]t�?             &@������������������������       ��Cc}�?             ,@                          �5@��F���?l            �e@                            �?�m%/[u�?<            �X@������������������������       �R���Q�?             4@������������������������       ��bs㷝�?/            �S@                           �7@h�ϱ���?0            �R@������������������������       ��h�*$��?             3@������������������������       �۶m۶m�?#             L@"       1                   �2@I�X�5�?�           @�@#       *                    �?Ev�Md�?�            �l@$       '                   �1@��	�g��?4            @V@%       &                     �?9��8���?             B@������������������������       �4%���?             1@������������������������       ��GcT!)�?
             3@(       )                     @�fXf��?            �J@������������������������       �zf<�n�?            �B@������������������������       �     ��?             0@+       .                    �?D��=�?T            `a@,       -                     �?*fW�Em�?"            �J@������������������������       ����Q��?             4@������������������������       ��(��r�?            �@@/       0                   �0@�撳g�?2            �U@������������������������       ��)x9/�?             ,@������������������������       ��������?+             R@2       9                   �=@;��P[�?R           `�@3       6                    �?�sx���?           Љ@4       5                   �5@dЅҶ9�?�             r@������������������������       ��!,*r�?A            @X@������������������������       ��??���?u             h@7       8                   �8@��QDBF�?V           ��@������������������������       �Z�ַ��?�            �v@������������������������       ���էR`�?q            �e@:       ;                    �?�H�K@��?F            �\@������������������������       �F]t�E�?             &@<       =                     �?~U98F��?@            �Y@������������������������       ���^B{	�?             B@������������������������       �bB�Fv6�?'            �P@?       ^                   �2@�����?t           ��@@       O                    �?�7^���?�           @�@A       H                   �1@ju�w�C�?�            pw@B       E                     �?�����W�?�             l@C       D                    @CbΊx�?"             M@������������������������       ����k���?             F@������������������������       �X�Cc�?	             ,@F       G                    @��dc� �?i            �d@������������������������       �P�|�@�?             A@������������������������       ��ͽ�n��?R            �`@I       L                     �?9EGr��?W            �b@J       K                    @���(\��?             D@������������������������       �K&:~��?             3@������������������������       ��3_<�?             5@M       N                    @�|@&|5�??            �[@������������������������       �[�&�p�?            �G@������������������������       �L���8�?"            �O@P       W                    @�ZƲ] �?�            s@Q       T                    @�(h�Ň�?J            @^@R       S                   �1@��}�f�?9            �V@������������������������       �v��n#�?$             O@������������������������       �~h����?             <@U       V                    @tF9i��?             ?@������������������������       �tk~X��?	             2@������������������������       �ݾ�z�<�?             *@X       [                    @���x�?{             g@Y       Z                   �1@�[��'��?V             `@������������������������       �t�c���?5            @S@������������������������       ��9J����?!             J@\       ]                     �?����?%            �K@������������������������       ����.�?             3@������������������������       ��Kh/��?             B@_       n                    @>�^:�y�?�           t�@`       g                   �9@���44�?�           ��@a       d                     �?��X����?.           ��@b       c                    �?8E�\@��?C           ��@������������������������       ��'�7O�?b             e@������������������������       �-<�Z�?�            �v@e       f                    �?��b�J��?�            �w@������������������������       ��N�u��?l            �e@������������������������       �Z�(�?            `j@h       k                   �:@FҊQ��?�             k@i       j                     �?&]^z���?#             M@������������������������       �      �?             @@������������������������       �;�;��?             :@l       m                    �?�)v+<J�?f            �c@������������������������       ��AE	��?(            @P@������������������������       ����{���?>            �W@o       v                     �? ��s'��?           @{@p       s                    �?��i���?�            �o@q       r                    @E��x���?F            �\@������������������������       �ôH�^�?>            �Y@������������������������       �Y�����?             &@t       u                    @�W����?Y            @a@������������������������       ��(AZs�?B            �Y@������������������������       �B{	�%��?             B@w       z                    �?��a���?w             g@x       y                   �8@��IU���?3            �R@������������������������       ������?&             K@������������������������       ��3_<�?             5@{       |                   �3@p��L��?D            @[@������������������������       ��q�q�?	             (@������������������������       ������?;            @X@�t�bh�h4h7K ��h9��R�(KK}KK��h��B8J       �~@     �R@     @v@      <@     @Q@      <@      T@     X�@     ��@     @U@     �R@     `b@     ��@     �x@      *@      N@      I@      a@      S@     �l@      ?@     �g@      (@     �E@      4@     �G@      ^@     �g@      C@     �G@      S@     �n@      g@      $@     �B@      @@      Q@     �J@      Y@      @     �H@      @      0@      "@      &@      C@     @Q@      @      @      *@      S@     �H@      �?      (@      &@      .@      &@      K@      @      3@      �?       @              @      6@      C@       @       @      @     �@@      2@      �?      @      @      @      @      2@      @      @                                      (@      =@       @      �?      @      *@      "@              @      @       @       @      "@              �?                                      @      *@                               @      �?                      @                      @              �?                                      @                                      @      �?                                              @                                                              *@                              @                              @                      "@      @      @                                      @      0@       @      �?      @      @       @              @               @       @      "@                                                      @      �?       @              @                                               @                      @      @                                      @      .@              �?              @       @              @                       @      B@      @      .@      �?       @              @      $@      "@              �?      @      4@      "@      �?       @              @      �?      6@      �?      .@      �?       @              @      $@      @                      @      1@      "@      �?      �?              @      �?      .@              *@      �?      �?              @      $@      �?                      @      &@      �?              �?              �?              @      �?       @              �?                              @                              @       @      �?                      @      �?      ,@       @                                       @              @              �?              @                      �?                              @       @                                       @              @                                                                                       @                                                                              �?              @                      �?                              G@      �?      >@       @      ,@      "@      @      0@      ?@      @      @      @     �E@      ?@              @       @       @       @      2@              @              @               @      @      (@              �?       @      5@      *@              @      @      �?       @      .@              @               @              �?      @      (@                       @      3@      @              @      �?      �?       @      @                                              �?      �?      @                      �?       @       @                              �?              (@              @               @                      @      @                      �?      1@       @              @      �?               @      @                              �?              �?                              �?               @      "@              @      @                                                      �?              �?                                               @      @                                              @                                                                              �?                       @              @      @                      <@      �?      ;@       @      &@      "@      @      "@      3@      @       @      @      6@      2@                      @      @      @      6@              ,@              @      @              "@      3@      �?       @      �?      *@       @                              �?       @      @               @                                              @                      �?      @                                      �?              2@              (@              @      @              "@      (@      �?       @               @       @                                       @      @      �?      *@       @      @      @      @                       @              @      "@      $@                      @      @      @      �?               @              @      @                                              �?      �?      @                      @                      @      �?      &@       @      @      �?      @                       @               @       @      @                              @      @      `@      8@     �a@      "@      ;@      &@      B@     �T@     �]@     �@@      E@     �O@      e@     �`@      "@      9@      5@     �J@      E@      A@       @      <@              �?              �?     �E@     �D@      @      �?      @     �D@      ,@               @      �?      "@      �?      1@      �?      @                                      (@      5@      @      �?      @      1@      @                              @      �?      *@                                                      @      @      @              �?      @                                      �?              @                                                      @      @      @              �?       @                                                      "@                                                      @       @                              @                                      �?              @      �?      @                                      @      .@              �?       @      &@      @                              @      �?       @              @                                      @      $@              �?       @      $@                                                       @      �?                                                      @                              �?      @                              @      �?      1@      �?      6@              �?              �?      ?@      4@                      @      8@      &@               @      �?      @              $@      �?      @                                      0@      @                              *@       @              �?              �?              @      �?                                              �?      @                               @                                                      @              @                                      .@      �?                              @       @              �?              �?              @              3@              �?              �?      .@      ,@                      @      &@      "@              �?      �?      @               @              @                                      @      @                                                                                      @              .@              �?              �?      $@      &@                      @      &@      "@              �?      �?      @             �W@      6@      \@      "@      :@      &@     �A@     �C@     �S@      >@     �D@     �L@     �_@     @^@      "@      7@      4@      F@     �D@     @V@      5@     �Y@      @      0@      @      ?@     �C@     �P@      6@     �A@     �H@     @_@     @]@      @      .@      0@     �A@      ?@     �E@      @      @@              "@              "@      3@      0@      @       @      (@     �P@     �B@              �?      @      $@      (@      1@      @      $@              �?              @      $@      @      @      �?      &@      .@      &@                       @       @              :@       @      6@               @              @      "@      $@      @      @      �?     �I@      :@              �?       @       @      (@      G@      0@     �Q@      @      @      @      6@      4@      I@      .@      ;@     �B@     �M@      T@      @      ,@      (@      9@      3@     �A@      $@      G@      @      @      @      &@      3@      C@      @      6@      6@     �C@      N@              @       @      6@       @      &@      @      9@      �?      @              &@      �?      (@       @      @      .@      4@      4@      @      $@      $@      @      &@      @      �?      "@       @      $@      @      @              (@       @      @       @       @      @      @       @      @      "@      $@                                                                              �?                              �?      �?       @              @      �?      @      �?      "@       @      $@      @      @              (@      @      @       @       @      @      @      @      @      @      "@              �?       @      �?              @      @              @      �?      @      @               @               @       @      �?      @      @              @      �?      $@       @                       @      @      �?      @       @      �?      @      @       @      @      @     0p@     �E@     �d@      0@      :@       @     �@@     0{@     �y@     �G@      <@     �Q@      v@     �j@      @      7@      2@      Q@      7@     @S@      @     �@@                              @     @k@      d@      @      @      .@      W@     �F@              @      @      $@       @      D@      @      "@                               @      a@     �Y@      �?      �?      @     �G@      :@                                              :@       @      @                               @     �V@      N@              �?      �?     �@@      @                                               @                                              �?      ;@      5@              �?              @                                                       @                                              �?      6@      (@              �?              @                                                                                                              @      "@                                                                                      8@       @      @                              �?      P@     �C@                      �?      ;@      @                                              @                                                      @      *@                              @                                                      1@       @      @                              �?     �L@      :@                      �?      4@      @                                              ,@       @      @                                      G@     �E@      �?              @      ,@      6@                                              �?       @      �?                                      @      4@                      @      @      @                                                              �?                                      �?      (@                      @      �?                                                      �?       @                                               @       @                              @      @                                              *@              @                                     �E@      7@      �?                      $@      1@                                              &@              @                                      *@      "@                              @       @                                               @                                                      >@      ,@      �?                      @      "@                                             �B@       @      8@                              @     @T@      M@      @       @      $@     �F@      3@              @      @      $@       @      4@       @      1@                              �?      *@      7@      @       @      @      7@      "@                      �?       @              2@       @      ,@                                      *@      "@      @       @      @      2@      @                      �?                      $@      �?      ,@                                      "@      @               @      @      &@      @                                               @      �?                                              @       @      @                      @       @                      �?                       @              @                              �?              ,@                      �?      @      @                               @                              @                                              *@                                                                       @               @                                              �?              �?                      �?      @      @                                              1@              @                               @      Q@     �A@                      @      6@      $@              @       @       @       @      &@              @                              �?     �L@      7@                      @      *@      "@                              �?       @      @              �?                                      ?@      2@                      @       @      @                              �?              @              @                              �?      :@      @                      �?      @       @                                       @      @                                              �?      &@      (@                              "@      �?              @       @      @               @                                              �?      "@      �?                              �?                               @      @              @                                                       @      &@                               @      �?              @              @             �f@     �B@     �`@      0@      :@       @      <@      k@      o@     �E@      9@      L@     @p@     @e@      @      1@      .@      M@      5@     �^@      ;@     @U@      $@      0@       @      2@     �d@     �h@      =@      0@     �C@      i@     �`@       @      $@      @      @@      *@     �Z@      4@      O@      $@      @      @      .@      b@      g@      (@      *@      >@     `d@     @Y@      �?      @      @      6@       @      O@       @     �C@      @      �?      �?      $@     �Q@     �\@      $@      @      ,@      W@     �Q@              @      @      &@      @      1@      @      @                      �?       @      4@      K@       @      @      @      <@      8@              �?                      �?     �F@      @      @@      @      �?               @     �I@     �N@       @      @       @      P@     �G@              @      @      &@      @      F@      (@      7@      @      @      @      @     �R@     �Q@       @      @      0@     �Q@      >@      �?                      &@      @      1@      @      @      �?      �?                      H@      <@       @      @      "@      @@      *@                              @              ;@      @      0@      @      @      @      @      :@      E@               @      @     �C@      1@      �?                      @      @      0@      @      7@              "@      @      @      3@      (@      1@      @      "@     �B@     �@@      �?      @      @      $@      @      @              @                                      @      �?                       @      .@      *@              @              @      @      @              @                                              �?                              *@      @                              @               @              @                                      @                               @       @      @              @                      @      "@      @      0@              "@      @      @      .@      &@      1@      @      @      6@      4@      �?      @      @      @       @      @       @      @              @                      *@      @      �?      @      @      .@      @               @              @              @      @      $@              @      @      @       @      @      0@              @      @      0@      �?      �?      @      @       @      N@      $@     �H@      @      $@              $@     �J@      J@      ,@      "@      1@      N@      B@      �?      @       @      :@       @      @@       @      <@      @      @              �?     �F@     �@@      @      @      ,@      >@      5@              @      @      0@       @      2@               @      �?                              9@      5@       @      @      @      (@      &@               @              @              (@               @      �?                              9@      5@       @      @      @       @      &@              �?              @              @                                                                                              @                      �?                              ,@       @      4@       @      @              �?      4@      (@      @      �?      "@      2@      $@              �?      @      *@       @      @       @      1@       @       @              �?      ,@       @      @              @      1@      @                      @      *@      �?       @              @               @                      @      @              �?      @      �?      @              �?                      �?      <@       @      5@      @      @              "@       @      3@      "@       @      @      >@      .@      �?      @       @      $@      @      $@      @      @              �?               @      @      "@      @       @      �?      3@      @              �?              @              @              @              �?               @      @      "@      @       @      �?      &@      @                              @              @      @       @                                       @                                       @                      �?                              2@      @      ,@      @      @              @      @      $@      @               @      &@      (@      �?      @       @      @      @                                                      �?              @                                      @              �?                              2@      @      ,@      @      @              @      @      @      @               @      &@      @      �?       @       @      @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ(�ihG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKuhnh4h7K ��h9��R�(KKu��hu�B�         >                     @�^�6��?�	           ��@                          �2@�;��Z�?�           X�@                           �?%a����?�           @�@                           �?�����?�            Px@                           �?W�7�L\�?0             U@                            �?�8��8��?             8@������������������������       ���8��8�?             (@������������������������       ��8��8��?             (@	       
                    �?�i�6��?!             N@������������������������       ��>�>�?             >@������������������������       ��`�`�?             >@                          �1@9�����?�            s@                           @j|�����?~             h@������������������������       �����_�?+            �S@������������������������       �3�<�K��?S            �\@                           @��>4��?I             \@������������������������       �h�!Ԣ�?<            �V@������������������������       ���ճC��?             6@                          �0@���_N��?�            0v@                            �?"��K�[�?'             O@                           �?VUUUU��?             H@������������������������       �     ��?	             0@������������������������       �      �?             @@������������������������       ���X��?	             ,@                           @r���lL�?�            Pr@                            �?�W�3�?�            �j@������������������������       �E�ϣ1��?e             c@������������������������       �쌯�t��?'             O@                           �?\��nS��?0            �S@������������������������       ��]�`��?             *@������������������������       �Oq����?(            �P@        /                   �8@xZc�2��?�           �@!       (                    �?��O�B8�?Q           ��@"       %                   �5@��~�݇�?            |@#       $                    �?9\*�U�?�            �m@������������������������       ����2p �?H            @Z@������������������������       ���WƐ�?N            ``@&       '                   �7@Ƿ�.�S�?�            �j@������������������������       �Ľͫm��?]            @c@������������������������       �t�@��?&             N@)       ,                    �?���&��?8           �@*       +                    @'�qG���?�            0u@������������������������       ��@?�1��?�            �g@������������������������       �)[�0��?_            �b@-       .                    �?Ku�$��?V           P�@������������������������       ��M�j��?�             o@������������������������       �C���l�?�             s@0       7                   �=@-�1�?�           (�@1       4                    @�WϊF�?7            ~@2       3                    �?�=vQ�?�            �u@������������������������       �b���j��?k             e@������������������������       �H�5U��?v             f@5       6                    @���x�?V            �`@������������������������       ��Y]�S�?1            @S@������������������������       ��Rpo�?%             M@8       ;                     �?��j[v�?h            �d@9       :                    �?��hZ�?H             ]@������������������������       ���7���?            �G@������������������������       ���ؗ���?,            @Q@<       =                    @�3���?             �H@������������������������       �j�V���?            �@@������������������������       �     @�?             0@?       \                   �4@b��o���?�           t�@@       O                   �1@�\�PZ��?[           ��@A       H                    �?��+�M�?h            �c@B       E                    �?��3Q�?1            �Q@C       D                    �?c>���?             5@������������������������       ��q�q�?             (@������������������������       ������H�?             "@F       G                   �0@гY����?"             I@������������������������       �      �?             (@������������������������       �]��N��?             C@I       L                    �?h�b�{8�?7            �U@J       K                    �?�̿0�=�?             ?@������������������������       �r�q��?	             (@������������������������       �"P7��?             3@M       N                    @���>4��?#             L@������������������������       ��9����?             6@������������������������       ���'s�	�?             A@P       W                    �?]�R����?�            pw@Q       T                    @�L�_�?l            �c@R       S                   �3@�.k���?Z             a@������������������������       �K�'��n�?>            @X@������������������������       ��B�����?            �C@U       V                    �?'�%����?             7@������������������������       �z�G�z�?             $@������������������������       ��K8��?             *@X       [                    @zۧ���?�             k@Y       Z                    @�EG����?x            �g@������������������������       � jA��?a            @c@������������������������       ���¤�h�?             A@������������������������       �������?             <@]       j                    @�����W�?�           @�@^       e                    �?�ʆ'*��?C           �@_       b                    �?�ued��?           p{@`       a                    @�?��V��?h             e@������������������������       �ԥxP��?O            �^@������������������������       �Ĭ뉳��?             G@c       d                   �@@�"�n���?�            �p@������������������������       �    ���?�             p@������������������������       �d}h���?	             ,@f       i                    @���yZ�?+            �R@g       h                   �<@�I��i�?%            �O@������������������������       ����B���?            �G@������������������������       �     @�?             0@������������������������       �r�q��?             (@k       r                   �;@@��TM�?S            �`@l       o                   �5@��cԧ�?E            @[@m       n                    �?������?             ?@������������������������       �c>���?             5@������������������������       ��G�z��?             $@p       q                   �6@e(��#�?3            �S@������������������������       �ŕ�(�?             5@������������������������       �n�Y���?%            �L@s       t                   �=@p_�Q�?             9@������������������������       �I�$I�$�?             ,@������������������������       ��ˠT�?             &@�t�bh�h4h7K ��h9��R�(KKuKK��h��BxE       �z@     @U@     pu@      @@     �P@      9@     @S@     ��@     ��@     �Q@      S@      g@     ȃ@     0z@      2@     @R@     �J@     �^@     �M@      s@      J@     `n@      1@     �A@      "@      J@     �{@     p|@     �K@     �J@     �\@     �z@     �p@       @     �G@     �A@      T@      B@      W@      (@      :@              �?              (@     �k@     `d@      @      @      6@     �`@     �A@               @      �?      "@      @     �J@      @      "@                              @     �a@     �W@                      @     �L@      4@                              �?              6@       @      @                                      :@      (@                      @      "@      �?                                              @              @                                      *@      �?                      �?              �?                                              @              �?                                      @                                                                                                               @                                      @      �?                      �?              �?                                              1@       @      @                                      *@      &@                      @      "@                                                       @              @                                      $@      @                      @      @                                                      .@       @      �?                                      @      @                              @                                                      ?@      @       @                              @     �\@     �T@                       @      H@      3@                              �?              5@       @                                      @     �T@      I@                      �?      ?@       @                              �?              @       @                                       @      A@      8@                              @       @                              �?              ,@                                              �?      H@      :@                      �?      9@                                                      $@      �?       @                                      @@      @@                      �?      1@      1@                                              @               @                                      >@      6@                      �?      .@      .@                                              @      �?                                               @      $@                               @       @                                             �C@      @      1@              �?              "@     @T@     @Q@      @      @      .@     @S@      .@               @      �?       @      @      (@              �?                                      &@      1@                      �?      3@      �?                                              @              �?                                       @      1@                      �?      .@      �?                                              �?                                                      @      "@                              @                                                      @              �?                                      @       @                      �?      (@      �?                                              @                                                      @                                      @                                                      ;@      @      0@              �?              "@     �Q@      J@      @      @      ,@      M@      ,@               @      �?       @      @      6@      @      *@              �?              @      I@      @@      @      @      "@     �H@      @                      �?      @      @      5@      @      @              �?              @      =@      3@      @      @       @     �A@      @                      �?      @      @      �?              @                               @      5@      *@       @              �?      ,@      �?                                              @              @                              @      4@      4@      �?              @      "@      @               @              @      �?      �?              �?                                              @      �?               @       @                                                      @               @                              @      4@      ,@                      @      @      @               @              @      �?     �j@      D@      k@      1@      A@      "@      D@      l@     @r@     �H@     �H@     @W@     �r@     �l@       @     �F@      A@     �Q@      @@      e@      0@     @c@      $@      *@      �?      4@     @g@     �l@      7@      7@      H@     @j@     �b@      �?      8@      &@     �A@      3@      R@      @     @P@       @       @              &@     �@@      D@      $@      .@      1@     �M@     �Q@              &@      @      .@      (@      G@      �?      8@       @      �?              @      1@      <@      �?       @      &@      :@      C@              @              *@       @      =@              @              �?               @      @      ,@      �?      @      @      4@       @               @              �?       @      1@      �?      1@       @                      @      $@      ,@              �?      @      @      >@              @              (@      @      :@      @     �D@              @              @      0@      (@      "@      @      @     �@@     �@@              @      @       @      @      5@       @     �@@              @              �?      @      &@      @      @      @      <@      3@              @      @      �?       @      @      �?       @               @              @      "@      �?      @       @       @      @      ,@                              �?       @      X@      (@     @V@       @      @      �?      "@      c@     �g@      *@       @      ?@     �b@     �S@      �?      *@      @      4@      @     �@@      @      3@      @              �?      @      K@     �U@       @              $@      P@      E@               @              @      @      (@      @      &@      @              �?      �?      7@     �I@       @               @     �E@      9@               @              �?       @      5@      �?       @                               @      ?@      B@                       @      5@      1@              @              @      �?     �O@      @     �Q@      @      @              @     �X@      Z@      &@       @      5@     �U@     �B@      �?      @      @      .@      @      9@      �?      B@      �?                      �?     �K@     �K@      @       @      @     �B@      1@              �?      �?      @       @      C@      @      A@      @      @              @      F@     �H@      @      @      2@      I@      4@      �?      @      @      "@       @      F@      8@     �O@      @      5@       @      4@      C@     �N@      :@      :@     �F@     �U@     @T@      �?      5@      7@      B@      *@     �A@      3@      M@      @      *@       @      .@     �A@     �G@      1@      2@      7@      R@     �M@      �?      0@      *@      5@      (@      5@      0@     �G@      @      &@       @      "@      =@      D@      ,@      0@      (@      E@     �C@      �?      &@      *@      .@      @      (@      $@      2@       @      @      �?      @      @      .@      @      $@      "@      3@      6@      �?      @      &@       @      @      "@      @      =@      �?      @      �?      @      8@      9@      @      @      @      7@      1@              @       @      @      �?      ,@      @      &@      �?       @              @      @      @      @       @      &@      >@      4@              @              @       @      @       @      "@      �?      �?              @              @      �?      �?      @      1@      &@              @              @       @      &@      �?       @              �?               @      @      @       @      �?      @      *@      "@                                              "@      @      @      @       @      @      @      @      ,@      "@       @      6@      .@      6@              @      $@      .@      �?       @      @      @       @       @      @      @       @      (@      @      @      5@      @      0@              @      @       @      �?      @              �?               @              @       @      @      �?       @      @      @      "@              �?      �?       @      �?       @      @       @       @              @       @              @      @      @      0@       @      @              @      @      @              �?       @       @      �?      @       @              �?       @      @       @      �?      "@      @                      @      @              �?       @              �?      �?       @              �?              �?       @      �?      "@      @                      @      @                               @              @                               @       @                                                      �?      @             �^@     �@@      Y@      .@      ?@      0@      9@     �X@     �b@      .@      7@     �Q@     @i@      c@      0@      :@      2@     �E@      7@     @R@      @      G@       @      "@      �?      @     @Q@     �T@      @      *@      6@     �[@      L@              @       @      3@      @      <@              .@               @                     �A@      8@      @              @      7@      0@              @               @              2@              @               @                      (@      @      �?              @      @      *@              @              �?              @               @                                      @       @      �?              �?               @                              �?              @                                                      @       @      �?              �?                                                               @               @                                       @                                               @                              �?              *@              @               @                      @      @                       @      @      &@              @                              @              �?                                      �?       @                              �?       @                                               @              @               @                      @      �?                       @      @      "@              @                              $@               @                                      7@      3@       @              @      1@      @              �?              �?              @              @                                       @      @                      �?      $@      �?                                              �?               @                                      �?       @                              @                                                      @              @                                      �?      @                      �?      @      �?                                              @               @                                      5@      *@       @               @      @       @              �?              �?              �?               @                                      @      @       @                      @      �?                              �?              @                                                      2@      @                       @      �?      �?              �?                             �F@      @      ?@       @      @      �?      @      A@     �M@              *@      0@      V@      D@               @       @      1@      @      @              *@              @      �?      @      8@      <@              @      @      C@      6@                               @      �?      @              *@              @      �?      @      8@      ;@              @       @     �@@      &@                              @      �?      @              @                              @      4@      6@              �?       @      8@      "@                              @      �?      @              @              @      �?              @      @              @              "@       @                              �?              �?                                              �?              �?               @      �?      @      &@                              �?                                                                                                               @       @                                              �?                                              �?              �?               @      �?      @      @                              �?              C@      @      2@       @      @              @      $@      ?@              @      *@      I@      2@               @       @      "@      @      @@      @      2@       @      @              �?      @      8@              @      *@     �G@      0@              �?       @      @      @      ;@      @      .@       @      @              �?      @      5@              @      @     �C@      ,@              �?      �?      @      @      @              @                                              @                      "@       @       @                      �?      @              @                                               @      @      @                              @       @              �?               @              I@      ;@      K@      *@      6@      .@      2@      =@      Q@      (@      $@      H@     �V@     @X@      0@      4@      0@      8@      2@     �A@      3@      E@      *@      5@      .@      ,@      1@     �K@      (@      $@      F@      P@      R@      *@      4@      *@      1@      2@      >@      1@     �D@      &@      4@      .@      $@      (@      C@      $@      $@     �@@     �M@      O@      &@      2@      *@      ,@      .@      .@       @      1@      @      @      �?      @      @      1@      �?       @      (@      B@      8@       @      @      @      @      @      *@      �?      .@      @       @      �?      @      @      1@      �?      �?      "@      1@      .@      �?      @      @      @      @       @      �?       @       @       @                      @                      �?      @      3@      "@      �?              �?                      .@      .@      8@      @      0@      ,@      @      @      5@      "@       @      5@      7@      C@      "@      (@      "@       @      $@      .@      .@      8@      @      0@      ,@      @      @      5@      "@      @      4@      7@      C@       @      (@       @       @      @                                                                                       @      �?                      @              �?              @      @       @      �?       @      �?              @      @      1@       @              &@      @      $@       @       @              @      @      @       @      �?       @                      @      @      .@       @              @      @      "@       @       @              @      @      @       @      �?       @                      @      @      .@                              @       @                              �?      @                                                               @               @              @              �?       @       @               @               @                              �?                               @                      @              �?                                              .@       @      (@              �?              @      (@      *@                      @      ;@      9@      @              @      @              .@      @      @              �?              �?      (@      $@                      @      4@      9@      @              @      @              @               @                                       @                              @      @      @                       @      �?               @               @                                      @                                      @       @                       @      �?              @                                                       @                              @               @                                              $@      @      @              �?              �?      @      $@                              ,@      5@      @              �?      @               @                                                       @      @                              @      "@                                               @      @      @              �?              �?       @      @                              "@      (@      @              �?      @                      @      @                              @              @                      �?      @                                      @                       @       @                              @                                              @                                      @                      �?      @                                              @                      �?      @                                                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJS��DhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKqhnh4h7K ��h9��R�(KKq��hu�B�         4                    �?�h��?�	           ��@                          �2@��>"!�?           ��@       
                    �?-�xؙ��?�             u@       	                    @����X�?\             b@                           @��?"md�?R            �_@                          �0@|���g�?D            �Y@������������������������       �      �?             0@������������������������       ���Aw��?8            �U@������������������������       �36�v[�?             7@������������������������       �3�R�f�?
             3@                           �?� ���?�             h@                           �?bX�h��?#            �K@                             @���Mb�?             9@������������������������       ��g���e�?             &@������������������������       �h�����?             ,@                          �1@��.�?�?             >@������������������������       �F]t�E�?             6@������������������������       �      �?              @                            �?oZ���?]            @a@                           @p_�Q�?             I@������������������������       ��}�!��?            �C@������������������������       ����k���?             &@                           @����|��?B             V@������������������������       �333333�?             4@������������������������       �� =[y�?2             Q@       '                    �?���Z\=�?:           l�@                            �?�1'��?�             w@                          �=@��;�?P             ]@                           �?�#*�6�?J             [@������������������������       �����S��?%             L@������������������������       ���ջ���?%             J@������������������������       �      �?              @!       $                    �?���R�?�            �o@"       #                     @��۾%d�?D             ]@������������������������       �#>�֕�?(            �Q@������������������������       �"*w�?             G@%       &                   �5@d�&���?Y            @a@������������������������       ���&�'�?'             O@������������������������       �d{�ԍ�?2             S@(       -                    �?���/�O�?M           H�@)       ,                   @@@�C��2��?�             v@*       +                   �6@�}D��?�            @u@������������������������       �,^��K��?[             c@������������������������       �Qf]�?x            `g@������������������������       �      �?             (@.       1                    @�$K�DJ�?s           H�@/       0                     �?�����?\             b@������������������������       ����&��?            �A@������������������������       ������?B            �[@2       3                   �?@En���-�?           �{@������������������������       �D��R��?           �y@������������������������       �     ��?             @@5       T                    �?���fx��?�           ��@6       E                    @�ƓXA��?�           ��@7       >                   �2@ۙ>�m��?           @�@8       ;                    @�&���?�            �s@9       :                    @,VN�@�?{            �h@������������������������       �U���f��?Q            ``@������������������������       �&5DSb�?*             Q@<       =                   �0@{��r���?P            �\@������������������������       ��Q����?            �A@������������������������       ���Q���?9             T@?       B                   �9@,�ρ^�?M           p�@@       A                    �?��G*M�?           �y@������������������������       �����X��?�             l@������������������������       ��J/1i�?|            �g@C       D                   �=@�O�
��?@            @\@������������������������       ����,��?1            @W@������������������������       ��Q����?             4@F       M                     �?_LMEj�?�            �q@G       J                   �5@>�� =��?*             O@H       I                    @���?            �C@������������������������       �Z�K8�?             :@������������������������       �����W�?             *@K       L                    @\")�i��?             7@������������������������       �9��8���?	             (@������������������������       �b���i��?             &@N       Q                   �2@(w�r(�?�            �k@O       P                    @s
^N���?%             L@������������������������       ��:��aZ�?            �C@������������������������       ��P�n#�?             1@R       S                    @�8=���?h            �d@������������������������       �P1��w�?            �C@������������������������       ���h���?P            @_@U       d                     @�b}�?�           �@V       ]                   �5@HP��$S�?J           x�@W       Z                    @QM�����?X           `�@X       Y                   �0@ͿN,���?�            `o@������������������������       ��q�q�?             8@������������������������       �B��"�C�?�            `l@[       \                     �?.��� |�?�            q@������������������������       �?4ևƺ�?E             \@������������������������       ���=�1��?o             d@^       a                   �:@ށ?n���?�            0x@_       `                    @���d���?�            �p@������������������������       ��y/���?y            @g@������������������������       �w�_���?/            �S@b       c                     �?����6��?J            �^@������������������������       �z�:���?/            @U@������������������������       ���4mx�?            �B@e       j                   �3@��ZNA��?�            `m@f       i                    @�s��?@            �Y@g       h                    �?��+���?*            @Q@������������������������       ��>d?�?�?            �G@������������������������       �ֳC��2�?             6@������������������������       ��1�^��?             A@k       n                    �?�zv��?V            �`@l       m                   �6@�n(T��?            �@@������������������������       �UUUUUU�?             (@������������������������       ��3_<�?             5@o       p                   �7@�7�j���?A            �X@������������������������       �ڃ����?            �K@������������������������       �$��Z=;�?"             F@�t�bh�h4h7K ��h9��R�(KKqKK��h��BC       �|@     �V@     `w@      >@     @R@      8@     @T@     ��@     H�@      N@     �U@     �a@     ؂@     �y@      (@      Q@     �H@     �b@     �B@     �g@     �E@     �f@      *@      I@      5@      I@     @\@     �g@      ?@     �J@     @T@     �m@      i@      @      F@      @@     �U@      7@      I@      @      7@              �?              @      K@     �L@               @       @     �P@      6@              @      �?      ?@       @      9@      @       @                              �?      1@      9@              @      @      A@      @              @              .@       @      5@      @      @                              �?      1@      9@               @      @      :@      @              @              *@       @      5@      @      @                              �?      0@      0@               @      @      8@       @              @              @              @              �?                                      @      @                              �?                                                      0@      @       @                              �?      *@      $@               @      @      7@       @              @              @                               @                                      �?      "@                               @      �?                              @       @      @              @                                                               @               @                                       @              9@       @      .@              �?               @     �B@      @@              @      @     �@@      3@              @      �?      0@              @      �?                      �?                       @      $@              �?      �?      ,@      @                              $@               @      �?                                              @                                      @       @                              "@                                                                      @                                      @      �?                                               @      �?                                                                                      �?      �?                              "@              @                              �?                      �?      $@              �?      �?      $@       @                              �?              @                              �?                      �?      @                              "@       @                                                                                                              @              �?      �?      �?                                      �?              4@      �?      .@                               @      =@      6@              @       @      3@      .@              @      �?      @              $@      �?       @                              �?      *@      @               @              $@      @                                               @      �?       @                              �?      @      @               @              $@      @                                               @                                                      @                                               @                                              $@              *@                              �?      0@      2@              �?       @      "@       @              @      �?      @               @              @                              �?      @      @              �?                       @                              @               @              "@                                      (@      .@                       @      "@      @              @      �?      @             `a@      C@     �c@      *@     �H@      5@     �G@     �M@     �`@      ?@     �F@     @R@     @e@     @f@      @      C@      ?@      L@      5@     @Q@      $@     �B@       @      $@      �?      (@      0@     �J@       @      &@      ,@      G@     �F@              $@      @      *@      @      *@      @      @               @              @       @      <@      @      "@      �?      *@      *@              @      @      �?      �?      (@      @      @              �?              @       @      <@      @      @      �?      *@      &@              @      @      �?      �?      @      @      @                                      @      4@              �?      �?      "@      @               @              �?              @              �?              �?              @      @       @      @      @              @       @              @      @              �?      �?                              �?                                              @                       @                                              L@      @      >@       @       @      �?       @       @      9@      @       @      *@     �@@      @@              @      @      (@      @      >@       @      *@      �?      @              @              1@               @      @      .@      0@               @              @              2@               @      �?      @              @              $@               @      @      "@      @                              @              (@       @      @                                              @                              @      $@               @               @              :@      @      1@      �?      @      �?      @       @       @      @              "@      2@      0@              �?      @      @      @      3@       @      @                              @      @      @       @               @      @      @                              @              @      @      *@      �?      @      �?              �?      �?      @              @      (@      &@              �?      @      �?      @     �Q@      <@     �^@      &@     �C@      4@     �A@     �E@      T@      7@      A@     �M@      _@     �`@      @      <@      8@     �E@      .@      B@      @     �C@       @      (@      @      .@      :@     �F@      @      (@      1@      M@      D@      �?      ,@      &@      @      @      B@      @     �C@       @      @      @      *@      :@     �F@      @      &@      1@      M@      D@              (@      $@      @      @      3@              .@      �?      @      @      @      2@      2@      �?      @      @     �A@      4@              @              �?      �?      1@      @      8@      �?      @              "@       @      ;@       @      @      ,@      7@      4@               @      $@      @      @                                      @               @                              �?                              �?       @      �?                      A@      6@     �T@      "@      ;@      1@      4@      1@     �A@      4@      6@      E@     �P@     @W@      @      ,@      *@      B@      $@      @      @      $@      @       @       @      @      @      3@      @      @      @      8@      7@       @      @      �?      (@              �?      @      @              �?              �?      @      @              �?      �?      "@      @              @      �?                      @              @      @      @       @       @       @      0@      @      @      @      .@      2@       @      @              (@              ;@      3@     @R@      @      3@      .@      1@      (@      0@      0@      .@      B@      E@     �Q@      @       @      (@      8@      $@      ;@      3@      Q@       @      3@      (@      1@      (@      0@      .@      ,@      <@      E@     �Q@               @      $@      5@       @                      @      @              @                              �?      �?       @                      @               @      @       @      q@     �G@      h@      1@      7@      @      ?@     �|@     �x@      =@     �@@      N@     �v@     �j@      @      8@      1@      O@      ,@     �a@      2@     �T@      �?      @              &@      q@     �n@      &@      .@      6@     �f@     @U@              @      �?      5@      @      [@      $@     �L@              @              @     �i@     �i@      @      "@      1@     �_@     @P@              @      �?      $@      @      B@              5@                               @      `@     �P@      �?      �?      @      F@      &@                                              :@              4@                               @     �P@      E@              �?      @      ?@      @                                              4@              @                              �?     �G@      =@              �?      �?      4@      @                                              @              .@                              �?      4@      *@                       @      &@                                                      $@              �?                                     �N@      8@      �?              �?      *@      @                                              @              �?                                      6@      @                               @                                                      @                                                     �C@      3@      �?              �?      &@      @                                              R@      $@      B@              @              @     �S@     �a@      @       @      *@     �T@      K@              @      �?      $@      @     �H@      @      7@                              @     @P@     ``@      @      @      "@     �N@      G@              �?      �?       @      @      ?@      @      $@                              �?      :@     @R@               @      @     �B@      @@                      �?       @              2@              *@                              @     �C@      M@      @      @      @      8@      ,@              �?              @      @      7@      @      *@              @                      ,@      "@       @      @      @      6@       @               @               @              7@      @      "@              @                      *@      @       @       @      @      (@      @               @               @                              @                                      �?       @              �?              $@       @                                             �@@       @      :@      �?      �?              @     @P@     �D@      @      @      @     �K@      4@                              &@              0@              @                              �?      @      1@              �?              "@      @                                              @              @                                      @      .@                              "@      �?                                               @                                                       @      .@                              @      �?                                              @              @                                      �?                                      @                                                      $@               @                              �?      @       @              �?                      @                                              @               @                                      @      �?                                                                                      @                                              �?              �?              �?                      @                                              1@       @      3@      �?      �?              @     �M@      8@      @      @      @      G@      .@                              &@              @              @                                      7@      (@      �?              �?      $@       @                                              @              @                                      1@       @                              @       @                                              �?                                                      @      @      �?              �?      @                                                      *@       @      0@      �?      �?              @      B@      (@      @      @      @      B@      *@                              &@              �?       @       @                                      @      @                       @      &@      @                              �?              (@      @       @      �?      �?              @      >@       @      @      @       @      9@      "@                              $@             �`@      =@     @[@      0@      1@      @      4@     �g@     �b@      2@      2@      C@      g@      `@      @      5@      0@     �D@      &@     @Z@      7@     �R@      &@      ,@       @      &@     �d@     �]@      1@      ,@      =@      c@      Y@       @      4@      0@      ;@       @     �R@      @      7@              @      �?      @     �a@     �T@      �?       @      .@      T@      M@              @      @      *@      @      B@       @      @               @      �?      �?     �V@     �@@      �?      @      @      :@     �@@              �?      @      �?      @       @                                                      2@      @                              �?                                                      A@       @      @               @      �?      �?     @R@      >@      �?      @      @      9@     �@@              �?      @      �?      @      C@      @      0@               @              @     �I@     �H@              @       @      K@      9@              @      @      (@      �?      (@      �?      @                                      9@      ;@              �?      @      4@      $@               @      �?      @              :@       @      (@               @              @      :@      6@              @      @      A@      .@              �?       @      @      �?      ?@      2@      J@      &@      $@      �?      @      9@      B@      0@      @      ,@      R@      E@       @      0@      $@      ,@      @      6@      (@      :@      "@      @      �?      @      8@      >@      @      @      "@     �M@      <@      �?      (@      @       @              ,@       @      ,@      @      @      �?      @      3@      <@       @      @      @     �H@      .@      �?      @              @               @      @      (@      @       @                      @       @       @              @      $@      *@              @      @      @              "@      @      :@       @      @              �?      �?      @      (@      �?      @      *@      ,@      �?      @      @      @      @      @      @      3@               @                      �?              (@              @      (@      &@              @      @      @      �?      @      @      @       @       @              �?              @              �?      �?      �?      @      �?                      �?      @      <@      @      A@      @      @      �?      "@      6@      >@      �?      @      "@      @@      =@      @      �?              ,@      @      &@              8@      @      �?              �?      $@      .@              @      @      (@      (@                              @              $@              5@       @      �?              �?      "@      "@              �?      �?      @       @                                               @              .@       @      �?              �?       @      @              �?      �?      @       @                                               @              @                                      @      @                               @                                                      �?              @       @                              �?      @              @      @      @      @                              @              1@      @      $@      �?       @      �?       @      (@      .@      �?              @      4@      1@      @      �?              &@      @      @      @              �?      �?                      @      "@                      �?       @      @                              @       @       @                      �?                              @                                               @                              �?       @      �?      @                      �?                              "@                      �?       @      �?                              @              ,@      @      $@              �?      �?       @       @      @      �?               @      2@      ,@      @      �?              @      �?      "@              @              �?               @      @      @                      �?      0@      @       @                      @      �?      @      @      @                      �?      @      @       @      �?              �?       @      $@       @      �?              �?        �t�bub��     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJc��hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKihnh4h7K ��h9��R�(KKi��hu�B�         6                    �?�����?�	           ��@       !                     @����?z           ��@                            �?�W��}�??           ��@                           �?�@:��?6           |@                          �1@Ug-��?n            `e@                          �0@9��8�#�?             H@������������������������       ��5;j��?             5@������������������������       �0���?             ;@	       
                   �7@d�y2A��?R            �^@������������������������       �X�EQ]N�?:            �U@������������������������       ������?            �B@                           �?��G�?�            `q@                          �4@�O�f��?             �G@������������������������       ���ӭ�a�?             2@������������������������       �v��`��?             =@                           �?����!�?�            �l@������������������������       ��G�z��?             $@������������������������       ��pA��?�            �k@                           @0���:*�?	           ��@                           @̦��4�?�            @s@                          �4@��J�e-�?�            �q@������������������������       ��GXwk�?J            �^@������������������������       �W%c3���?m            @d@                           6@@��Z��?             7@������������������������       ��9����?             &@������������������������       ��q�q�?             (@                          �4@�	�'/�?E           �@                           �?ro->Ԓ�?�            Pq@������������������������       �Y��L/1�?Q            @_@������������������������       �UH�� �?c             c@                            @���ə5�?�            �m@������������������������       ��J�j�?^            �c@������������������������       �q=
ף��?3             T@"       )                   �1@�o}e�?;            @#       (                    @��OC��?0            �T@$       %                    �?     ��?&             P@������������������������       ��p=
ף�?             4@&       '                    �?��J���?             F@������������������������       ��q-�?             *@������������������������       �In�.P��?             ?@������������������������       ���Hx��?
             2@*       1                   �9@��k����?            z@+       .                    �?ĺ��z�?�            �u@,       -                   �2@�|v*���?D            @\@������������������������       ��p=
ף�?             4@������������������������       �u{����?9            @W@/       0                    @��{A���?�             m@������������������������       ����9��?y            �g@������������������������       �=;n,��?             F@2       3                    �?���&��?3            �Q@������������������������       �����>4�?	             ,@4       5                   �?@�Cc}h�?*             L@������������������������       �zk&{��?$            �H@������������������������       �4և����?             @7       J                   �5@�ˇW	�?W           ��@8       A                   �0@}�J��%�?�           (�@9       >                    @c�����?5            �S@:       ;                    �?F#߼��?'             N@������������������������       �������?             &@<       =                    �?�CkR��?            �H@������������������������       �9��8���?             8@������������������������       �^K�=��?             9@?       @                    @�)O�?             2@������������������������       �����X�?             @������������������������       ��zv��?             &@B       I                    @�L	Ƃ?�?�           ��@C       F                   �1@��˙?�?|           `�@D       E                    �?#���HJ�?�            `k@������������������������       �t�û��?             7@������������������������       �cC�B��?w            �h@G       H                    �?�7RM6h�?�           ��@������������������������       ��o��`�?�            �t@������������������������       ��n���?&           �|@������������������������       �     ��?
             0@K       Z                    �?\�2����?�           T�@L       S                    �?��rЛ�?d           ��@M       P                   �<@bB�Fv6�?}             i@N       O                     �?�t ����?d            �d@������������������������       ��Uzo ��?4            �U@������������������������       �P7����?0            @S@Q       R                    �?@�|���?            �B@������������������������       �ffffff�?             $@������������������������       �%�R�@��?             ;@T       W                   �@@�����?�            �v@U       V                    �?�3d`�?�            �t@������������������������       �_j�����?+             S@������������������������       ��M�S�?�            �o@X       Y                    @     P�?             @@������������������������       �"P7��?
             3@������������������������       ���1G���?             *@[       b                   �9@�F̶�<�?8            ~@\       _                    @B{	�%��?�             r@]       ^                   �7@�fXf�Z�?�            �j@������������������������       ��)�/�?P            @^@������������������������       ��v����?6            �V@`       a                    @����U�?:             S@������������������������       ����u���?(             K@������������������������       ���.���?             6@c       f                    @JL<�Z�?x            @h@d       e                     @(��ʼ�?N            �_@������������������������       �F�V15�?<            @X@������������������������       � �^�@��?             =@g       h                     @�}2��?*             Q@������������������������       �k�y�ʍ�?             G@������������������������       ��#��Z=�?             6@�t�bh�h4h7K ��h9��R�(KKiKK��h��BX>       �z@     �U@     Pu@      C@     @S@      C@     @T@     �@     0�@      M@     �V@      e@     ��@     p|@      0@      O@      E@     �_@     �L@     �g@      =@      `@      @      4@      $@      A@     �t@     �t@      &@     �A@      N@     �r@      g@      �?      4@      *@      J@      *@      a@      5@     �U@       @      (@              9@     �p@     �p@       @      ;@      E@     `i@     @_@              "@      @      ?@      $@      I@      &@      ;@      �?      @              "@      P@      X@      �?      @      5@     �R@     �L@              @      �?      0@      @      5@              &@                               @      ;@      G@      �?      @      *@      8@      5@                      �?                      $@              @                                      6@      @               @      �?       @       @                                              @              �?                                      @       @               @               @                                                      @              @                                      .@      @                      �?               @                                              &@              @                               @      @     �D@      �?       @      (@      6@      3@                      �?                      @              @                              �?      @      6@               @      $@      5@      ,@                                              @                                              �?      �?      3@      �?               @      �?      @                      �?                      =@      &@      0@      �?      @              @     �B@      I@              @       @     �I@      B@              @              0@      @      @      @       @                                      �?      @                      �?      1@      "@              �?              @      �?      @                                                      �?                              �?      &@                                                              @       @                                              @                              @      "@              �?              @      �?      8@       @      ,@      �?      @              @      B@      G@              @      @      A@      ;@              @              *@      @      �?       @      �?                                               @                                                                      @              7@      @      *@      �?      @              @      B@      F@              @      @      A@      ;@              @              "@      @     �U@      $@      N@      �?      "@              0@      i@      e@      @      4@      5@      `@      Q@              @      @      .@      @     �B@      @     �@@              @              @     �G@      K@      @      *@      $@      G@     �@@              @              @      @      =@      @      ?@              @              @     �F@     �J@      @      *@      $@     �D@      ?@              @              @      @      $@              @                              �?      A@     �B@      �?               @      2@      &@              �?              @              3@      @      <@              @              @      &@      0@       @      *@       @      7@      4@               @              �?      @       @               @               @                       @      �?                              @       @                              �?              @              �?               @                              �?                               @       @                                              @              �?                                       @                                      @                                      �?              I@      @      ;@      �?       @              $@      c@     �\@      @      @      &@     �T@     �A@              �?      @       @      �?      =@       @      "@                              @     �Z@      J@      @               @     �H@      1@                              @              "@      �?      @                                      N@      9@                              5@      @                                              4@      �?      @                              @     �G@      ;@      @               @      <@      (@                              @              5@      @      2@      �?       @              @      G@     �O@      �?      @      "@     �@@      2@              �?      @      @      �?      @      �?      &@              �?              @     �@@     �G@      �?      @      @      :@      &@                      @      @              ,@       @      @      �?      �?                      *@      0@              @      @      @      @              �?               @      �?     �J@       @      E@      @       @      $@      "@     �P@     �P@      @       @      2@     @X@      N@      �?      &@      "@      5@      @      3@               @                                      5@      ,@       @              �?      6@      �?                                              0@              �?                                      (@      &@       @              �?      4@      �?                                               @                                                      @      @       @              �?      @                                                      ,@              �?                                      @       @                              .@      �?                                              @                                                       @      �?                              @                                                      @              �?                                      @      @                              (@      �?                                              @              �?                                      "@      @                               @                                                      A@       @      D@      @       @      $@      "@      G@     �J@      �?       @      1@     �R@     �M@      �?      &@      "@      5@      @      9@       @      >@      �?      @      $@       @      G@      I@      �?      @      .@     �L@     �J@              @      @      4@       @      ,@      �?       @              @      @              $@      (@                              6@      9@              �?              (@              @      �?      @                                                                              �?      @                              @              &@              @              @      @              $@      (@                              5@      5@              �?              @              &@      �?      6@      �?      @      @       @      B@      C@      �?      @      .@     �A@      <@              @      @       @       @      &@      �?      5@      �?      @      @      @      ?@      @@              @      ,@      8@      1@              @      @      @       @                      �?                              @      @      @      �?              �?      &@      &@              �?              @              "@      @      $@       @      �?              �?              @               @       @      2@      @      �?      @      @      �?      �?       @              �?                              �?                                              @       @                                      �?      @      @      "@       @      �?                              @               @       @      &@      @      �?      @      @      �?              @      @      "@       @                                      @                       @      &@      @               @       @      �?                                              �?                                               @                              �?       @      �?                     `m@      M@     �j@     �@@     �L@      <@     �G@     @j@     @o@     �G@     �K@     @[@     �t@     �p@      .@      E@      =@     �R@      F@     �b@      $@     �V@      &@      .@       @      2@     `d@     `d@      (@      3@      E@     @h@     �a@              2@      @      <@      4@      0@      �?      �?                                      ;@      *@                       @      (@      @                                              *@      �?      �?                                      6@      @                       @      &@      @                                              @      �?                                              �?                                      @                                                      @              �?                                      5@      @                       @       @      @                                              @                                                       @      @                              @      �?                                                              �?                                      *@       @                       @      @      @                                              @                                                      @      @                              �?       @                                                                                                       @      @                                                                                      @                                                      @       @                              �?       @                                             �`@      "@     �V@      &@      .@       @      2@      a@     �b@      (@      3@      D@     �f@     �`@              2@      @      <@      4@     ``@      "@     �V@      &@      .@       @      2@     �`@     �b@      (@      3@      D@     `f@     �_@              2@      @      <@      1@      <@      �?       @              @               @     �B@     �C@      �?      "@      @     �I@      7@              �?      �?      @      �?      @                                                       @      @      �?               @      @      �?                              @              6@      �?       @              @               @     �A@      B@              "@      @     �G@      6@              �?      �?      @      �?     �Y@       @     �T@      &@      &@       @      0@     �X@     �[@      &@      $@      A@      `@     �Y@              1@      @      5@      0@     �C@       @      G@       @      @       @       @      *@     �A@       @      @      6@     �K@      L@              @              1@      @      P@      @      B@      "@      @               @     @U@      S@      @      @      (@     @R@     �G@              $@      @      @      &@      �?                                                      �?                                      @       @                                      @     �U@      H@     @^@      6@      E@      :@      =@     �G@     �U@     �A@      B@     �P@     �`@     @`@      .@      8@      9@      G@      8@     �E@      4@     �R@      &@      ;@      2@      0@      ,@      @@      3@      8@     �F@     �N@     @Q@      "@      1@      2@      9@      4@      8@      @      3@               @              @      "@      (@      @      @      $@     �@@      8@              @      $@      *@       @      7@      @      .@              @              �?       @       @      @      @      @     �@@      6@              @      @      "@      @      "@       @      @              @              �?      @      @               @      @      9@      &@              @       @      @      �?      ,@      �?      "@              @                      @      @      @      @               @      &@              �?      @      @      @      �?      @      @              �?              @      �?      @              �?      @               @              �?      @      @       @                                                      @              @              �?                       @                                              �?      @      @              �?               @      �?      �?                      @                              �?      @      @       @      3@      ,@      L@      &@      3@      2@      "@      @      4@      ,@      2@     �A@      <@     �F@      "@      $@       @      (@      (@      3@      ,@     �K@      $@      0@      2@      "@      @      3@      ,@      0@      8@      <@     �F@      �?      $@      @      (@      "@       @      @      0@      @      @       @              @      @       @              @      "@      @                      �?      @      @      &@      $@     �C@      @      *@      0@      "@       @      0@      (@      0@      1@      3@      D@      �?      $@      @      @      @                      �?      �?      @                              �?               @      &@                       @               @              @                      �?              @                                               @      @                      @               @               @                              �?                                      �?                      @                      @                              �?      F@      <@      G@      &@      .@       @      *@     �@@     �K@      0@      (@      6@     @R@     �N@      @      @      @      5@      @     �@@      .@      =@      "@      @               @      4@     �F@      @      $@      &@      K@      :@      @      @      @      $@              6@      (@      4@      @      �?               @      2@      E@      @      $@      "@     �B@      2@       @                      @              3@      @      "@              �?              @      .@      .@      @       @      @      6@      0@                              @              @      @      &@      @                      @      @      ;@               @      @      .@       @       @                                      &@      @      "@      @      @                       @      @                       @      1@       @      @      @      @      @              &@       @      @      @      �?                      �?      @                              (@      @      �?       @       @      @                      �?      @               @                      �?                               @      @      @       @      �?      �?                      &@      *@      1@       @      &@       @      @      *@      $@      *@       @      &@      3@     �A@      �?      @      @      &@      @       @      @      @       @      &@      @      �?      (@      @      "@       @      @      ,@      9@      �?      @      @      @       @      @      @      @       @      "@      @              &@      @      @       @      @      ,@      ,@               @      @      @       @      �?      �?                       @              �?      �?      @       @                              &@      �?       @              @              @      "@      (@                       @      @      �?      @      @               @      @      $@                      �?      @       @      @      @      (@                              �?      �?       @      @              @      �?       @                      �?       @       @              @                               @      @              �?                      @      @       @                               @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��ahG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKwhnh4h7K ��h9��R�(KKw��hu�B         >                    �?�l`����?�	           ��@                          �1@M�-��?K           ��@                           @q�F�:�?�            @q@                           �?��&k��?H             ]@                          �0@�R�����?             �H@                            �?r�q��?             8@������������������������       �$߼�x�?             .@������������������������       �VUUUUU�?             "@	       
                    �?J+��?             9@������������������������       ��(\����?             $@������������������������       �
ףp=
�?             .@                            �?/��R��?(            �P@                           @�s����?             5@������������������������       ���8��8�?             (@������������������������       ���E���?             "@                           �?������?             G@������������������������       �?4և���?             <@������������������������       �����H�?
             2@                           @p=
ף��?o             d@                            �?�m۶m[�?Q             \@                           @0�����?             5@������������������������       ����!pc�?             &@������������������������       ����Q��?             $@                           @,c8�C�?C            �V@������������������������       �n۶m۶�?(             L@������������������������       ���P���?            �A@                          �0@�������?             H@������������������������       ����Q��?             $@                            �?6��P^C�?             C@������������������������       �1�G�2��?             ;@������������������������       ���!pc�?             &@        /                     �?1���E�?�           ��@!       (                    @L$e?�:�?�             w@"       %                    �?|��{`�?�            �q@#       $                   �;@�]�N��?2            @U@������������������������       �FmW7@��?,            �R@������������������������       ���Q��?             $@&       '                   �5@�Q�|�?w             i@������������������������       �=�ܻb�?7            �V@������������������������       ������?@            �[@)       ,                   �6@C�`PI�?;            �T@*       +                   �4@d�_p�<�?%             K@������������������������       �     ��?             @@������������������������       ��4_�g�?             6@-       .                   �9@�(�I�8�?             =@������������������������       ��.�s�?             3@������������������������       ���(\���?             $@0       7                    @�t4��.�?�           �@1       4                    @;�Kۄ�?�           @�@2       3                    �?���ғ�?�           ��@������������������������       �e�o�W�?�            pq@������������������������       �g'�R��?           Pz@5       6                    @.�I�w��?5             S@������������������������       �     ��?-             P@������������������������       ��q�q�?             (@8       ;                    @]/��P��?�             s@9       :                     �?��"e���?             B@������������������������       �VUUUUU�?             "@������������������������       �rJ�:��?             ;@<       =                    �?���y���?�            �p@������������������������       ����!pc�?4             V@������������������������       �6nK8��?v            �f@?       Z                    �?�������?E           �@@       O                   �9@>;K��?�           ��@A       H                   �2@���W�?W           X�@B       E                    @�o��x��?w            @h@C       D                     �?O��:�?S            @a@������������������������       �:&5�-�?            �D@������������������������       ��^�X�?;            @X@F       G                     �?��>4և�?$             L@������������������������       �V4�ͫ�?             >@������������������������       ��HPS!��?             :@I       L                   �7@3+2m�?�            �v@J       K                     @�I��Z�?�            Pr@������������������������       ���g����?�             k@������������������������       ���(��V�?4            @S@M       N                     �?1�!���?'             Q@������������������������       �     ��?	             0@������������������������       ��.y0���?             J@P       U                   �;@B���J�?=            @Y@Q       T                    @��;�\`�?             E@R       S                   �:@$I�$I��?             <@������������������������       ���>4և�?             ,@������������������������       ��Cc}�?
             ,@������������������������       �I�$I�$�?	             ,@V       Y                    @:���W�?$            �M@W       X                   �=@�46<�?             I@������������������������       ��F���H�?             5@������������������������       �e�$O�?             =@������������������������       ���E���?             "@[       h                   �3@^\�"��?�           �@\       c                    @U�z�  �?6           h�@]       `                     @��
Ŋ�?�            �u@^       _                   �2@������?y             j@������������������������       ����P��?Q            �a@������������������������       �U��5m�?(            �P@a       b                    @�Нq,�?P            @a@������������������������       ��\5ݓ�?(            �P@������������������������       �F��ӭ��?(             R@d       e                    �?��̦G��?m            @f@������������������������       �      �?             0@f       g                   �0@���}�?b            @d@������������������������       ��6�i��?             >@������������������������       �>v�禺�?P            �`@i       p                   �>@ʶc��1�?{           p�@j       m                   �9@ᰐo�?D           ��@k       l                     @ʨ�|��?�           ��@������������������������       �u��h)��?           `|@������������������������       ��.k���?�            �i@n       o                    @����*�?�            Pp@������������������������       ���(��?�            �k@������������������������       �{�G�z�?             D@q       t                     �?�n��i�?7            �U@r       s                   �?@�]�"R�?            �C@������������������������       �h/�����?             "@������������������������       ���2Tv�?             >@u       v                     @UUUUU��?!             H@������������������������       �r�q��?	             (@������������������������       �O��E��?             B@�t�bh�h4h7K ��h9��R�(KKwKK��h��B�F       p|@     �U@     `t@      C@     �T@      ;@     �S@     X�@     ��@     �Q@     @S@     �f@     ��@      {@      @     �U@      B@     �`@      C@     �k@      ;@     �^@      @      @@      @      8@     �s@     pr@      0@     �B@     �L@     `r@      d@      �?      ?@      *@      J@      ,@      D@       @      "@                              �?     �[@      M@      @       @      @     �B@      @                              �?              9@               @                                      >@      5@      @       @       @      :@      @                              �?              1@              �?                                      $@      $@      �?       @       @      @                                                      "@              �?                                      @      @               @              �?                                                      @              �?                                      �?      @               @                                                                      @                                                      @      �?                              �?                                                       @                                                      @      @      �?               @      @                                                      @                                                       @       @      �?               @                                                              @                                                      @       @                              @                                                       @              �?                                      4@      &@       @                      4@      @                              �?                                                                      $@       @                               @                                      �?                                                                      @      �?                              @                                                                                                              @      �?                               @                                      �?               @              �?                                      $@      "@       @                      (@      @                                              @              �?                                      "@      @                              @      @                                              @                                                      �?      @       @                      @                                                      .@       @      @                              �?     @T@     �B@                      @      &@      @                                              @       @      @                              �?     @P@      9@                      �?      @      �?                                                              �?                                      .@      @                      �?                                                                                                                       @      @                                                                                                      �?                                      @      �?                      �?                                                              @       @      @                              �?      I@      5@                              @      �?                                               @       @      �?                              �?      A@      $@                              @                                                      @              @                                      0@      &@                              �?      �?                                              $@               @                                      0@      (@                       @      @       @                                              �?                                                      @      �?                              �?                                                      "@               @                                      "@      &@                       @      @       @                                              @                                                      @      &@                       @      @      �?                                              @               @                                       @                                              �?                                             �f@      9@     �\@      @      @@      @      7@      j@     �m@      *@     �A@      J@     p@     @c@      �?      ?@      *@     �I@      ,@      I@      (@      9@       @      @              @      ;@     @P@      @      *@      .@     �Q@      D@              @      �?      8@      @     �E@      "@      1@       @      @              @      1@     �G@              (@      (@      O@      5@              @      �?      8@      @      2@              @       @      �?              @       @      5@              @      @      7@      @                      �?                      *@              @       @      �?              �?       @      3@              @       @      7@      @                      �?                      @                                               @               @                      �?                                                              9@      "@      ,@               @                      .@      :@              "@      "@     �C@      0@              @              8@      @      3@       @      @              �?                      &@      &@               @       @      5@       @               @              @      @      @      @      &@              �?                      @      .@              @      �?      2@      ,@              @              5@      �?      @      @       @                                      $@      2@      @      �?      @      "@      3@              �?                              @      @      @                                       @      .@       @      �?       @      @      @              �?                              @      @      @                                       @      @       @                      @      @              �?                               @                                                      @      "@              �?       @       @                                                       @              �?                                       @      @       @              �?      @      .@                                              �?              �?                                       @       @                              @      $@                                              �?                                                              �?       @              �?              @                                             @`@      *@     @V@      @      =@      @      4@     �f@     �e@      "@      6@     �B@     @g@     �\@      �?      8@      (@      ;@       @     @Z@      "@     �R@      @      <@      @      3@     �Z@      Z@      @      0@      ?@     @`@      T@      �?      2@      (@      6@      @     �W@      "@      M@      @      9@      @      3@      V@     �X@      @      ,@      ?@      ^@      R@      �?      2@      (@      6@      @     �G@      @      6@              &@              @      7@      C@       @      "@      @     �I@      @@      �?      $@              ,@      �?     �G@      @      B@      @      ,@      @      *@     @P@      N@       @      @      9@     @Q@      D@               @      (@       @      @      &@              1@              @                      2@      @      �?       @              $@       @                                              &@              1@                                      0@      @      �?      �?              "@      @                                                                              @                       @                      �?              �?      @                                              9@      @      ,@              �?              �?     �R@      Q@      @      @      @      L@      A@              @              @      �?      @              �?                                      6@       @                              @      @                                              @              �?                                      @                                              �?                                                                                                      2@       @                              @      @                                              6@      @      *@              �?              �?     �J@     �P@      @      @      @      J@      >@              @              @      �?      *@               @                                      "@      <@              �?       @      3@      ,@                                              "@      @      &@              �?              �?      F@      C@      @      @      @     �@@      0@              @              @      �?     `m@     �M@     `i@     �@@     �I@      6@     �K@     �m@     pq@     �K@      D@     �_@     �t@     q@      @      L@      7@     @T@      8@     �R@      (@      C@      @      4@       @      0@     �W@      ]@      3@      ,@      :@     �V@     �S@              (@      @      2@      @     �Q@      "@     �@@      @      "@      @      (@     �W@     �[@      (@      @      1@     �S@     �M@              (@      @      (@      @      5@      �?      (@              �?              @     �H@      C@       @      @      �?     �C@      .@                              @       @      2@      �?      &@              �?              @      8@      <@       @      @              ?@      $@                              @       @       @                                                      @      ,@              �?              *@      @                              @              0@      �?      &@              �?              @      4@      ,@       @       @              2@      @                                       @      @              �?                               @      9@      $@                      �?       @      @                              �?              @                                               @       @      "@                      �?      @      @                              �?                              �?                                      1@      �?                              @       @                                             �H@       @      5@      @       @      @      @     �F@     @R@      $@      @      0@      D@      F@              (@      @      @      @      F@      @      0@      @       @      @       @      E@     �L@      @      @      .@      :@      B@              (@      @      @      @      A@       @      ,@               @      �?       @     �C@      G@               @      $@      3@      <@               @       @      @      �?      $@       @       @      @      @      @              @      &@      @      �?      @      @       @              @      @      �?       @      @      @      @                      �?      @      @      0@      @      �?      �?      ,@       @                                                               @                               @       @      @      �?                      @                                                      @      @      @                      �?      @      �?      *@      @      �?      �?       @       @                                              @      @      @      @      &@       @      @      �?      @      @      @      "@      (@      3@                      �?      @       @       @       @       @       @      @                      �?               @              @      $@      (@                                               @              �?       @      �?                                      �?              @      "@      "@                                              �?              �?       @                                                                      @      @                                              �?                              �?                                      �?              @      @      @                                                       @      �?              @                      �?              �?                      �?      @                                               @      �?      @      �?      @       @      @              @      @      @      @       @      @                      �?      @       @       @              @      �?      @       @      @              @      @      @      @       @       @                      �?      @       @                       @               @              @              @      �?      @                      �?                              �?       @       @              �?      �?      @       @                              @       @      @       @      �?                      �?      @                      �?                                                       @                                      @                              �?              d@     �G@     �d@      ;@      ?@      ,@     �C@     �a@     `d@      B@      :@      Y@      n@     `h@      @      F@      1@     �O@      1@     �R@       @      K@      @      @              @     @V@     @U@      @      @      2@     �T@     �K@               @      @      4@      @     �G@      @     �E@      @      @              @      C@      J@      @      @      (@      O@      G@              @       @      .@      @      ;@       @      ;@       @       @              @      ;@     �A@      �?               @      F@      3@              @      �?      @      @      ,@      �?      4@                              @      5@      5@      �?              @     �C@      ,@                      �?       @              *@      �?      @       @       @                      @      ,@                      @      @      @              @              @      @      4@      @      0@       @      @                      &@      1@       @      @      @      2@      ;@                      �?      $@              @      @      (@      �?      @                      @      "@               @              .@      @                              �?              ,@              @      �?                              @       @       @      �?      @      @      4@                      �?      "@              ;@       @      &@       @                             �I@     �@@       @      @      @      5@      "@              @      �?      @              &@      �?                                              �?                                      �?       @                                              0@      �?      &@       @                              I@     �@@       @      @      @      4@      @              @      �?      @              @              �?                                      ,@      �?                              @      �?                               @              $@      �?      $@       @                              B@      @@       @      @      @      .@      @              @      �?      @             �U@     �C@     �[@      5@      :@      ,@      B@      J@     �S@      ?@      4@     �T@     �c@     �a@      @      B@      ,@     �E@      ,@      U@      B@     �W@      0@      7@      "@      B@      J@     �R@      :@      0@      O@     �c@      a@       @     �@@      $@     �D@      (@     @R@      7@     �R@      "@      0@      @      4@      D@     �M@      3@      .@      F@      ]@     �V@      �?      ,@      @      ?@      @      I@      0@     �K@      @      *@      �?      "@      @@      E@      ,@      ,@      =@      U@     �E@              (@      @      ;@      @      7@      @      3@       @      @      @      &@       @      1@      @      �?      .@      @@      H@      �?       @       @      @      �?      &@      *@      5@      @      @      @      0@      (@      .@      @      �?      2@      D@     �F@      �?      3@      @      $@       @      @      $@      *@      @      @      @      *@      (@      .@      @      �?      2@      B@     �D@      �?      3@      �?      @      @      @      @       @       @                      @                      @                      @      @                      @      @      �?      @      @      0@      @      @      @                      @      @      @      4@      �?      @      @      @      @       @       @      @              @      @       @                               @      �?              1@      �?                              �?       @                              @                                                                      @                                      �?                      @               @      @       @                               @      �?              *@      �?                                       @                      @      $@      �?      �?      @                       @      @      @      @              @      @      @      @               @               @      @              �?                              �?      �?                              �?                       @                              �?      @      �?              @                      �?      @      @      @              @      @      @      �?               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�L�|hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKmhnh4h7K ��h9��R�(KKm��hu�B�         8                   �4@"B�GG��?�	           ��@                            @�t��'M�?o           T�@                            �?�~��T��?!           �@                           �?��|p�/�?J           x�@                          �1@�9��9��?�            �q@                           @_ޛ�T��?@            @Y@������������������������       �v_����?3            �T@������������������������       ��KM�]�?             3@	       
                    �?o
Z.��?q            @g@������������������������       �)\�����?6             T@������������������������       ��b-����?;            �Z@                           @yÏ��?�           ��@                           @�_m�WT�?	           pz@������������������������       �ʀ1d��?�            �u@������������������������       �^U�'"��?5            @R@                            �?���!<0�?�             m@������������������������       �
^N��)�?F             \@������������������������       ���'d��?J            @^@                           @bW��"?�?�            pu@                           @�Q�}e��?�             j@                           @�C"�b��?r            �d@������������������������       ��*9�b��?5            @S@������������������������       �d��K|��?=            �U@                           �?(&ޏ��?             F@������������������������       �        	             7@������������������������       ���kv�?
             5@                          �3@|2֟3�?R            �`@                          �2@��ϭ�*�?G             ]@������������������������       ���a�2�?2            �T@������������������������       �%�Էr�?            �@@������������������������       ��}�+r��?             3@        )                   �0@���;��?N           x�@!       $                    �?�Qk�?'            �L@"       #                    @��WV��?             :@������������������������       ��X�C�?
             ,@������������������������       �9��8���?	             (@%       &                    �?p��N�?             ?@������������������������       ���!pc�?             &@'       (                    @�Q����?             4@������������������������       �r�q��?             (@������������������������       �      �?              @*       1                    �?	������?'           `}@+       .                    @����r��?y            @g@,       -                    @CG�:�?_            �b@������������������������       �M�h���?A             Z@������������������������       ������?            �G@/       0                   �2@p�_�Q�?            �A@������������������������       �lv�"��?             5@������������������������       ��>4և��?             ,@2       5                    @�&���?�            �q@3       4                   �1@0	>.r�?�            �m@������������������������       �/ 6����?,            �Q@������������������������       �j��6���?l             e@6       7                    @ڤ�:�^�?            �F@������������������������       �r�q��?             (@������������������������       ��B#�E�?            �@@9       T                     @]
Zi�?#           h�@:       I                   �<@�7����?�           ��@;       B                    �?�d����?           l�@<       ?                    @A���'��?b           X�@=       >                    @���'�%�?           @{@������������������������       ���<�!�?�            �y@������������������������       �^�:|z�?
             5@@       A                    @���t�9�?\            �b@������������������������       �P(�y#�?*            �O@������������������������       �n,�Ra�?2             V@C       F                   �5@SI\6���?�           ��@D       E                    �?���� �?_            �a@������������������������       �������?"            �J@������������������������       �D����0�?=            �U@G       H                    �?��0"��?]            �@������������������������       �     ��?�             p@������������������������       �`��rB��?�            @t@J       Q                    @_E�|�?�            �i@K       N                    �?Ri�D�?s             f@L       M                    �?�|��0��?)            @Q@������������������������       ��o^M<+�?             .@������������������������       �l����?"             K@O       P                   �>@�S����?J             [@������������������������       ����ߎD�?#            �H@������������������������       �KHݒ��?'            �M@R       S                   �@@4և����?             <@������������������������       �     ��?             0@������������������������       �r�q��?	             (@U       ^                    �?<�M`gZ�?{           `�@V       ]                    @��'c�	�?D            �Z@W       Z                   �8@p�N�-�?:            @U@X       Y                    �? �$D4�?"            �G@������������������������       ��ܤ��?             5@������������������������       ���?�(�?             :@[       \                   �:@� u#��?             C@������������������������       �:���I�?             1@������������������������       �wKnR�?             5@������������������������       �lv�"��?
             5@_       f                   �<@ѺO7[I�?7            ~@`       c                    �?���{���?            y@a       b                    @W���N��?t            `g@������������������������       ��k�΋��?S             `@������������������������       ���Bb��?!             M@d       e                    �?aG.��?�            �j@������������������������       �LU��$�?             �H@������������������������       �-���@L�?n            �d@g       j                   �>@     ��?5             T@h       i                    �?�Rͦ$�?            �B@������������������������       �ܶm۶m�?             5@������������������������       �      �?             0@k       l                   �@@J1|w���?            �E@������������������������       �6�;Nё�?             9@������������������������       �~X�<��?             2@�t�bh�h4h7K ��h9��R�(KKmKK��h��B�@       p}@      Q@      t@      4@     �O@      ?@     �U@     ��@     ��@      R@     @V@      f@     ؃@      z@      "@     �Q@      I@     @\@     �L@     �m@      &@      ^@              *@      �?      7@     z@     �t@      0@      ;@     �Q@     �s@     �a@              5@       @      J@      &@      e@      @     �P@              @              .@     Pu@     `o@      &@      3@     �J@     `i@      W@              (@      @     �@@      @     @a@      @     �E@              �?              &@     �j@     �f@      @      3@     �G@     @d@     �P@              &@      @      :@      @     �J@      �?      2@              �?              @      J@     �B@      @      &@      .@     �K@      7@               @              $@      @      1@              @                              �?      =@      *@       @      @      @      2@      @                              @              1@              @                              �?      6@       @              @      @      .@      @                              @                                                                      @      @       @              �?      @      �?                                              B@      �?      .@              �?               @      7@      8@      �?      @      "@     �B@      2@               @              @      @      1@      �?      �?              �?                      *@      $@      �?      @       @      5@       @               @                       @      3@              ,@                               @      $@      ,@                      @      0@      0@                              @      �?     @U@      @      9@                               @     `d@     �a@      @       @      @@     �Z@     �E@              "@      @      0@      @     �G@       @      *@                              @     @^@      U@              @      .@     �S@      ?@              @      �?      "@      @     �A@      �?      $@                              @     �Z@     �R@              @      &@     �P@      9@               @              @      @      (@      �?      @                              @      ,@      $@                      @      (@      @              @      �?      @              C@      �?      (@                              �?      E@     �M@      @       @      1@      <@      (@              @      @      @      �?      0@      �?      @                              �?      3@     �B@      @              @      ,@      @                       @      @              6@               @                                      7@      6@               @      *@      ,@      @              @      @      @      �?      >@       @      7@               @              @     �_@     �Q@      @              @     �D@      :@              �?              @              ,@              *@               @              @     @U@      ?@      @               @      ;@      7@                              @              ,@              *@               @              @     �K@      <@      @               @      :@      *@                              @               @              @               @              @      8@      (@                       @      @      @                              @              @              @                                      ?@      0@      @                      3@      @                                                                                                      >@      @                              �?      $@                                                                                                      7@                                                                                                                                                      @      @                              �?      $@                                              0@       @      $@                                     �D@      D@      �?              @      ,@      @              �?              @              "@              @                                     �C@      C@      �?              @      *@      @                               @              @              @                                      :@     �@@                      @      @       @                                               @               @                                      *@      @      �?                      @      �?                               @              @       @      @                                       @       @                              �?                      �?              �?              Q@      @      K@              $@      �?       @      S@     �S@      @       @      1@     �\@     �H@              "@       @      3@      @      *@              @               @                      3@      &@                              @      @                                              @                                                      $@      @                              @      �?                                              @                                                       @      �?                               @                                                      @                                                       @      @                              @      �?                                              @              @               @                      "@      @                                      @                                               @                                                      @       @                                      �?                                              @              @               @                      @      @                                       @                                              @               @                                              @                                      �?                                                              �?               @                      @      �?                                      �?                                             �K@      @     �I@               @      �?       @     �L@     �P@      @       @      1@     @[@     �F@              "@       @      3@      @      1@      �?      8@                      �?       @      B@      :@       @       @      @      A@      6@              @               @      �?      *@      �?      2@                      �?      �?      A@      3@                      @      ?@      3@               @              @      �?       @      �?      ,@                      �?      �?      0@      &@                      @      9@      *@               @              @      �?      @              @                                      2@       @                              @      @                                              @              @                              �?       @      @       @       @       @      @      @              �?               @              @              @                                       @      @       @                       @                      �?                                              @                              �?                               @       @      �?      @                               @              C@      @      ;@               @              @      5@     �D@      @      @      $@     �R@      7@              @       @      &@      @      @@      @      ;@               @               @      0@      >@      @      @      @     �P@      5@               @       @      $@       @      ,@              @               @                      (@      @               @       @      *@      @              �?              @              2@      @      4@              @               @      @      8@      @      @      @      K@      ,@              �?       @      @       @      @                                              @      @      &@                      @       @       @              @              �?      �?       @                                              �?      @       @                      @                                                      �?      @                                              @       @      "@                               @       @              @              �?             `m@     �L@     @i@      4@      I@      >@     �O@     �b@     �p@      L@      O@     �Z@     �s@     0q@      "@      I@      E@     �N@      G@     @g@     �C@     �c@      $@      B@       @     �E@      \@     �j@     �E@     �I@     �O@     `n@     �f@      @      =@      9@     �F@      9@     �d@      A@     �_@      "@      7@      @      A@     �[@     �h@      >@      F@     �F@     `l@     @d@       @      5@      0@      C@      1@     �R@      (@      N@      @      @              ,@     �N@      ]@      @      1@      1@     �Y@     @R@              @      @      $@      @      M@      &@     �M@      �?      @              ,@      E@     �P@      @      "@      (@     �R@      N@              @      @       @       @     �L@      &@      L@      �?      @              ,@      ?@     �P@      @      "@      (@     �Q@      M@              @      @       @       @      �?              @                                      &@      �?                              @       @                                              1@      �?      �?       @       @                      3@     �H@               @      @      <@      *@                       @       @       @      (@      �?                                              &@      0@              �?              $@      $@                       @                      @              �?       @       @                       @     �@@              @      @      2@      @                               @       @     �V@      6@     �P@      @      0@      @      4@      I@     �T@      7@      ;@      <@     @_@     @V@       @      1@      &@      <@      *@      7@      �?       @                              "@      1@      =@              @      @      *@      3@                              @      @      @                                              @      @      3@               @       @       @      "@                               @       @      2@      �?       @                              @      &@      $@               @      @      &@      $@                              @      @     �P@      5@     �M@      @      0@      @      &@     �@@     �J@      7@      7@      6@      \@     �Q@       @      1@      &@      6@       @      A@      (@      ;@      �?      $@       @       @      @      "@      (@      0@      *@      J@      ?@      �?      $@      @      "@      @     �@@      "@      @@      @      @       @      "@      =@      F@      &@      @      "@      N@     �C@      �?      @      @      *@       @      5@      @      ?@      �?      *@      @      "@      �?      .@      *@      @      2@      0@      2@      �?       @      "@      @       @      2@      @      ?@      �?      *@      @      @              *@      (@      @      0@      .@      *@      �?      @       @      @      @      "@      @      &@              "@              �?               @      @      @      �?       @      @                      �?              @                      @              @                               @      @                      �?      �?                                      �?      "@      @      @              @              �?              @       @      @      �?      @      @                      �?              @      "@       @      4@      �?      @      @      @              @      @      @      .@      @      @      �?      @      @      @      �?       @      �?      @      �?       @      �?       @              �?       @       @       @      @      @      �?      @      @      @      �?      �?      �?      ,@               @       @       @              @      @      �?      *@      @      �?              @      @      �?              @                                      �?      @      �?       @      �?      �?       @      �?      @              �?      �?       @      @      �?                                      �?      @      �?       @              �?              �?       @              �?      �?       @               @                                              �?                      �?               @              @                                      @     �H@      2@      F@      $@      ,@      6@      4@     �B@      L@      *@      &@     �E@     �R@     �W@      @      5@      1@      0@      5@       @      @      "@              @      �?       @      "@       @      @       @      @      5@      $@              �?      @       @      @      @      @      "@              @      �?      �?      @       @      @       @      @      .@      @              �?      @       @      @      @       @      @               @      �?      �?      @       @      @      �?      @              @              �?      @       @       @              �?      @                      �?              �?      @      @              @              �?              �?       @                      @      �?      �?               @              �?      @      @       @      �?      �?               @                      �?       @       @      �?      �?      @               @                       @              �?      �?      @      .@      @                      @              �?                       @              �?                                                              &@                              @                      �?      �?       @              �?                       @              �?      �?      @      @      @                                      �?      @                                              �?      @                                      @      @                                      @     �D@      .@     �A@      $@      $@      5@      2@      <@      H@      @      "@      B@      K@     @U@      @      4@      &@      ,@      ,@      B@      (@      =@      $@      @      0@      ,@      ;@      G@      @      @      >@      I@     �S@      @       @      "@      &@      @      2@      @      (@      @       @      �?       @      6@      3@       @              ,@      @@     �@@       @      @      @      @       @      *@       @       @      @       @      �?       @      "@      1@                      ,@      0@      :@       @      @      @      @      �?      @       @      @                                      *@       @       @                      0@      @              �?      �?      @      �?      2@       @      1@      @      @      .@      (@      @      ;@      @      @      0@      2@     �F@       @      @      @      @       @       @      @      @      �?      @      @      �?              @      �?              @      @      @              �?      @      �?              0@      @      (@      @       @       @      &@      @      5@       @      @      $@      *@      E@       @      @              @       @      @      @      @              @      @      @      �?       @       @      @      @      @      @       @      (@       @      @      $@      @              @                              @               @                       @      @      @               @              @       @      @              �?                              @                                              @      @               @               @       @      �?              @                                               @                       @      �?                      @              �?              �?      @       @              @      @              �?               @      @      @              @       @      @       @               @      �?      @       @                      @              �?               @      �?      �?              @              �?       @              @                                      @      �?                                       @      @                       @      @                      @�t�bub��e      hhubh)��}�(hhhhhKhKhKhG        hh.hNhJn�ihG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmK{hnh4h7K ��h9��R�(KK{��hu�B�         >                   �2@��o���?�	           ��@                           @ض�����?�           �@                           �?��L��w�?+           �}@                          �1@�Ğ4���?�            pt@                           �?	T�B���?n            �e@                           �?      �?+             R@������������������������       �l~X�<�?             B@������������������������       �l~X�<�?             B@	       
                    �?�_<�l��?C            �Y@������������������������       ��� =[�?             A@������������������������       �C%��N��?,            @Q@                           �?���|�?a             c@                            �?�A�f���?             I@������������������������       �     ��?             0@������������������������       ��@�m�?             A@                           �?�������?C            �Y@������������������������       ��DR���?             G@������������������������       �����S�?$             L@                            �?o����?\            �b@                           �?� _���?&            �O@                          �0@Iє�?             A@������������������������       �H�z�G�?             $@������������������������       ��q�q�?             8@                           @΃�\�?             =@������������������������       ��.�?�P�?             .@������������������������       �����S�?             ,@                           @�z�b��?6            �U@                           �?�d��1��?*            �Q@������������������������       �R~��#��?            �G@������������������������       ���/��@�?             7@������������������������       �     ��?             0@        /                   �0@hz���M�?\           (�@!       (                     �?������?K             _@"       %                    �?�paRC�?)             Q@#       $                    �?ۛ�xt�?            �C@������������������������       �:���I�?             1@������������������������       ��A�0�~�?             6@&       '                    �?c��gS~�?             =@������������������������       ��)x9/�?             ,@������������������������       ��������?	             .@)       ,                     @���X�?"             L@*       +                    @����S��?             <@������������������������       ��������?             (@������������������������       �     ��?
             0@-       .                    @��X��?             <@������������������������       �      �?
             0@������������������������       ��������?             (@0       7                     �?������?           �z@1       4                   �1@'���?P            ``@2       3                    @�5ɬ?�?+            �R@������������������������       ���zv��?             F@������������������������       �k�Y�H��?             >@5       6                    �?\:��?%            �L@������������������������       ��5;j��?             5@������������������������       �~X�<��?             B@8       ;                     @ID~��?�            `r@9       :                    @x|T
�?�            `k@������������������������       �F�h�6�?n             d@������������������������       ��y��*�?              M@<       =                    @hE#߼�?3            �R@������������������������       �      �?%             L@������������������������       ����,�?             3@?       ^                     @����K��?6           ��@@       O                    �?��:�g��?           ��@A       H                    �?^����?G           x�@B       E                    @��,c�?�            �s@C       D                   �4@&Tc^ӝ�?}            �h@������������������������       �������?            �H@������������������������       ��?�|��?`            �b@F       G                    @H�]qb��?G            @]@������������������������       �^���� �?            �D@������������������������       �.窷u�?2             S@I       L                    @�ߍ�}�?�           ��@J       K                    @�M��aD�?�            �q@������������������������       ��/k���?R            �_@������������������������       ��l�o�?f            @c@M       N                   �=@�N��r�?�            �s@������������������������       ��;��;A�?�            �r@������������������������       �*�8�G��?             1@P       W                    �?<�׿0�?�           ��@Q       T                    �?
�-@��?            �{@R       S                    �?rfg�Ka�?t             f@������������������������       �Nb&����?!            �H@������������������������       �     5�?S             `@U       V                     �?����~�?�            �p@������������������������       ��ћ=4��?c            �c@������������������������       ���Au���?I            �Z@X       [                    @�aĳ�?�           8�@Y       Z                    @L?��[�?=           0�@������������������������       ��[r��G�?7           �@������������������������       ��G�z��?             $@\       ]                   �>@��V����?g             d@������������������������       ��������?a            �b@������������������������       �}��7�?             &@_       l                    �?�1�3�'�?+           Ȋ@`       g                    @;�\E^�?�            Pu@a       d                    @KP�H��?�            �p@b       c                   �9@G�I@��?l            �d@������������������������       �P,�Ս��?S            �_@������������������������       ����Q��?             D@e       f                    �?���b� �?E            �Y@������������������������       �h�UF$��?;            �U@������������������������       ��M�]��?
             1@h       i                    �?�2�tk~�?-             R@������������������������       ���ٴ��?             ;@j       k                    @�"����?            �F@������������������������       �؉�؉��?
             *@������������������������       �      �?             @@m       t                    �?,掷dm�?M            �@n       q                    �?��bD}��?�            �u@o       p                    @-�R�C��?<            @X@������������������������       �����>4�?"             L@������������������������       ����p�?            �D@r       s                    �?k�P�N��?�             o@������������������������       ��h70V�?-             O@������������������������       �����^Q�?~            `g@u       x                    @Y�R���?f            @e@v       w                   �<@4�����?I             ]@������������������������       �U$	��$�?A            �X@������������������������       �Iє�?             1@y       z                    @�|ew���?             K@������������������������       �p_�Q�?             9@������������������������       ��V�D.(�?             =@�t�bh�h4h7K ��h9��R�(KK{KK��h��BI       �{@      Q@     �r@      J@     �R@      6@     @T@     p�@     8�@     �R@     @W@      c@     ��@      {@      *@      R@      L@      b@      J@      b@      "@     �J@       @      @              &@     �p@     `j@      @      (@      9@     �b@     �S@               @      @      >@      @      U@      @      ;@       @      @              @     �Q@     @Z@       @      "@      ,@     �S@     �C@              @      @      3@      @      K@      @      3@       @      @              @      D@     �N@       @      @      (@     �O@      ;@              @       @      1@      @     �A@      �?      &@              @              �?      <@      4@       @       @      @      C@      .@              @       @      @      @      (@              @                                      1@      ,@      �?              �?      1@      @                                               @              �?                                      "@      $@      �?              �?      @      �?                                              @              @                                       @      @                              (@      @                                              7@      �?      @              @              �?      &@      @      �?       @      @      5@      "@              @       @      @      @      $@      �?                      @                      @       @                              $@      @                                      �?      *@              @                              �?      @      @      �?       @      @      &@      @              @       @      @       @      3@      @       @       @                      @      (@     �D@              @      @      9@      (@               @              (@      �?      "@      @      �?                                      @      (@                      �?       @      @              �?              $@              �?                                                               @                      �?              @                              @               @      @      �?                                      @      @                               @       @              �?              @              $@              @       @                      @       @      =@              @      @      7@      @              �?               @      �?      @              @                                      @      *@              @      @      "@      @                                      �?      @              @       @                      @      @      0@                              ,@      @              �?               @              >@               @                                      >@      F@              @       @      .@      (@              �?       @       @              @               @                                      ,@      8@              @       @      @      @              �?              �?               @               @                                      &@      &@              @       @       @                                      �?                                                                      �?      @              @                                                                       @               @                                      $@      @                       @       @                                      �?              @                                                      @      *@                              @      @              �?                              @                                                       @      �?                              @      @              �?                                                                                      �?      (@                              �?                                                      8@              @                                      0@      4@                              "@       @                       @      �?              6@              @                                      0@      &@                               @      @                       @                      0@               @                                      &@      $@                              @      @                                              @               @                                      @      �?                              @      @                       @                       @               @                                              "@                              �?      �?                              �?             �N@      @      :@              �?              @      i@     �Z@      @      @      &@      R@     �C@               @      �?      &@              5@               @              �?                     �O@      0@                      �?      (@      @                               @              ,@               @                                      :@      *@                      �?       @       @                               @              @               @                                      2@      $@                              @                                                      �?               @                                      &@                                      @                                                      @                                                      @      $@                                                                                       @                                                       @      @                      �?      @       @                               @              @                                                      @       @                              @                                                      @                                                      @      �?                      �?      �?       @                               @              @                              �?                     �B@      @                              @      @                                               @                                                      5@       @                               @      �?                                                                                                      $@      �?                                      �?                                               @                                                      &@      �?                               @                                                      @                              �?                      0@      �?                               @      @                                              @                              �?                      &@      �?                                                                                       @                                                      @                                       @      @                                              D@      @      8@                              @     @a@     �V@      @      @      $@      N@     �@@               @      �?      "@              (@       @      �?                              @     �A@     �B@               @      @      2@      *@                      �?      @              @              �?                                      >@      5@               @      �?      &@       @                              �?              @                                                      4@      0@               @              �?       @                                               @              �?                                      $@      @                      �?      $@                                      �?              @       @                                      @      @      0@                      @      @      &@                      �?       @                                                              @      �?      @                              @      @                                              @       @                                              @      $@                      @      @      @                      �?       @              <@      �?      7@                              @     �Y@     �J@      @      �?      @      E@      4@               @              @              3@      �?      $@                              @      U@      D@      @              @      ?@      1@               @              @              @      �?      @                              �?      R@      <@      �?               @      >@      (@                                              (@              @                               @      (@      (@      @              �?      �?      @               @              @              "@              *@                              �?      3@      *@              �?      @      &@      @                               @              @              *@                                      0@      @              �?      @       @       @                                               @                                              �?      @      @                              @      �?                               @             �r@     �M@      o@      I@     �Q@      6@     �Q@     �q@     @y@     �P@     @T@     �_@     `|@     @v@      *@      P@     �I@     �\@      H@     �l@     �B@     �f@      <@     �C@       @      I@     @n@     �s@     �F@     �L@     �T@      t@     �k@      @      E@      <@      T@      <@     �Z@      0@      R@      @      "@              5@      `@     @f@      $@      >@      :@      d@     �Y@              &@       @      3@      "@     �E@      @      9@       @      @              @      9@     @V@      �?      (@      *@      K@      ;@              �?      @      @       @      8@      @      &@       @      @              @      @     �P@      �?       @      &@      ?@      ,@              �?      @      @       @      �?              �?                                       @      2@                      @      ,@       @                                              7@      @      $@       @      @              @      @      H@      �?       @      @      1@      @              �?      @      @       @      3@              ,@                                      3@      7@              @       @      7@      *@                                              @              @                                      @      @              @       @      ,@      @                                              .@              $@                                      0@      0@              �?              "@      "@                                             �O@      $@     �G@      @      @              0@      Z@     @V@      "@      2@      *@     �Z@     �R@              $@      @      0@      @      =@      @      7@              @              @      ?@      ;@      @      &@      "@      P@     �C@              @      @      &@      @      $@      @      (@                              @      0@      @      @      @       @      6@      3@              @       @      "@      @      3@      @      &@              @               @      .@      4@      �?       @      �?      E@      4@               @      �?       @      @      A@      @      8@      @       @              "@     @R@      O@      @      @      @      E@      B@              @       @      @      �?      @@      @      5@      @      �?              "@     @R@      O@      @      @      @      D@      <@              @       @      @               @              @              �?                                                               @       @                                      �?     �^@      5@      [@      7@      >@       @      =@     @\@     �`@     �A@      ;@     �L@      d@     �]@      @      ?@      4@     �N@      3@     �H@      *@     �I@      &@      1@      @      ,@      =@      >@      0@      1@      7@     �F@     �L@       @      .@      (@      6@      (@      4@      @      0@              "@      �?      @      "@      0@      @      @      (@      9@      4@              @      @      "@      @      @               @              @              @       @      "@              @       @      @      @              @      �?       @      �?      *@      @      ,@              @      �?      @      @      @      @       @      $@      5@      .@              @       @      @      @      =@      @     �A@      &@       @      @      @      4@      ,@      &@      &@      &@      4@     �B@       @       @      "@      *@      @      4@      @      4@       @      @      @      @      @      &@      @      "@      @      &@      4@       @      @      @      @      @      "@      �?      .@      @      �?               @      .@      @       @       @      @      "@      1@              @      @      @      @     @R@       @     �L@      (@      *@       @      .@      U@      Z@      3@      $@      A@     �\@     �N@       @      0@       @     �C@      @     �J@      @      D@      $@      "@       @      (@     �N@     �X@      .@       @      5@     @X@      D@       @      &@      @      7@      @     �J@      @      D@      @      @       @      &@     �M@     �X@      .@       @      5@      X@      D@       @      &@      @      7@      @                              @       @              �?       @                                      �?                                                      4@       @      1@       @      @              @      7@      @      @       @      *@      2@      5@              @      @      0@       @      4@       @      *@       @      @               @      7@      @      @       @      &@      2@      5@              @      @      (@       @                      @                              �?                                       @                                              @             �R@      6@      Q@      6@      @@      ,@      4@     �F@      W@      6@      8@      F@     �`@      a@      "@      6@      7@      A@      4@      :@       @      =@      @      (@      �?      @      :@      B@      @      *@      &@     @S@      K@       @      "@      &@      "@      @      7@      �?      :@      @      (@      �?      @      3@     �@@      @      "@      &@     �L@     �A@       @      @      &@      @      @      3@              2@      �?      @                      ,@      6@      @      @      @      <@      9@       @      @      @      @       @      (@              @      �?      @                      ,@      6@      @      �?      �?      9@      5@       @      @      @      @              @              (@               @                                              @      @      @      @               @                       @      @      �?       @      @      @      �?      @      @      &@              @      @      =@      $@                      @       @      @      @               @      @      @      �?      @      @      $@              @      @      2@      "@                      @       @      @              �?                                                      �?                      �?      &@      �?                       @                      @      �?      @                              @      @      @      @      @              4@      3@              @               @              �?      �?                                              �?      @                              $@      &@                                               @              @                              @      @              @      @              $@       @              @               @              �?              �?                                      @                      �?              @      �?              �?                              �?               @                              @      @              @      @              @      @              @               @              H@      4@     �C@      2@      4@      *@      *@      3@      L@      0@      &@     �@@     �L@     �T@      @      *@      (@      9@      ,@      6@      .@      >@      (@      ,@      *@      @      "@      >@      .@      &@      6@     �A@      L@      @      &@      (@      2@      (@      "@      �?       @               @              �?      @      @      @      @      @      @      6@              @       @      @      @              �?      @                                      @      @      @      @      @      @      2@              @      @      @              "@              @               @              �?      �?       @      @      �?      @       @      @                      @              @      *@      ,@      6@      (@      (@      *@      @       @      8@      "@      @      .@      >@      A@      @       @      @      ,@      "@      @      @      @      @      @      @               @       @      �?              @       @      �?               @      @      �?      @      @      $@      0@       @      @       @      @              0@       @      @      (@      6@     �@@      @      @      �?      *@      @      :@      @      "@      @      @              @      $@      :@      �?              &@      6@      :@      @       @              @       @      5@      @       @      @       @              @       @      *@      �?              "@      0@      1@       @       @              @      �?      3@      @       @      @       @              @       @      *@                       @      ,@      0@               @              �?      �?       @                                                                      �?              @       @      �?       @                       @              @              �?       @      @              @       @      *@                       @      @      "@       @                      @      �?       @                       @                      �?      �?      @                              @      @                              �?      �?      @              �?              @               @      �?      @                       @      �?      @       @                      @        �t�bubhhubehhub.