���      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�Ch                                                                	       
                     �t�b�
n_classes_�h�scalar���h"�i8�����R�(Kh&NNNJ����J����K t�bC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h/�C       �t�bK��R�}�(h	K�
node_count�K�nodes�hhK ��h��R�(KK��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hLh/K ��hMh/K��hNh/K��hOh"�f8�����R�(Kh&NNNJ����J����K t�bK��hPhZK ��hQh/K(��hRhZK0��uK8KKt�b�B�                              @�{:<k@I           ��@       	                    @�2S�@           �@                           @������@z           �@                           �?���k~w@�           �@������������������������       ���B�@�           `|@������������������������       ��~:�@�            �g@                          �0@f��MG@�           ��@������������������������       ��VOF�@             7@������������������������       �\x���-@�           �@
                           @�g�漹@�           4�@                           @Q4��(@�           ��@������������������������       �sE��MK@�           �@������������������������       �@x皐@�            �n@                          �7@�P��^@�           �{@������������������������       �4��=��@9           �s@������������������������       ��I�@�            ``@                          �6@Ԁ�\@B           �@                           @�����@�           H�@                          �5@D���c�@�            @������������������������       �x�Ŏ
w@�           pz@������������������������       ��c�ю�@I            @R@                           @����y	@�             c@������������������������       �w�(��@7            �K@������������������������       ������	@b            �X@                          �8@�Ҏ�h@�           �{@                           �?,b���^@�             d@������������������������       �n����Z@             8@������������������������       ���2�>�@�             a@                           �?=��[�@           �q@������������������������       �(�°@@             P@������������������������       �M��2�6@�             k@�t�b�values�hhK ��h��R�(KKKK��hZ�B�        ?@     �V@     ��@     @]@     (�@     ��@     �J@     �r@      2@      @@      @@     �x@      �@      6@     �K@     �z@     �S@     px@     �|@      C@     �i@      *@      3@      .@      q@     ȉ@      (@      :@      l@      @@     �e@     �k@      &@     �X@       @      $@      @     �]@     @}@      @      *@     �W@      (@     �U@      V@      @      C@      �?      @             �P@     �l@       @      "@     �Q@      "@     @P@      O@       @      ;@              �?             �B@     @e@       @      @      8@      @      6@      :@      @      &@      �?      @              >@     �M@       @      *@     @`@      4@      V@     �`@      @     �N@      �?      @      @     �I@     �m@      @              @              @                      @                              �?       @      @      *@     �_@      4@     @U@     �`@      @      L@      �?      @      @      I@     �l@      $@      =@     �i@      G@      k@     �m@      ;@     @Z@      &@      "@      &@     �c@     Pv@      @      9@     @a@      A@     �b@     @e@      5@      O@      &@       @      "@     @]@     `l@      @      8@     �W@      9@      \@      `@      3@      H@      @      @      "@      V@     @e@      @      �?      F@      "@     �B@     �D@       @      ,@      @      �?              =@     �L@      @      @      Q@      (@     �P@      Q@      @     �E@              �?       @     �C@     @`@      @      @      H@      &@     �F@      G@      @      <@              �?             �@@     �U@                      4@      �?      6@      6@              .@                       @      @     �E@      "@     �A@      a@     �C@     �g@     �b@      .@     �X@      @      *@      1@     @^@     pp@      @      8@     @R@      2@     �]@     �T@      $@     �R@      @      $@      ,@     �T@     �`@      @      3@     �L@      .@      U@     �P@      @      K@       @      "@       @      P@     �[@      @      0@     �G@      (@     �R@      O@       @      D@       @       @       @      N@      V@              @      $@      @      "@      @      @      ,@              �?              @      6@      @      @      0@      @     �A@      0@      @      5@       @      �?      @      2@      6@      @              @              1@      @      �?      $@                      �?      "@      @              @      $@      @      2@      *@      @      &@       @      �?      @      "@      1@      @      &@     �O@      5@     �Q@     �P@      @      8@      �?      @      @     �C@     ``@              @      8@      "@      >@      1@      @       @               @      �?      @     �J@                      @      @      @      @       @      �?                                      @              @      5@      @      :@      (@       @      @               @      �?      @      H@      @      @     �C@      (@     �D@     �H@      �?      0@      �?      �?       @      @@     �S@       @      �?      @       @      &@      @      �?      @      �?              �?      (@      1@      �?      @      @@      $@      >@     �E@              *@              �?      �?      4@     �N@�t�bub�_sklearn_version��1.1.3�ub.