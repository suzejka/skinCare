���0      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�CX                                                                	       
       �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K�
node_count�KO�nodes�hhK ��h��R�(KKO��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�BH         F                    @�Eѽb�?s            �\@       3                    @ j�^
�?c            �X@       ,                    @�%69��?E            @Q@                           @9��8���?0             H@       
                     �?�HP��?             9@       	                    �?      �?              @                           6@r�q��?             @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �      �?              @                             @U��6���?             1@                           �?������?             @������������������������       �                     @                           �?      �?             @������������������������       �      �?              @������������������������       �                      @                           �?{�G�z�?
             $@                          �1@      �?              @������������������������       �                     �?                           3@������?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                          �4@���Q��?             @������������������������       �                     �?                           �?      �?             @������������������������       �      �?              @������������������������       �      �?              @������������������������       �                      @       '                      @x�W��#�?             7@       &                    �?������?             .@        %                     �?X�<ݚ�?	             "@!       $                    @���Q��?             @"       #                    3@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �      �?              @������������������������       �      �?             @������������������������       �                     @(       )                   �2@      �?              @������������������������       �                      @*       +                    �?�8��8��?             @������������������������       �      �?              @������������������������       �      �?             @-       0                    �?؇���X�?             5@.       /                   �2@�<ݚ�?	             "@������������������������       �                     @������������������������       ��q�q�?             @1       2                     �?�8��8��?             (@������������������������       �r�q��?             @������������������������       �                     @4       ;                    @k�Y�H��?             >@5       6                   �2@�m۶m��?             ,@������������������������       �                     &@7       :                    �?�q�q�?             @8       9                   �5@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?<       ?                     �?     @�?             0@=       >                    @r�q��?             @������������������������       �z�G�z�?             @������������������������       �                     �?@       C                    4@���Q��?
             $@A       B                    �?r�q��?             @������������������������       �                      @������������������������       �      �?             @D       E                    �?      �?             @������������������������       �      �?              @������������������������       �                      @G       H                    �?     ��?             0@������������������������       �                     @I       N                    @�z�G��?
             $@J       K                   �2@�q�q�?	             "@������������������������       �                     �?L       M                     �?      �?              @������������������������       �      �?              @������������������������       ��q�q�?             @������������������������       �                     �?�t�b�values�hhK ��h��R�(KKOKK��hV�B(        *@      �?      ,@      @      9@      *@      5@      @       @      0@      �?      *@      �?      ,@      @      6@      *@      5@      @       @      @      �?       @              ,@      @      .@       @      5@               @      @      �?       @              ,@      @      (@       @      @               @      @      �?                      @              @       @      �?               @      @      �?                                      �?      @      �?              �?                                                      �?      @                                                                                      @                                                                              �?       @                                                                                              �?              �?                                      @              @      @                      �?      @      �?                      @              �?                                      @                                                                                      @                              @              �?                                                                      �?              �?                                                                       @                                                                                                      @      @                      �?              �?                                      @      @                      �?              �?                                                                      �?                                                      @      @                                      �?                                              �?                                      �?                                              �?                                                                                                                              �?                                      @       @                                                                              �?                                                                                       @       @                                                                              �?      �?                                                                              �?      �?                                                                               @                                                       @              &@      @      @               @                                                      &@              @                                                                      @              @                                                                       @              @                                                                      �?               @                                                                                      �?                                                                      �?              �?                                                                      �?              �?                                                                      @              �?                                                                      @                                                                       @                      @      �?               @                                                                                       @                                       @                      @      �?                                                      �?                              �?                                                      �?                      @                                                                                              @              2@                                                                       @              @                                                                                      @                                                                       @              @                                                                      �?              &@                                                                      �?              @                                                                                      @                                      &@      �?                      @      @              @                              &@      �?                       @                                                      &@                                                                                              �?                       @                                                              �?                      �?                                                              �?                                                                                                              �?                                                                                      �?                                                                                      @      @              @                                                              �?      @                                                                              �?      @                                                                                      �?                                                                              @                      @                                                              �?                      @                                                                                       @                                                              �?                      @                                                              @                      �?                                                              �?                      �?                                                               @                                                                                      @                                      *@                                                                                      @                                              @                                      @                                              @                                      @                                                                                      �?                                              @                                      @                                              �?                                      �?                                               @                                      @                                                                                      �?        �t�bub�_sklearn_version��1.1.0�ub.