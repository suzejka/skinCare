���H      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K.�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C`                                                                	       
              �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K	�
node_count�Ks�nodes�hhK ��h��R�(KKs��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B(         *                    �?fY�eY��?�             e@                          �5@R=6�z�?A            @P@       
                    �?Z�K8�?             :@                           �?:/����?             @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?       	                   �4@      �?             @������������������������       �                      @������������������������       �      �?              @                           @|�ʒ���?             3@                           @�X�C�?             ,@                          �4@�$I�$I�?             @������������������������       ����Q��?             @������������������������       �      �?              @                           �?և���X�?             @                           3@�q�q�?             @������������������������       �                     �?������������������������       �                      @                            �?      �?             @������������������������       �                      @������������������������       �      �?              @������������������������       �                     @       %                     @>L�*:�?'            �C@                           @��kv�?             5@������������������������       �        	             "@                           �?�������?             (@                           9@      �?             @������������������������       �                     @������������������������       �                     �?       $                    A@      �?              @        !                   �7@؇���X�?             @������������������������       �                     @"       #                    <@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?&       '                    <@0�����?             2@������������������������       �                     0@(       )                   @@@      �?              @������������������������       �                     �?������������������������       �                     �?+       d                    @���r�?g            �Y@,       O                    @(��(���?T             U@-       @                    @�2�,E�?5            �J@.       7                    @{��?��?             ?@/       2                    5@޾�z�<�?             *@0       1                     �?؇���X�?             @������������������������       ��q�q�?             @������������������������       �                     @3       4                     �?�q�q�?             @������������������������       �                     @5       6                      @�q�q�?             @������������������������       �                     �?������������������������       �      �?              @8       =                    @VUUUUU�?             2@9       <                    �?�eP*L��?             &@:       ;                   �2@���Q��?
             $@������������������������       �      �?             @������������������������       ��q�q�?             @������������������������       �                     �?>       ?                   �2@������?             @������������������������       �      �?             @������������������������       ��q�q�?             @A       L                   �5@"pc�
�?             6@B       K                    @R���Q�?             4@C       J                   �2@     ��?             0@D       G                     @d}h���?             ,@E       F                    �?"pc�
�?             &@������������������������       �؇���X�?             @������������������������       �      �?             @H       I                    �?�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                      @������������������������       �                     @M       N                    @      �?              @������������������������       �                     �?������������������������       �                     �?P       [                    �?�5�`���?             ?@Q       Z                    !@/y0��k�?             *@R       S                    @���!pc�?             &@������������������������       �                     @T       Y                    @      �?             @U       V                   �3@���Q��?             @������������������������       �                     �?W       X                    @      �?             @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @\       a                   �;@��Hx��?             2@]       `                   �2@�Q����?             .@^       _                     �?��Q��?
             $@������������������������       ��q�q�?             @������������������������       �      �?             @������������������������       �                     @b       c                   �?@�q�q�?             @������������������������       �                      @������������������������       �                     �?e       n                   �8@�p9W���?             3@f       i                   �2@.y0��k�?             *@g       h                    �?      �?              @������������������������       �                     �?������������������������       �                     �?j       m                   �4@�C��2(�?             &@k       l                    �?r�q��?             @������������������������       �                      @������������������������       �      �?             @������������������������       �                     @o       p                    @�8��8��?             @������������������������       �                     @q       r                   �;@�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�b�values�hhK ��h��R�(KKsKK��hV�B +        �?      .@      9@      �?      @      4@       @      I@      $@      <@      &@       @      �?      @              �?      @      0@               @      @      0@      $@       @              @              �?                               @              .@               @              @                                                               @               @                                                                              �?               @                                                                                               @                                                                              �?                              @                                                              �?                               @                                                                                              �?                                                              �?                              @              �?                               @              *@                              @              �?                               @               @                                              �?                               @              @                                                                               @              @                                              �?                                              �?                              @                                                              @                               @                                                              �?                                                                                              �?                               @                                                                                              �?                                                              @                                                                                               @                              �?                                                              �?                                                                                              @                      �?      �?                      @      0@                      @      �?      $@                      �?                      @                              @              $@                                                                                              "@                      �?                      @                              @              �?                                              @                              �?                                                              @                                                                                                                              �?                                      �?                                                      @              �?                      �?                                                      @                                                                                              @                                      �?                                                       @                                      �?                                                                                                                                                       @                                                                                                              �?              �?                                      0@                              �?                                                              0@                                                      �?                                                                      �?                      �?                                                                                                                                                                      �?                               @      9@                      @       @      H@      @      (@      �?                       @      ,@                       @       @      G@              &@      �?                       @      @                                      A@               @                               @      @                                      0@              @                                      �?                                      $@               @                                      �?                                      @                                                      �?                                       @                                                                                              @                                                                                              @               @                                                                              @                                                                                              �?               @                                                                                              �?                                                                              �?              �?                               @       @                                      @               @                              @                                              @                                              @                                              @                                               @                                               @                                              @                                               @                                                                                              �?                                               @       @                                      �?               @                              �?       @                                      �?                                              �?                                                               @                                                                              2@              @                                                                              1@              @                                                                              *@              @                                                                              &@              @                                                                              "@               @                                                                              @              �?                                                                              @              �?                                                                               @              �?                                                                              �?              �?                                                                              �?                                                                                               @                                                                                              @                                                                                              �?              �?                                                                                              �?                                                                              �?                                                      &@                       @       @      (@              @      �?                               @                               @      @                                                       @                                      @                                                      @                                                                                              @                                      @                                                      @                                       @                                                      �?                                                                                               @                                       @                                                       @                                      �?                                                                                              �?                                                                                              �?                                                                                       @                                                              @                       @              "@              @      �?                              @                                      "@              @                                      @                                      @              @                                       @                                      @                                                      �?                                                      @                                                                              @                                                                               @                                      �?                                                       @                                                                                                                                      �?                              &@                       @               @      @      �?                                      &@                                      �?              �?                                      �?                                                      �?                                      �?                                                                                                                                                      �?                                      $@                                      �?                                                      @                                      �?                                                       @                                                                                              @                                      �?                                                      @                                                                                                                       @              �?      @                                                                                              @                                                                       @              �?                                                                                              �?                                                                               @                                                �t�bub�_sklearn_version��1.1.0�ub.