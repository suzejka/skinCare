���O      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�Ch                                                                	       
                     �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K�
node_count�Ky�nodes�hhK ��h��R�(KKy��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�Bx         f                   �9@6�����?�             e@       E                   �5@�[N����?�            �a@       4                     @���4��?c            �X@       1                    @�%�e��?I            @R@                           �?�����k�?E            @Q@                           �?������?             .@                           3@      �?             @������������������������       �                     �?	       
                    �?�q�q�?             @������������������������       �      �?              @������������������������       �                     �?                           �?"pc�
�?             &@������������������������       ��q�q�?             @������������������������       �                     @       "                    @�-����?6             K@                          �1@�ʻ����?"             A@                           @�eP*L��?             &@                           �?X�<ݚ�?	             "@������������������������       ����Q��?             @������������������������       �      �?             @������������������������       �                      @                           �?D%��N��?             7@                            �?�<ݚ�?             2@������������������������       �      �?              @                            �?     ��?             0@������������������������       �                     @                           �?���!pc�?             &@������������������������       �                     �?                           @z�G�z�?
             $@������������������������       ����Q��?             @������������������������       �                     @        !                   �3@{�G�z�?             @������������������������       �                     �?������������������������       �      �?             @#       $                    @���(\��?             4@������������������������       �                      @%       *                    @X�<ݚ�?             2@&       )                    2@      �?              @'       (                    �?�q�q�?             @������������������������       �      �?              @������������������������       �      �?             @������������������������       �                      @+       .                    �?���Q��?
             $@,       -                     �?      �?             @������������������������       �      �?              @������������������������       �      �?              @/       0                    @�q�q�?             @������������������������       ��q�q�?             @������������������������       ��q�q�?             @2       3                    !@      �?             @������������������������       �                      @������������������������       �      �?              @5       >                    @
j*D>�?             :@6       =                    �?�q�q�?             2@7       8                    �?և���X�?             ,@������������������������       �                     @9       :                    @���!pc�?             &@������������������������       �                     �?;       <                    �?�z�G��?
             $@������������������������       �      �?             @������������������������       ��q�q�?             @������������������������       �                     @?       D                   �3@      �?              @@       C                   �2@���Q��?             @A       B                    @      �?             @������������������������       �      �?              @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     @F       ]                     @X�EQ]N�?+            �E@G       X                    @ �o_��?             9@H       M                   �7@ԍx�V�?             3@I       J                    �?:/����?             @������������������������       �                      @K       L                   �6@���Q��?             @������������������������       �                     @������������������������       �                      @N       W                   �8@�q�q�?             (@O       V                    @���!pc�?             &@P       U                    @և���X�?             @Q       T                    @�q�q�?             @R       S                    �?���Q��?             @������������������������       �      �?             @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?Y       Z                     �?VUUUUU�?             @������������������������       �                      @[       \                    @      �?             @������������������������       �                      @������������������������       �                      @^       a                    �?�Kh/��?             2@_       `                    @VUUUUU�?             @������������������������       �      �?              @������������������������       �                     �?b       c                    �?���Q��?             .@������������������������       ��q�q�?             @d       e                     @�8��8��?             (@������������������������       �r�q��?             @������������������������       �                     @g       l                     �?��k����?             :@h       k                    @      �?              @i       j                   �@@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @m       x                     @����H�?             2@n       w                    @�"�O�|�?             1@o       r                    �?      �?              @p       q                    �?�q�q�?             @������������������������       �                     �?������������������������       �      �?              @s       v                    �?���Q��?             @t       u                    �?      �?             @������������������������       �      �?              @������������������������       �      �?              @������������������������       �                     �?������������������������       �        	             "@������������������������       �                     �?�t�b�values�hhK ��h��R�(KKyKK��hV�B(1        2@      Q@      4@       @      @       @      ;@      *@       @       @       @      @      @      2@      Q@      @       @      @       @      7@      *@       @      �?               @      �?      .@     �M@       @      �?      @              0@                      �?                      �?      @      F@       @      �?      @              0@                      �?                      �?      @      F@       @              @              ,@                                              �?      @      &@                                                                                               @       @                                                                                                      �?                                                                                               @      �?                                                                                              �?      �?                                                                                              �?                                                                                                       @      "@                                                                                               @      @                                                                                                      @                                                                                                     �@@       @              @              ,@                                              �?              5@                                      (@                                              �?              @                                      @                                                              @                                      @                                                              @                                       @                                                               @                                       @                                                                                                       @                                                              0@                                      @                                              �?              ,@                                      @                                                              �?                                      �?                                                              *@                                      @                                                              @                                                                                                       @                                      @                                                                                                      �?                                                               @                                       @                                                              @                                       @                                                              @                                                                                                       @                                       @                                              �?                                                                                                      �?               @                                       @                                                              (@       @              @               @                                                                       @                                                                                              (@                      @               @                                                              @                                       @                                                              @                                       @                                                              �?                                      �?                                                              @                                      �?                                                               @                                                                                                      @                      @                                                                               @                       @                                                                              �?                      �?                                                                              �?                      �?                                                                              @                       @                                                                               @                      �?                                                                               @                      �?                                                                                              �?                       @                      �?                                                                               @                                                                              �?                                              �?                              &@      .@                                                                                              @      (@                                                                                              @       @                                                                                              @                                                                                                      @       @                                                                                                      �?                                                                                              @      @                                                                                              �?      @                                                                                               @      @                                                                                                      @                                                                                              @      @                                                                                               @      @                                                                                               @       @                                                                                              �?      �?                                                                                              �?      �?                                                                                                      �?                                                                                              @                                                                                                      @      "@       @      �?       @       @      @      *@       @                       @               @       @       @               @       @      @               @                      �?                       @                               @      @               @                      �?                                                       @      @               @                                                                                                       @                                                                               @      @                                                                                                      @                                                                                               @                                                                       @                                      @                                      �?                       @                                      @                                                              @                                      @                                                              @                                       @                                                              @                                       @                                                              @                                      �?                                                                                                      �?                                                              �?                                                                                                                                              �?                                                              @                                                                                                                                                                                      �?               @               @               @                                                                       @                                                                                                                       @               @                                                                                       @                                                                                                                       @                                                                      �?      �?              �?                      �?      *@                              �?              �?      �?                                      �?                                                              �?                                      �?                                                      �?                                                                                                                              �?                              *@                              �?                                      �?                               @                                                                                                      &@                              �?                                                                      @                              �?                                                                      @                                                              0@                              @                      �?       @      �?       @                       @                              @                               @                                       @                              @                                                                                                      @                                                                       @                                                                                                                                                                       @                                      ,@                                                      �?              �?       @                      ,@                                                      �?                       @                      @                                                      �?                       @                       @                                                      �?                                              �?                                                                                                      �?                                                      �?                                              @                                                                               @                       @                                                                               @                      �?                                                                              �?                      �?                                                                              �?                      �?                                                                                                      "@                                                                                                                                                                              �?        �t�bub�_sklearn_version��1.1.0�ub.