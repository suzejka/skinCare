����      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K
�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C�                                                                	       
                                                                                           �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K
�
node_count�K��nodes�hhK ��h��R�(KK���h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�Bh         R                   �5@�^<��@�             c@       ;                    @ �X��@g            �Y@       $                     @�?aO @N            �S@                           �?e���@0             H@                            �?7�nt�?             ,@                           �?�+��&�?             (@������������������������       �                     @       	                    �?�t�I�|�?	             "@������������������������       �_�z|�X�?             @
                           3@|%��b�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                      @       !                   �4@I`1*ĸ @"             A@                           �?X��ܳ�?             ?@                           @Ո����?             0@                           @      �?              @                            �?      �?             @������������������������       �|%��b�?             @������������������������       �                     �?                            �?�c�����?             @������������������������       �                     �?������������������������       �|%��b�?             @                           �?c�YB�d�?              @������������������������       ��c�����?             @������������������������       �                     @                            �?�n$����?             .@                            �?���'���?             @������������������������       �|%��b�?             @������������������������       �                     �?                            �?c�YB�d�?              @������������������������       ��c�����?             @������������������������       �                     @"       #                    !@|%��b�?             @������������������������       �                     �?������������������������       �                      @%       *                    �?y�*p{��?             >@&       '                   �2@���� ��?             @������������������������       �                     @(       )                    4@h���\�?             @������������������������       �                     �?������������������������       �      �?              @+       0                    �?!}=�K�?             8@,       -                    �?���xp��?             .@������������������������       �                      @.       /                   �1@�9>����?             @������������������������       �                      @������������������������       ��Z���?             @1       :                   �4@t�&-�?	             "@2       3                    @��b}�?              @������������������������       �      �?              @4       5                    @      �?             @������������������������       �                     �?6       7                    @��&��?             @������������������������       �                      @8       9                    �?|%��b�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?<       ?                   �0@&MI`@             9@=       >                    �?�Z���?             @������������������������       �                     �?������������������������       ��c�����?             @@       K                   �4@Se���?             4@A       B                     �?/��PL��?             (@������������������������       �                     �?C       D                   �1@Ҙ�W���?             &@������������������������       �                     �?E       J                    @
����3�?
             $@F       I                    �?|%��b�?	             "@G       H                     �?�c�����?             @������������������������       �|%��b�?             @������������������������       �                     �?������������������������       ���&��?             @������������������������       �                     �?L       M                    @��'4���?              @������������������������       �                     �?N       O                    �?������?             @������������������������       �                     �?P       Q                    @|%��b�?             @������������������������       �      �?              @������������������������       ��c�����?             @S       j                    �?�)'@2             I@T       c                   �8@dHRb�	@             7@U       ^                     �?|R��>@             0@V       Y                    �?      @              @W       X                    @      �?             @������������������������       �      �?              @������������������������       �      �?              @Z       [                   �6@      �?             @������������������������       �                      @\       ]                   �7@      �?              @������������������������       �                     �?������������������������       �                     �?_       b                    7@�1H����?              @`       a                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @d       g                    >@.��Zz�?             @e       f                   �:@|%��b�?             @������������������������       �                     �?������������������������       �                      @h       i                   �@@�c�����?             @������������������������       �                     �?������������������������       �                     @k       x                    �?f�>��@             ;@l       q                   �6@���@             (@m       p                     @h���\�?             @n       o                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?r       w                    @oS�<��?	             "@s       v                    @��'4���?              @t       u                     @�Z���?             @������������������������       �                     @������������������������       �      �?              @������������������������       �h���\�?             @������������������������       �                     �?y       �                     �?��9�s@             .@z       }                    7@�,�4�?             @{       |                     �?|%��b�?             @������������������������       �                      @������������������������       �                     �?~                           :@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �9@|R��>@              @�       �                    @>���i��?             @������������������������       �                     �?�       �                    @�c�����?             @������������������������       �                      @�       �                   �8@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �;@|%��b�?             @������������������������       �                     �?������������������������       �                      @�t�b�values�hhK ��h��R�(KK�KK��hV�B�c        "@      9@      1@      @      "@       @      @      @      1@       @      9@      @      �?       @       @       @       @       @      @      @      �?       @       @       @      6@      1@               @              @              $@              8@                              �?       @                              @      �?              �?       @      0@      1@               @                              @              8@                              �?       @                              @      �?                       @      $@      1@              @                               @              @                              �?       @                                                               @      @       @                                                              @                                                                                                              @       @                                                              @                                                                                                                                                                                      @                                                                                                              @       @                                                              @                                                                                                              �?       @                                                              @                                                                                                               @                                                                      �?                                                                                                              �?                                                                                                                                                                                      �?                                                                      �?                                                                                                       @                                                                                                                                                                                              @      .@              @                               @                                              �?       @                                                                      @      .@              @                               @                                                                                                                              @      @              @                               @                                                                                                                               @      @                                               @                                                                                                                              �?      �?                                               @                                                                                                                              �?                                                       @                                                                                                                                      �?                                                                                                                                                                              �?      @                                                                                                                                                                                      �?                                                                                                                                                                              �?       @                                                                                                                                                                              �?                      @                                                                                                                                                              �?                      @                                                                                                                                                                                      @                                                                                                                                                              @      &@                                                                                                                                                                              @      @                                                                                                                                                                               @      @                                                                                                                                                                              �?                                                                                                                                                                                      �?      @                                                                                                                                                                              �?      @                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                      �?       @                                                                                                                                                                              �?                                                                                                                                                                                               @                                                                      @                      �?                              �?              1@                                                                      @      �?                              �?                                                      �?                                                                                      @      �?                                                                                                                                                                              @                                      �?                                                      �?                                                                                              �?                                                                                                                                                                                      �?                              �?                                                      �?                                                                                                                              @                      �?                                              1@                                                                      �?                                      �?                                                                      ,@                                                                                                                                                                                       @                                                                                                              �?                                                                      @                                                                                                                                                                                       @                                                                                                              �?                                                                      @                                                                                                              @                      �?                                              @                                                                      �?                                      @                      �?                                              @                                                                                                              �?                      �?                                                                                                                                                              @                                                                      @                                                                                                                                                                                      �?                                                                                                              @                                                                       @                                                                                                               @                                                                                                                                                                                      �?                                                                       @                                                                                                                                                                                       @                                                                                                              �?                                                                                                                                                                                                                                                                                                                                      �?                              @      @                                      @              @                                                                                      �?                      �?              �?                                      @                                                                                                                                                                                      �?                                                                                                                                              �?                                      @                                                                                                                                      @      @                                                      @                                                                                      �?                      �?      �?      @                                                      @                                                                                                              �?                                                                                                                                                                                      �?      �?      @                                                      @                                                                                                                      �?                                                                                                                                                                                              @                                                      @                                                                                                                              @                                                      @                                                                                                                              �?                                                      @                                                                                                                              �?                                                       @                                                                                                                                                                                      �?                                                                                                                               @                                                      @                                                                                                                                                                                      �?                                                                                                                      @       @                                                                                                                                              �?                                                                                                                                                                                      �?                              @       @                                                                                                                                                                              �?                                                                                                                                                                                      @       @                                                                                                                                                                              �?      �?                                                                                                                                                                              @      �?                                                                                                                                                                              �?      @              @      �?       @       @      @      @       @      �?      @      �?       @      �?               @       @      @       @               @      �?              �?              �?               @               @      �?       @              @      �?                               @              @       @                                      �?                               @               @      �?                                                               @              @       @                                                                       @               @      �?                                                               @                      �?                                                                       @                                                                                       @                                                                                              �?                                                                                      �?                                                                                              �?                                                                                      �?                                                                                                               @      �?                                                                                      �?                                                                                       @                                                                                                                                                                                              �?                                                                                      �?                                                                                              �?                                                                                                                                                                                                                                                                              �?                                      �?                                                                                                                                      @      �?                                      �?                                                                                                                                              �?                                                                                                                                                                                      �?                                      �?                                                                                                                                                                                                                                                                                                                              @                                                              �?                                               @              @      �?                                                                                                              �?                                               @                                                                                                                                      �?                                                                                                                                                                                                                                       @                                                                                                                                                                                                      @      �?                                                                                                                                                                                      �?                                                                                                                                                                              @                                                                                              �?       @              @      �?               @      @      @              �?                       @      �?                       @                               @      �?               @                                      �?      �?      @              �?                                                                                              �?                                                              �?      �?              �?                                                                                                                                                              �?      �?                                                                                                                                                                                      �?                                                                                                                                                                              �?                                                                                                                                                                                                              �?                                                                                                               @                                      �?              @                                                                                                              �?               @                                      �?              @                                                                                                                              �?                                                      @                                                                                                                                                                                      @                                                                                                                              �?                                                      �?                                                                                                                              �?                                      �?              �?                                                                                                                                                                                                                                                                                                      �?      �?                      @      �?              �?       @                                               @      �?                       @                               @                                                                                                                       @      �?                       @                               @                                                                                                                              �?                                                       @                                                                                                                                                                                       @                                                                                                                              �?                                                                                                                                                                               @                               @                                                                                                                                                       @                                                                                                                                                                                                                       @                                              �?                      @      �?              �?       @                                                                                                                              �?                      @      �?                                                                                                                                                      �?                                                                                                                                                                                                              @      �?                                                                                                                                                                               @                                                                                                                                                                                      �?      �?                                                                                                                                                                                      �?                                                                                                                                                                              �?                                                                                                                                                                                                              �?       @                                                                                                                                                                              �?                                                                                                                                                                                               @                                                                                                                        �t�bub�_sklearn_version��1.1.0�ub.