��u      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C(                                    �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K�
node_count�K9�nodes�hhK ��h��R�(KK9��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�Bx                              @�������?s            �\@                            �?�R$�?Q            @T@                           @��w+��?2             I@                           3@b�$�?%            �B@       
                    @���l��?             0@                            �?"S,f�B�?             &@������������������������       �                      @       	                    �?�Q$��?	             "@������������������������       �|%��b�?             @������������������������       �|%��b�?             @������������������������       �                     @                           �?��0\^�?             5@������������������������       �                      @                          �4@vׯD�"�?             3@                            �?���'���?             @������������������������       �                     @������������������������       �                     @������������������������       �                     (@                           @���q"
�?             *@������������������������       �                     (@������������������������       �                     �?                           7@�3>�f�?             ?@������������������������       �                     ;@                           �?      �?             @������������������������       �                      @������������������������       �                      @       0                    @(�����?"             A@       )                    �?i�q]�?             4@       &                   �4@l�ɾ���?
             $@       #                    �?_�z|�X�?             @                           �1@|%��b�?             @������������������������       �                     �?!       "                    �?      �?              @������������������������       �                     �?������������������������       �                     �?$       %                     @|%��b�?             @������������������������       �                     �?������������������������       �      �?              @'       (                    �?�c�����?             @������������������������       �      �?              @������������������������       �                      @*       +                    �?��Yo��?
             $@������������������������       �                     �?,       /                   �2@M�)9��?	             "@-       .                    @�Z���?             @������������������������       �                     @������������������������       �      �?              @������������������������       �                     @1       2                    @�9>����?             ,@������������������������       �        	             "@3       8                    �?��&��?             @4       5                   �3@|%��b�?             @������������������������       �                     �?6       7                   �5@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�t�b�values�hhK ��h��R�(KK9KK��hV�B�        (@      F@     �@@      �?      9@       @      F@      9@              $@       @      .@      7@              $@       @      @      7@              "@                      @              "@                      @              @                       @                                      @              @                      �?               @                      @               @                                      @       @      @      0@                       @                                              @      0@                              @      @                              @                                              @                                      (@                              (@                      �?              (@                                                              �?              =@       @                              ;@                                       @       @                               @                                               @                      $@               @      �?      .@      $@              @      �?      @       @              @              @      �?               @              @                       @              �?                      �?                                      �?              �?                      �?                                                      �?      �?                               @                                      �?      �?                              �?      �?              @                      �?              �?                                       @                       @              �?      �?                              �?                       @                      �?              @                      �?              @                                      �?                      �?              @                                                       @              (@                                      "@                       @              @                       @              �?                      �?                                      �?              �?                                      �?                      �?                                                       @�t�bub�_sklearn_version��1.1.0�ub.