��B^      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K&�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C�                                                                	       
                                          �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K�
node_count�K}�nodes�hhK ��h��R�(KK}��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�BX         N                   �5@�5;j��?�             e@       9                     @䃞ͪ��?d             Y@       0                    @h�m��?J            �R@       	                   �0@     D�?@             P@                           �?z�G�z�?
             $@������������������������       �                      @                           @      �?              @������������������������       �z�G�z�?             @������������������������       ��q�q�?             @
                          �1@���e/�?6             K@                            @r�q��?             (@������������������������       �                     �?                           �?"pc�
�?             &@������������������������       �r�q��?             @������������������������       �z�G�z�?             @       #                    @~VC�1��?*             E@                           �?UUUUUU�?             8@                            �?�T�6|��?             *@                          �4@VUUUUU�?	             "@������������������������       ����Q��?             @                           �?      �?             @������������������������       �      �?              @������������������������       �                      @                           �?      �?             @������������������������       �      �?              @������������������������       �                      @       "                   �4@j�V���?             &@       !                    @z�G�z�?
             $@                            �?����X�?             @                            �?���Q��?             @������������������������       ��q�q�?             @������������������������       �      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     �?$       )                    @2�tk~X�?             2@%       (                    �?      �?             (@&       '                    3@�q�q�?	             "@������������������������       ��q�q�?             @������������������������       ��q�q�?             @������������������������       �                     @*       +                    @�q�q�?             @������������������������       �                      @,       /                   �3@      �?             @-       .                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @1       2                   �0@p=
ףp�?
             $@������������������������       �                     �?3       8                    @�<ݚ�?	             "@4       5                   �2@      �?             @������������������������       �                     �?6       7                     �?�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                     @:       I                    @pƵHPS�?             :@;       >                    �?g\�5�?             *@<       =                   �3@      �?             @������������������������       �                      @������������������������       �      �?              @?       H                    �?�n���?	             "@@       E                    @      �?              @A       D                    �?���Q��?             @B       C                    �?      �?             @������������������������       �      �?              @������������������������       �      �?              @������������������������       �                     �?F       G                    �?VUUUUU�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     �?J       M                    �?$�q-�?             *@K       L                     @�����H�?	             "@������������������������       �؇���X�?             @������������������������       �                      @������������������������       �                     @O       \                    �?}�@�m�?D             Q@P       Y                   �:@s
^N���?             ,@Q       V                    �?�<ݚ�?	             "@R       S                     �?�$I�$I�?             @������������������������       �      �?             @T       U                    @�q�q�?             @������������������������       �      �?              @������������������������       �                     �?W       X                    @      �?              @������������������������       �                     �?������������������������       �                     �?Z       [                    �?���Q��?             @������������������������       �                     @������������������������       �                      @]       f                   �6@�}���?6             K@^       a                    �?      �?              @_       `                    @      �?             @������������������������       �                     �?������������������������       �                     @b       e                    @      �?             @c       d                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @g       r                    @��	,UP�?.             G@h       m                   �<@�q-��?             *@i       j                    �?      �?              @������������������������       �                     @k       l                    :@      �?              @������������������������       �                     �?������������������������       �                     �?n       q                    �?
ףp=
�?             @o       p                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       ��q�q�?             @s       t                    �?ҿЈ:G�?!            �@@������������������������       �                     3@u       |                   �9@>4և���?             ,@v       w                    �?      �?              @������������������������       �                     @x       y                    @�Q����?             @������������������������       �                      @z       {                     �?VUUUUU�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                     @�t�b�values�hhK ��h��R�(KK}KK��hV�B�>        *@       @       @       @      @      9@       @      G@      �?      �?      @       @      =@      7@      �?      &@      "@                               @      5@       @      @                                      <@      6@              $@       @                               @      ,@       @      @                                      (@      6@              $@       @                               @      (@       @      @                                      (@      6@              @                                               @                                                               @                                                                                                                               @                                                               @                                                              @                                                              �?                                                              @                                                              �?                                                               @                       @                               @      $@       @      @                                      (@      ,@              @                                               @                                                      "@      �?                                                                                                                              �?                                                               @                                                      "@                                                                      �?                                                      @                                                                      �?                                                      @                               @                               @       @       @      @                                      @      *@              @       @                                      @               @                                      @      @              @                                              @              �?                                      @      @              @                                              @                                                      @      @                                                               @                                                      @                                                                      �?                                                              @                                                              �?                                                              �?                                                                                                                               @                                                                              �?                                                              @                                                              �?                                                              �?                                                                                                                               @       @                                       @              �?                                                                       @                                       @                                                                                      @                                       @                                                                                      @                                       @                                                                                       @                                      �?                                                                                      �?                                      �?                                                                                       @                                                                                                                              @                                                                                                                                                                                      �?                                                                                                       @      @       @      �?                                              $@                                                              @                                                              "@                                                              @                                                              @                                                              �?                                                               @                                                               @                                                              @                                                                                                                              @                                                       @               @      �?                                              �?                                                                       @                                                                                                               @                      �?                                              �?                                                                              �?                                              �?                                                                              �?                                                                                                                                                                              �?                                                       @                                                                                                                                       @              �?                                                              @                                                              �?                                                                                                               @                                                                              @                                               @                                                                               @                                                                                                                              �?                                               @                                                                              �?                                              �?                                                                                                                              �?                                                                              �?                                                                                                                              @      �?                                      @               @                                      0@                              �?                                      @               @                                      @                              �?                                      @                                                                                                                               @                                                                                      �?                                      �?                                                                                                                              @               @                                      @                                                                      @              �?                                      @                                                                       @                                                      @                                                                       @                                                       @                                                                      �?                                                      �?                                                                      �?                                                      �?                                                                                                                              �?                                                                      �?              �?                                      �?                                                                      �?                                                      �?                                                                                      �?                                                                                                                              �?                                                                                                              �?                                                      (@                                                                      �?                                                       @                                                                      �?                                                      @                                                                                                                               @                                                                                                                              @                              @       @       @       @      @      @              D@      �?      �?      @       @      �?      �?      �?      �?      @                                       @               @                      @       @                              �?      @                                       @               @                                                              �?      @                                      �?               @                                                                      @                                      �?                                                                                      �?                                                       @                                                                      �?                                                      �?                                                                                                                              �?                                                                                                              �?                                                                              �?                                              �?                                                                                                                                                                                                              �?                                                                                      @       @                                                                                                                      @                                                                                                                                       @                                               @       @       @      @       @              C@      �?      �?                      �?      �?      �?                                       @              �?              @                                      �?              �?                                                                      @                                      �?                                                                                                                              �?                                                                                      @                                                                                               @              �?                                                                      �?                                                      �?                                                                      �?                                                      �?                                                                                                                                                                                                      �?                                       @                                                                                                               @       @              @      �?             �A@      �?      �?                              �?                               @       @                                      @      �?      �?                                                              �?                                              @                                                                                                                              @                                                                              �?                                              �?                                                                              �?                                                                                                                                                                              �?                                                                              �?       @                                              �?      �?                                                                                                                      �?      �?                                                                                                                      �?                                                                                                                                      �?                                                              �?       @                                                                                                                                              @      �?              <@                                              �?                                                                              3@                                                                                                      @      �?              "@                                              �?                                                      @      �?              @                                              �?                                                                              @                                                                                                      @      �?                                                              �?                                                       @                                                                                                                              �?      �?                                                              �?                                                      �?                                                                                                                                      �?                                                              �?                                                                              @                                                                �t�bub�_sklearn_version��1.1.0�ub.