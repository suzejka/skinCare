���y      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C�                                                                	       
                                                                                           �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K
�
node_count�K}�nodes�hhK ��h��R�(KK}��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�BX         8                   �4@��f��@�             e@       )                    @��H�	@Y            @V@                            @Ok��@F            �Q@                           �?�5�� @-            �F@                          �2@>���i��?
             $@������������������������       �                     @������������������������       �n���?             @                           �?�p����?#            �A@	                           @H:�$s>�?             2@
                           @���G�?             @                            �?|%��b�?             @������������������������       �                      @������������������������       �                     �?                           2@�c�����?             @������������������������       �                      @������������������������       �      �?              @                           �?��Ȓ���?             &@������������������������       �V�T����?             @������������������������       ��Z���?             @                            �?~��kp��?             1@                           2@������?             @������������������������       ��Z���?             @������������������������       �      �?              @                           �?���?
             $@������������������������       �V�T����?             @������������������������       �                     @       &                    @H�X���?             9@                           �?t�r�v��?             &@������������������������       �                      @       %                    �?h���\�?	             "@       "                    �?J��MY.�?             @        !                     @|%��b�?             @������������������������       �      �?              @������������������������       �                     �?#       $                   �2@      �?             @������������������������       �                     �?������������������������       �h���\�?             @������������������������       �                      @'       (                    �?���;E��?             ,@������������������������       �                      @������������������������       �V�T����?             @*       /                    �?+5��/��?             3@+       .                    �?�c�����?             (@,       -                    @�9>����?             @������������������������       ��c�����?             @������������������������       �                     @������������������������       ���&��?             @0       3                    @��Z-�@             @1       2                     �?|%��b�?             @������������������������       �                     �?������������������������       �                      @4       5                     �?      �?             @������������������������       �                     �?6       7                    �?|%��b�?             @������������������������       �                     �?������������������������       �      �?              @9       n                   �8@�5m��@O            �S@:       [                   �6@���ES@:             M@;       D                     �?�����	@             <@<       ?                    �?�K�܏?@	             "@=       >                    @|%��b�?             @������������������������       �      �?              @������������������������       �                     �?@       A                   �5@h���\�?             @������������������������       �                      @B       C                    @      �?             @������������������������       �                      @������������������������       �                      @E       P                     �?mJ�X��@             3@F       O                    @3chd���?             (@G       N                   �5@�ڰ`+��?
             $@H       I                    �?�!]]t�?	             "@������������������������       �                     @J       K                    @|%��b�?             @������������������������       �                     �?L       M                    @��&��?             @������������������������       �      �?              @������������������������       �|%��b�?             @������������������������       �                     �?������������������������       �                      @Q       T                   �5@*��Q@             @R       S                    @|%��b�?             @������������������������       �                     �?������������������������       �                      @U       X                     @       @             @V       W                    �?      �?              @������������������������       �                     �?������������������������       �                     �?Y       Z                     @      �?              @������������������������       �                     �?������������������������       �                     �?\       k                     @u���9@             >@]       b                    �?��̎�@             .@^       a                    @���G�?             @_       `                    @�Z���?             @������������������������       ��c�����?             @������������������������       �                     �?������������������������       �      �?              @c       f                    �?|R��>@              @d       e                   �7@�c�����?             @������������������������       �                     @������������������������       �                     �?g       h                    @      �?             @������������������������       �                      @i       j                    @      �?              @������������������������       �                     �?������������������������       �                     �?l       m                    �?Lִ�e�?             .@������������������������       �                     *@������������������������       �      �?              @o       t                   �<@U���v @             5@p       s                    @z&F�Y�?             @q       r                    �?|%��b�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @u       v                    @�1H����?             0@������������������������       �                     &@w       z                   �?@|���7��?             @x       y                    @      �?              @������������������������       �                     �?������������������������       �                     �?{       |                    A@|%��b�?             @������������������������       �                      @������������������������       �                     �?�t�b�values�hhK ��h��R�(KK}KK��hV�B�Y         @      6@      4@       @      $@       @      @      @      5@      �?      9@      ,@       @       @      �?       @      �?       @      *@      @      @       @       @              0@      4@              "@               @              (@              6@       @                                                               @      @              �?              (@      4@              "@                               @              6@                                                                       @      @                               @      4@              "@                               @              @                                                                                                               @       @                                                              @                                                                                                                                                                                      @                                                                                                               @       @                                                              @                                                                                                              @      2@              "@                               @                                                                                                                              @      @              "@                               @                                                                                                                              �?      @                                               @                                                                                                                                      �?                                               @                                                                                                                                                                                       @                                                                                                                                      �?                                                                                                                                                                              �?      @                                                                                                                                                                                       @                                                                                                                                                                              �?      �?                                                                                                                                                                               @                      "@                                                                                                                                                              �?                      @                                                                                                                                                              �?                      @                                                                                                                                                              @      ,@                                                                                                                                                                               @      @                                                                                                                                                                              �?      @                                                                                                                                                                              �?      �?                                                                                                                                                                              �?      "@                                                                                                                                                                              �?      @                                                                                                                                                                                      @                                                                                                                                                                              @                                                                      0@                                                                       @      @                              @                                                                      @                                                                       @      @                                                                                                                                                                               @                                      @                                                                      @                                                                              @                              �?                                                                      @                                                                              @                                                                                                      �?                                                                               @                                                                                                      �?                                                                              �?                                                                                                                                                                                      �?                              �?                                                                       @                                                                              �?                                                                                                      �?                                                                                                              �?                                                                      �?                                                                              �?                               @                                                                                                                                                                                      �?                                                                      *@                                                                                                                                                                                       @                                                                                                              �?                                                                      @                                                                                                              @                                       @              $@                       @                                                                                      �?              @                                                      "@                                                                                                                              �?                                                      @                                                                                                                              �?                                                      @                                                                                                                                                                                      @                                                                                                                               @                                                      @                                                                                                                              �?                                       @              �?                       @                                                                                      �?                                                                                               @                                                                                      �?                                                                                                                                                                                      �?                                                                                               @                                                                                                      �?                                       @              �?                                                                                                                                                                                      �?                                                                                                                              �?                                       @                                                                                                                                                                                      �?                                                                                                                                              �?                                      �?                                                                                                                                       @      @               @      �?       @      �?      @      "@      �?      @      (@       @       @      �?       @      �?       @      *@      @               @      �?       @      @                      �?       @      �?      @      "@              @                       @      �?       @      �?              *@      @               @              @      @                               @              @      �?              @                              �?       @      �?                      @               @                                                       @               @                       @                                              �?                                       @                                                       @                                                                                      �?                                                                                              �?                                                                                      �?                                                                                              �?                                                                                                                                                                                                       @                       @                                                                                       @                                                                                               @                                                                                                                                                               @                                                                                                               @                                                                                                                                                                                       @                                                                       @                                                                                                                              @      @                                              �?      �?              �?                              �?       @                              @                              @       @                                                                                                      �?       @                                                              @       @                                                                                                      �?                                                                      @       @                                                                                                                                                                              @                                                                                                                                                                                      @       @                                                                                                                                                                              �?                                                                                                                                                                                      @       @                                                                                                                                                                              �?      �?                                                                                                                                                                               @      �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                               @                                                                      �?                                              �?      �?              �?                                                                      @                                                                                              �?                                                                                       @                                                                                              �?                                                                                                                                                                                                                                                                               @                                      �?                                              �?                      �?                                                                      �?                                      �?                                                                                                                                              �?                                                                                                                                                                                      �?                                      �?                                                                                                                                                                                                                                      �?                      �?                                                                                                                                                              �?                                                                                                                                                                                                              �?                                                                                                      �?      @                      �?              �?               @                                       @                                      *@      �?                              �?       @                      �?              �?              @                                       @                                              �?                                       @                                      �?              @                                                                                                                              �?                                                      @                                                                                                                              �?                                                      @                                                                                                                                                                                      �?                                                                                                                              �?                                      �?                                                                                                                                      �?                              �?                              @                                       @                                              �?                                                                                              @                                                                                      �?                                                                                              @                                                                                                                                                                                                                                                                              �?                              �?                              �?                                                                       @                                                                                                                                                                                       @                                                                              �?                              �?                                                                                                                                                                                      �?                                                                                                                                                      �?                                                                                                                                                                                              �?                                                      �?                                                                              *@                                                                                                                                                                                      *@                                              �?                                                      �?                                                                                                                                               @                              �?              �?              (@       @                                       @                                      �?                               @                                              �?                                                               @                                                                       @                                              �?                                                                                                                                                                                      �?                                                                                                                                       @                                                                                                                                                                                                                                                                                                       @                                                                                                      �?                              (@       @                                                                              �?                                                                                              &@                                                                                                                                                      �?                              �?       @                                                                              �?                                                              �?                                                                                                                      �?                                                                                                                                                                                      �?                                                              �?                                                                                                                                                                                                                      �?       @                                                                                                                                                                                       @                                                                                                                                                                              �?                                                                                        �t�bub�_sklearn_version��1.1.0�ub.