��2K      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C�                                                                	       
                                                               �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K
�
node_count�KW�nodes�hhK ��h��R�(KKW��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B         "                    �?���e��?�             c@                            �?�������?0             H@                           >@46<�R�?             9@                           @P���� �?             7@������������������������       �                     ,@                           �?X�<ݚ�?	             "@������������������������       �                     @       	                   �6@{�G�z�?             @������������������������       �                      @
                          �7@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           A@      �?              @������������������������       �                     �?������������������������       �                     �?                           7@L$e?���?             7@                           �?�|�j��?             .@                           �?      �?              @                          �4@�q�q�?             @������������������������       �                      @������������������������       �                     �?                          �3@z�G�z�?             @������������������������       �                      @                          �5@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?                             @:/����?             @������������������������       �                      @                           �?���Q��?             @������������������������       �                     @������������������������       �                      @        !                     @      �?              @������������������������       �                      @������������������������       �                     @#       0                    @n�����?i            @Z@$       -                    @�q�q�?             8@%       &                    �?�eP*L��?             6@������������������������       �                     (@'       *                    5@���Q��?
             $@(       )                      @      �?              @������������������������       �                     @������������������������       �                     �?+       ,                    @      �?              @������������������������       �                     �?������������������������       �                     �?.       /                     �?      �?              @������������������������       �                     �?������������������������       �                     �?1       J                    @T�Xnt�?Q            @T@2       G                     @��Z�O{�?9            �L@3       8                   �4@4F�b-�?&             C@4       7                   �0@HP�s��?             9@5       6                    �?���Q��?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     4@9       B                    @ƵHPS!�?             *@:       ;                   �5@{�G�z�?             @������������������������       �                     �?<       A                   �8@      �?             @=       @                    �?�q�q�?             @>       ?                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?C       F                    �?      �?              @D       E                    @���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @H       I                    �?p�ݯ��?             3@������������������������       �                     (@������������������������       �                     @K       P                     �?      �?             8@L       O                    9@{�G�z�?             @M       N                   �4@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @Q       R                    @��y4F�?             3@������������������������       �                     0@S       T                   �:@VUUUUU�?             @������������������������       �                     �?U       V                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�t�b�values�hhK ��h��R�(KKWKK��hV�B�3        2@      �?      ,@       @      @      �?      �?     �@@      8@      @      @      @      :@      @       @      @       @       @      �?       @               @              @      �?                               @      �?      @      8@      @              @                      �?                                              �?                               @      �?      �?      4@                                                                                                                               @      �?              4@                                                                                                                                                      ,@                                                                                                                               @      �?              @                                                                                                                                                      @                                                                                                                               @      �?               @                                                                                                                               @                                                                                                                                                              �?               @                                                                                                                                      �?                                                                                                                                                                       @                                                                                              �?                                              �?                                                                                                      �?                                                                                                                                                                                                      �?                                                               @               @              @                                                       @      @      @              @                      �?       @               @              @                                                              @                      @                      �?                                                                                                      @                      @                      �?                                                                                                                               @                      �?                                                                                                                               @                                                                                                                                                                              �?                                                                                                      @                      �?                                                                                                                               @                                                                                                                                                       @                      �?                                                                                                                              �?                      �?                                                                                                                              �?                                                       @               @              @                                                                                                                       @                                                                                                                                                                       @              @                                                                                                                                                      @                                                                                                                                       @                                                                                                                                                                                                                               @              @                                                                                                                                       @                                                                                                                                                                      @                                              0@      �?      (@       @                      �?     �@@      8@      @       @      @       @               @               @       @                      �?                                      �?              3@      �?       @                                                                              �?                                                      3@      �?      �?                                                                                                                                      (@                                                                                              �?                                                      @      �?      �?                                                                              �?                                                      @                                                                                                                                                      @                                                                                              �?                                                                                                                                                                                                                      �?      �?                                                                                                                                                      �?                                                                                                                                              �?                                                                                                                              �?                              �?                                                                                                                                                      �?                                                                                                                      �?                                                                                                      0@              (@       @                             �@@      @       @              @       @               @               @       @                              (@                                     �@@      @       @               @                       @                      �?                                                                      :@      @       @               @                       @                      �?                                                                      7@       @                                                                                                                                              @       @                                                                                                                                              �?                                                                                                                                                       @       @                                                                                                                                              4@                                                                                                                                                      @      @       @               @                       @                      �?                                                                                                       @                       @                      �?                                                                                                      �?                                                                                                                                                      �?                       @                      �?                                                                                                                               @                      �?                                                                                                                              �?                      �?                                                                                                                              �?                                                                                                                                                                              �?                                                                                                                              �?                                                                                                                              �?                                                                                                                      @      @       @                                                                                                                                      @               @                                                                                                                                                       @                                                                                                                                      @                                                                                                                                                              @                                                                                                      (@                                      @                                                                                                              (@                                                                                                                                                                                              @                                                                                              0@                       @                                                              �?       @                               @      �?                                       @                                                                      �?                               @                                               @                                                                      �?                                                                                                                                                      �?                                                                               @                                                                                                                                                                                                                                                               @                      0@                                                                                      �?      �?                                      �?              0@                                                                                                                                                                                                                                              �?      �?                                      �?                                                                                                      �?                                                                                                                                                              �?                                      �?                                                                                                              �?                                                                                                                                                                                              �?        �t�bub�_sklearn_version��1.1.0�ub.