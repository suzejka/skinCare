��v      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K
�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C�                                                                
                                                                                                  �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K	�
node_count�Ky�nodes�hhK ��h��R�(KKy��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�Bx         0                    �?�?CV�@�             c@                          �6@k=B��r@0             H@                          �4@JYS��@!            �@@                          �3@��Vw@             2@       
                    �?�v���?
             $@                           �?�c�����?             @������������������������       �                      @       	                   �1@      �?              @������������������������       �                     �?������������������������       �                     �?                            �?_�z|�X�?             @������������������������       �                     @                           �?|%��b�?             @������������������������       �      �?              @������������������������       �                     �?                           @�1H����?              @                           �?�9>����?             @������������������������       �                     �?������������������������       �V�T����?             @������������������������       �                     �?                           @�Du�q@             .@                             @�t�I�|�?	             "@                           �?��&��?             @������������������������       �                      @������������������������       �                     @                           �?�c�����?             @������������������������       �                     @������������������������       �                     �?                           �?|%��b�?             @������������������������       �                     @������������������������       �                      @        -                    >@��qa@             .@!       (                     �?�)���?             &@"       %                    @|���7��?             @#       $                   �7@      �?              @������������������������       �                     �?������������������������       �                     �?&       '                   �:@|%��b�?             @������������������������       �                     �?������������������������       �                      @)       ,                    @|%��b�?             @*       +                     @      �?             @������������������������       �|%��b�?             @������������������������       �                     �?������������������������       �                      @.       /                   �@@�c�����?             @������������������������       �                     �?������������������������       �                     @1       >                     �?�Օ�H�	@i            @Z@2       9                    @�F�Ze�?             3@3       8                    @܂��D��?             ,@4       5                    6@���q"
�?             *@������������������������       �        
             $@6       7                    �?|%��b�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?:       =                    9@z&F�Y�?             @;       <                   �4@|%��b�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @?       ^                    @���U'@V            �U@@       M                    @8t��n@5            �J@A       F                     @}�-j� @             :@B       E                     �?�v���?
             $@C       D                   �2@_�z|�X�?             @������������������������       ��c�����?             @������������������������       �                      @������������������������       �                     @G       H                    @      �?             0@������������������������       �                      @I       J                   �1@���'���?             ,@������������������������       �                      @K       L                    �?      �?             (@������������������������       ����'���?             @������������������������       ���&��?             @N       U                    �?]��[T @             ;@O       T                     @BL�F�0�?             0@P       S                    3@JQe1���?             ,@Q       R                   �1@      �?             @������������������������       ��c�����?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @V       [                    @6�DmU��?             &@W       Z                    @h���\�?             @X       Y                    4@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?\       ]                    <@c�YB�d�?              @������������������������       �                     @������������������������       �                     �?_       b                   �4@lh#2@!            �@@`       a                   �1@V�-���?             0@������������������������       �                     @������������������������       �        
             $@c       r                   �8@Ji��G@             1@d       g                     �?EA��W�?             *@e       f                    @������?             @������������������������       �                      @������������������������       �                     @h       o                    @���V��?             @i       l                    @      �?             @j       k                   �5@      �?              @������������������������       �                     �?������������������������       �                     �?m       n                    7@      �?              @������������������������       �                     �?������������������������       �                     �?p       q                   �7@      �?              @������������������������       �                     �?������������������������       �                     �?s       v                   �:@       @             @t       u                    @      �?              @������������������������       �                     �?������������������������       �                     �?w       x                    <@      �?              @������������������������       �                     �?������������������������       �                     �?�t�b�values�hhK ��h��R�(KKyKK��hV�B�V         @      6@       @       @      @      @       @      @      �?       @      @      �?      2@       @       @      @      �?      �?      ,@      @      �?      8@      0@               @               @      �?      @       @      @              �?      @                       @       @      @                      @      @               @                       @               @              @       @                              @                       @              @                      @                      �?                       @                              �?      @                                                                      @                      @                      �?                       @                                      @                                                                      @                                              �?                                                              �?                                                                      @                                                                                                                                                                                       @                                                                                                              �?                                                                      �?                                                                                                                                                                                      �?                                                                                                              �?                                                                                                                                               @                                      @                                                                                                                      �?                                                              @                                                                                                                                               @                                                                                                                                                              �?                      �?                                                                                                                                                              �?                      �?                                                                                                                                                                                                                      �?                                                                              �?                      @                                                                              �?                                                                                                      @                                                                                                                                                                                      �?                                                                              �?                                                                                                      @                                                                                                                                                              �?                                                                                       @              @      @                              @                       @                                                                                                       @              @      @                                                                                                                                                               @                      @                                                                                                                                                               @                                                                                                                                                                                                              @                                                                                                                                                                              @      �?                                                                                                                                                                              @                                                                                                                                                                                              �?                                                                                                                                                                                                                      @                       @                                                                                                                                                              @                                                                                                                                                                                                               @                                                                                                              �?                      @              �?                                       @      �?                              @              �?                                              �?                                                                               @      �?                              @              �?                                              �?                                                                                      �?                               @              �?                                              �?                                                                                      �?                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                       @              �?                                                                                                                                                                                      �?                                                                                                                                                                       @                                                                                                                                               @                                      @                                                                                                                                               @                                       @                                                                                                                                              �?                                       @                                                                                                                                              �?                                                                                                                                                                                                                               @                                                                                      @              �?                                                                                                                                                                                      �?                                                                                                                                                                      @                                                                                                                               @      4@       @      @       @                      �?      �?      �?      �?      �?      2@                              �?      �?       @      �?      �?      6@      0@       @                                                              �?                                                              �?      �?                              ,@                                                                                                                                              �?      �?                              (@                                                                                                                                                      �?                              (@                                                                                                                                                                                      $@                                                                                                                                                      �?                               @                                                                                                                                                                                       @                                                                                                                                                      �?                                                                                                                                                                              �?                                                       @                                                              �?                                                                                                       @               @                                                              �?                                                                                                                                                                                      �?                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                               @                      4@       @      @       @                      �?              �?      �?      �?      2@                                               @      �?      �?       @      0@              4@      �?      @       @                                              �?      �?      (@                                               @              �?              @              $@              @                                                                      �?                                               @                              @               @              @                                                                      �?                                                                              @               @              @                                                                      �?                                                                                                              @                                                                      �?                                                                                               @                                                                                                                                                                                                                                                                                                                                                              @               @                                                                                                                                       @                                               @                                                                                                                                                                                      @                                                                                                                                       @                                                                                                                                                                                       @                                              @                                                                                                                                      @                                              @                                                                                                                                      @                                               @                                                                                                                                      @                                              $@      �?               @                                              �?      �?      &@                                                              �?                              @                       @                                                              &@                                                                                              @                                                                                      &@                                                                                              @                                                                                      @                                                                                              �?                                                                                      @                                                                                               @                                                                                                                                                                                                                                                                               @                                                                                                                       @                                                                                                                                                              @      �?                                                              �?      �?                                                                      �?                                      �?                                                                      �?                                                                      �?                                                                                                              �?                                                                      �?                                                                                                              �?                                                                                                                                                                                                                                                              �?                                      �?                                                                                                                                                                              @                                                                      �?                                                                                                              @                                                                                                                                                                                                                                                              �?                                                                                                                      �?      @                              �?              �?                      @                                                      �?               @      (@                                                                                                                                                                              @      $@                                                                                                                                                                              @                                                                                                                                                                                              $@                      �?      @                              �?              �?                      @                                                      �?               @       @                              @                                                                      @                                                                       @       @                               @                                                                      @                                                                                                               @                                                                                                                                                                                                                                                              @                                                                                                              �?                                                                      �?                                                                       @       @                                                                                                      �?                                                                       @      �?                                                                                                      �?                                                                      �?                                                                                                                                                                                      �?                                                                                                              �?                                                                                                                                                                                                                                                              �?      �?                                                                                                                                                                                      �?                                                                                                                                                                              �?                                      �?                                                                                                                                                      �?                              �?                                                                                                                                                                                                                                                                                                                                              �?                      �?                                      �?              �?                                                                              �?                                              �?                                      �?                                                                                                                                                                                      �?                                                                                                                                              �?                                                                                                                                                                                                                                              �?                                                                              �?                                                                                                      �?                                                                                                                                                                                                                                                                      �?                        �t�bub�_sklearn_version��1.1.0�ub.