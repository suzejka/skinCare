���0      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K
�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C@                                                         �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K	�
node_count�K_�nodes�hhK ��h��R�(KK_��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B�         ,                    @7j�P�e�?s            �\@                             @r�q��?0             H@                          �4@��2Tv�?             >@                           �?ffffff�?             4@                          �2@      �?             @������������������������       �                      @������������������������       �      �?              @                            �?     @�?             0@	                           2@      �?              @
                           �?�Q����?             @������������������������       �                      @������������������������       �VUUUUU�?             @������������������������       ��q�q�?             @                           �?      �?              @                           @r�q��?             @������������������������       �                      @������������������������       �      �?             @������������������������       �      �?              @                            �?{�G�z�?
             $@                           �?�$I�$I�?             @                           �?z�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �      �?              @                           �?VUUUUU�?             @������������������������       �      �?              @������������������������       �                     �?       +                   �6@<ݚ�?             2@       $                    �?     @�?             0@       !                    3@      �?              @                           �1@�q�q�?             @������������������������       �                     �?������������������������       �                      @"       #                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @%       &                    �?      �?              @������������������������       �                     �?'       (                    �?������?             @������������������������       �                     �?)       *                   �2@�8��8��?             @������������������������       �      �?              @������������������������       �      �?             @������������������������       �                      @-       P                     @�(M?�e�?C            �P@.       K                   �5@	�̮�r�?3            �I@/       F                   �4@�<DC%�?.             G@0       =                    �?��r._�?)            �D@1       8                     �?�p=
ף�?             4@2       7                    @��S���?             .@3       6                    @*x9/��?             ,@4       5                    �?X�<ݚ�?	             "@������������������������       ��q�q�?             @������������������������       �      �?             @������������������������       ��Q����?             @������������������������       �                     �?9       :                    @�Q����?             @������������������������       �      �?              @;       <                    2@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @>       A                    @Tg�x�P�?             5@?       @                    �?��Q��?
             $@������������������������       ��8��8��?             @������������������������       �      �?             @B       E                   �2@�C��2(�?             &@C       D                   �0@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @G       H                    @{�G�z�?             @������������������������       �                      @I       J                    �?�q�q�?             @������������������������       �      �?              @������������������������       �                     �?L       O                    �?���Q��?             @M       N                    @�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                      @Q       V                    �?     ��?             0@R       U                    �?x�5?,�?	             "@S       T                    �?      �?              @������������������������       �      �?             @������������������������       �      �?             @������������������������       �                     �?W       ^                   �5@������?             @X       ]                   �2@�8��8��?             @Y       Z                    �?      �?             @������������������������       �                     �?[       \                    @�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�t�b�values�hhK ��h��R�(KK_KK��hV�B�        @      1@     �B@      <@      &@       @      @      &@      @      @      @      *@      @       @      @      "@              �?      @       @      @              �?      "@                       @      @      @              �?      "@                              �?       @              �?                                               @                                                      �?                      �?                               @      @      �?                      "@                       @       @      �?                      @                              �?      �?                      @                                                               @                              �?      �?                      �?                       @      �?                                                               @                              @                              �?                              @                                                               @                              �?                              @                              �?                              �?              �?      @      @      �?                                              @       @      �?                                              @      �?                                                       @      �?                                                       @                                                                      �?      �?                                      �?      �?      �?                                              �?              �?                                                      �?                                              @      @              @               @      @              @      �?              @               @      @              �?                      �?               @      @                                      �?               @                                              �?                                                                               @                      �?                                              @              �?                                                                                                              @              @      �?              @                                                              �?                                      @      �?              @                                      �?                                                               @      �?              @                                              �?              �?                                       @                       @                                               @                                                              *@      >@      .@      @                       @              &@      ;@      "@       @                       @               @      ;@      @       @                       @               @      9@      @       @                                      @      $@      @      �?                                       @      $@      @                                               @      "@      @                                              �?      @       @                                                       @      �?                                              �?      @      �?                                              �?      @      �?                                                      �?                                                      @              �?      �?                                      �?              �?                                               @                      �?                                      �?                                                              �?                      �?                                      @      .@       @      �?                                       @      @       @      �?                                              @       @      �?                                       @       @                                                      �?      $@                                                      �?      @                                                              @                                                      �?                                                                      @                                                               @      �?                               @                       @                                                                      �?                               @                              �?                              �?                                                              �?              @               @                                              �?               @                                                              �?                                              �?              �?                                               @                                                               @      @      @      @                                      �?              @      @                                      �?              @      @                                      �?              �?       @                                                       @       @                                                              �?                                      �?      @      @                                              �?       @      @                                              �?       @      �?                                              �?                                                                       @      �?                                                      �?      �?                                                      �?                                                                       @                                                      �?                                        �t�bub�_sklearn_version��1.1.0�ub.