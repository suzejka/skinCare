��e&      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K
�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C@                                                         �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K	�
node_count�KI�nodes�hhK ��h��R�(KKI��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B�                             �?.���@s            �\@                           �?���� �?             ;@                          �2@       @              @                           �?h���\�?             @������������������������       �                     �?                          �1@      �?              @������������������������       �                     �?������������������������       �                     �?	       
                    �?�Z���?             @������������������������       �      �?              @������������������������       �                     @                           �?��l�?             3@������������������������       �                     @                           @JQe1���?             ,@                           �?V�-���?              @                           3@|%��b�?             @������������������������       �                     �?������������������������       �                      @                            �?�Z���?             @������������������������       �                     @������������������������       �      �?              @������������������������       �                     @       @                    @h$�w!5�?X             V@       5                    @� K���?H             R@       *                    @�;�t�m�?4             J@       #                     �?"�\�?!            �@@                            @w���Q�?             3@                            �?�Z���?
             $@                           6@|%��b�?             @������������������������       �|%��b�?             @������������������������       �                     @������������������������       �                     @!       "                    �?|%��b�?	             "@������������������������       �|%��b�?             @������������������������       ����V��?             @$       )                    @!,�Wj}�?             ,@%       &                     @҂�26��?
             $@������������������������       �      �?             @'       (                   �4@�c�����?             @������������������������       �                      @������������������������       �      �?              @������������������������       �      �?             @+       4                   �5@vׯD�"�?             3@,       3                    �?M�)9��?             2@-       .                      @��Ȓ���?             &@������������������������       �                     @/       2                   �3@|%��b�?             @0       1                     @��&��?             @������������������������       ��c�����?             @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?6       ;                    �?x1���?             4@7       8                    @��Ȓ���?             &@������������������������       �                      @9       :                     �?|%��b�?             @������������������������       �                     �?������������������������       �      �?              @<       ?                    @�t�I�|�?	             "@=       >                     �?�Z���?             @������������������������       �|%��b�?             @������������������������       �                      @������������������������       ��c�����?             @A       D                   �2@��e����?             0@B       C                    �?      �?              @������������������������       �                     �?������������������������       �                     �?E       H                   �4@�9>����?             ,@F       G                    �?�c�����?              @������������������������       �                      @������������������������       �|%��b�?             @������������������������       �                     @�t�b�values�hhK ��h��R�(KKIKK��hV�B@        �?      .@      <@      �?      E@      :@      �?      �?      �?       @              �?              .@      �?      �?      �?                      �?              @      �?      �?      �?                                              �?      �?                                                              �?      �?                                              �?                                                              �?              �?                                                                                      �?              @                                              �?              �?                                                              @                               @                              &@                              @                                                              @                              &@                              @                              @                               @                              �?                                                              �?                               @                                                              �?                              @                                                              @                              �?                              �?                                                              @                              @      <@              E@      &@                              @      .@              D@      $@                              @      @              A@      @                              @      @              2@      @                               @      @              (@      �?                                       @               @                                               @              @                                               @              �?                                                              @                                                              @                                       @       @              @      �?                              �?                       @                                      �?       @               @      �?                              @                      @      @                              @                      @      �?                              @                      @                                                              @      �?                                                       @                                                              �?      �?                               @                               @                                                      0@      @                                                      0@       @                                                      "@       @                                                      @                                                              @       @                                                      @       @                                                      @      �?                                                              �?                                                      �?                                                              @                                                                      �?                                      &@              @      @                                      "@               @                                               @                                                              �?               @                                                              �?                                              �?              �?                                               @              @      @                                      �?              @                                              �?               @                                                               @                                              �?                      @                                      *@               @      �?                                      �?                      �?                                      �?                                                                                      �?                                      (@               @                                              @               @                                               @                                                              @               @                                              @                                        �t�bub�_sklearn_version��1.1.0�ub.