���?      �!sklearn.neighbors._classification��KNeighborsClassifier���)��}�(�n_neighbors�K�radius�N�	algorithm��auto��	leaf_size�K�metric��	minkowski��metric_params�N�p�K�n_jobs�N�weights��uniform��n_features_in_�K�outputs_2d_���classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C�                                                                	       
                                                               �t�b�_y�hhK ��h��R�(KMI��h �i4�����R�(Kh$NNNJ����J����K t�b�B$=                                                                    	                                                                                                                                                                     	                              
                                                                                                     
                                              	                                      
                                                                    	                                                                                 	                   
                                                                                                                                                                                                                                                                   	                             	                                                                                                                                                                                                                                                       	                                                                                                  	                                                                                                         
                                                                                                                                              
                  	                                                                                                                 	         
                                                                                                                                                                              
             
                                           	                                                                                       	         
               	                                                                                                                                                                                
         
                                  	                                                      	            	                                    
         
                                                                                
            
                	                                                                                    	                                                                                                                                                                                      	         
                            	                                                                                                  
                    
                                    	                                    	                                                                                                                          	                
                                   	                                                                                                                                                                               
                                                                                                                                         
                         	                                                                                                                         	                                                                               
                                 	                                        
                                                  	                       
                   
         
                                             	                               
      	                                           	                                          	                   
   
                                         
                                                                                                                                 	                                                                            
         	                              	                                                   
                                                                          
         
                                                                                                          	            	                                                                                                                                     
                                             	                                                                                                	                                     	                                          
                                                                                                                                                          
                                                           
                   
                                                                                                                          	                                                                                                                                                                                                                                              
                                                                                                                                        
                                                                               	                                                                                              
                                                     	            
                                     
                                                                                                                                                                                                                                                                                                                                                                  	                     
                                                                                    
                         
                                     	                        	                                                                                                                                                                                                  
            	                   	                
      	            
                                                                                                                                                                                        	                                    
                                                         	                                                    
                                               	                                                    	   
                                                       
                                                                                              	         	                                                                                                                                                                                       	                                                                                                               
                                                                                               
                          	      
                                          	                       
   
                                      
                                                                                             	                                                                                                                                                    
                                                         	                                                                                                                     
                                                                                                                                                             	            	                                                                                          	                                                                                
            	                                                	                                                                                          
               
               	                                                                                                                                                                                                          	         
                                                                                                                                                                                                                                                               	                  
                                       	   
                                             	                                                                                                                      	                                                        	                                                                                                                	                                                  	                                                                           	                                             
                                                          
                                                                                 
   	               
                                                                                               	                                                                                                                                    
            	                             	                     
                                                                       
                                                                       	                            
                                                                                                                                                                                                                               
                                        	                            	                                                                                                                                                            	                                                      	                                                                    
      
                        
                                                                          
                      	                                                       	                                                                                                                                    
                             	                                                        
                                                                                                                                                                                                                           
                                                                                                                                                     	         
      
                                                       
      	   
       
                                                                                                    
                                                                                                                                          
                         	                                                                                                                               �t�b�effective_metric_params_�}��effective_metric_��	euclidean��_fit_method��kd_tree��_fit_X�hhK ��h��R�(KMIK��h#�Bhc                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         "                                                                                                                                                                                                                                                           #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    $                                                                                                                                                                                                                                                                                                                                                                          %                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          %                                                                                                                                                                                                                                                          "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             #                                                                                                                                                                                                                                                                                                                                                                                                                                                                               !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 #                                                                                                                                                                                                                                                                                                                                                                                                                                                     "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 	                                                                                                                   !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    %                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       $                                                                                                                                                                                                                                                           	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            "                                                                                                                                                                                                                                                                                                !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             #                                                                                                                                                                                     "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 "                                                                                                            !                                                                                                                                                                                                                                                       %                                                                                                                                                                                      #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               $                                                                      !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              	       $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     !                                                                                                                                                                                   #                                                                                                                                                                                                                                                                                                                                                                        $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 $                                                                                                                                                                                                                                                                                                       #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "                                                                                                          !                                                                                                                                                                                                                                                                                                                                       #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       !                                                                                                                                                                                                                        $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      $                                                                                                                                                    !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            #                                                                                                                                                                                                                                                                                                   "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   !                                                                                                             !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "                                                                                                                                                                                                                                                                                                   %                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               %                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  !                                   !                                    !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               	                                                                                                                                                         #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           	                                                                              "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ��       �t�b�n_samples_fit_�MI�_tree��sklearn.neighbors._kd_tree��newObj���hB�KDTree�����R�(hhK ��h��R�(KMIK��h �f8�����R�(Kh$NNNJ����J����K t�b�Bhc       @                      @      6@              �?      �?              8@              �?              @      3@      @                              1@       @      �?      @              1@                      @      @      0@              �?      �?      @      ;@              �?              @      8@      @      �?      �?      @      >@                       @              4@      �?      �?       @      @      2@      @      �?      �?       @      =@      @      �?      @      �?      2@       @               @      "@      7@       @      �?       @      @      7@       @              @              2@      �?                      @      7@      @      �?      �?              0@                       @              :@       @      �?       @      @      >@      �?      �?      @      @      9@      �?      �?              @      <@       @              @              5@              �?      @      @      <@      �?                              3@      @      �?      �?      @      6@      �?      �?      @              5@      �?      �?              @      8@       @      �?       @      @      6@      @      �?      @      @      4@       @                              3@              �?       @      @      2@      �?              @      @      4@                       @              4@                      @       @      1@              �?      @      @      2@       @      �?                      9@      �?              @              4@      �?              @      @      9@                                      3@      @                       @      0@       @              @      @      ;@      �?      �?                      9@                      @      @      =@              �?      �?      @      ;@      @      �?      �?              6@       @              �?      @      9@                      �?      @      8@                      @      @      ;@              �?      �?      @      4@      @      �?      �?      @      0@                                     �@@      @              �?              :@      @      �?      �?              4@      @              �?      @      3@       @              @      @      =@      @      �?      �?      @      8@      �?                              7@      @              @              7@      �?      �?       @      @      4@              �?       @              0@      @               @      @      0@      @                       @      8@              �?      �?      @      6@              �?      �?      @      ;@      @              @      @      6@                      �?      @      2@              �?      @      @      4@                       @      @      3@              �?      @       @      7@       @      �?       @      @      3@      @              @      @      6@      @               @              ;@       @      �?      @      @      1@      �?              @              5@      �?      �?       @              1@      @      �?      @      @      A@                      �?      @      @@      @      �?      @       @      3@      @      �?      @      @      7@      @      �?       @      @      0@      �?      �?      @              0@      �?      �?               @      1@              �?      �?      @     �A@       @              @      @      6@      �?              @              8@      @      �?      @      @      4@      �?      �?      @       @      3@       @      �?      @              7@      @              @       @      2@      @      �?      �?      @      4@      @      �?      �?       @      8@      @      �?              @      5@      �?               @      @      6@                      @       @      8@       @              @      @      8@       @               @      @      9@      �?              @              2@       @              @      @      6@                      �?      @      3@      @              @      @      1@                      @      @      2@      �?      �?      @              5@                      �?      @      5@              �?      �?      @      =@      �?      �?                      4@                      �?      @      3@      @              �?      �?      B@      @      �?       @              :@       @              @      @      <@                      �?      @      5@      @      �?      @              7@      @              �?       @      3@      @              @              0@                      @              3@      @      �?      @              2@      @      �?      �?      @      7@      �?      �?      �?      @     �B@      �?      �?      �?      @      4@                              @      1@              �?      @      @      4@                      @              3@       @              @              7@       @      �?      @       @      7@                      @      @      1@      @      �?      @              ;@      �?      �?                      1@      �?      �?      �?              2@      @              @      @      3@      �?              �?              9@       @      �?      @      @      7@                       @      @      7@      @      �?       @              :@      �?              @      @      >@      @              �?              2@      �?      �?      �?              1@      @              �?      @      ;@      �?      �?       @      @      2@      @                              3@      @      �?      �?              <@              �?       @              3@                      �?              0@              �?      @       @      =@      �?      �?      �?      @      4@      �?              @      @      3@                      @      @      1@              �?      @      @      9@      @                      @      7@      @      �?      �?       @      6@      �?      �?              @      2@      @              @      @      :@       @              @              0@              �?      @       @      9@       @      �?      @      @      2@      @              �?      @      6@      @               @              1@      @              �?      @      2@                      �?       @      4@      �?              @              9@              �?      @      @      9@              �?      @              8@                      @      @      8@                       @              4@      �?              @      @      1@      @               @              5@              �?              @      9@      �?               @      @      2@              �?      @      @      1@      @      �?      �?      @      0@              �?       @      @      1@      �?              @      @      6@      @               @      @      4@       @      �?       @      @      6@      @              @      �?      7@      @              @      �?      6@      @      �?      �?             �B@      @      �?      �?       @      8@      �?      �?      @       @      2@                      @              1@      @      �?       @      �?      2@      �?              �?      @      6@      �?      �?      @      @      5@      @              �?      @      A@                      @              4@      @      �?      �?      @      3@       @              @              3@      @      �?      @      �?      2@       @      �?      �?      @      ?@      �?      �?      �?      @      4@              �?      @      @      7@              �?              @      8@              �?      �?      @      1@      @      �?      @              8@      �?                              5@      @      �?      @              4@      �?      �?      �?      @      3@      �?      �?      �?              9@      @      �?      �?      @      2@                       @              7@              �?      �?      @      :@              �?       @      @      :@       @      �?      @      @      0@      @      �?      @              4@      �?              @              8@                              @      ;@       @      �?      @      @      2@      �?      �?       @      @      1@              �?      @              :@      �?              @      @      0@      �?              @      @      3@      �?                              2@      @      �?       @      @      :@      �?              @              7@              �?      @              ?@      @      �?      �?      @      2@      �?              @              4@      @      �?      �?      @      9@      @              @      @      6@              �?                      2@      �?      �?              @      <@      �?               @              4@       @      �?      @      @      3@      �?              �?      @      1@      �?              @              3@      @      �?              @      2@      �?      �?      @      @      8@       @              @              4@      @                       @      <@                      @              4@      @              @       @      3@      @      �?      �?      �?      8@                       @              2@              �?                      0@                      @              ;@       @              @              8@       @      �?              @     �A@              �?      @      @      4@              �?       @      �?      4@              �?      �?      @      9@              �?                      0@      �?      �?      @       @      >@       @              @      @      5@       @      �?                      3@       @      �?              @      0@                              @      7@       @              @      @      2@                      @      @      0@      @      �?      �?              6@              �?                      4@                      �?              5@              �?      �?      @      3@       @              @      @      0@       @      �?      �?      @     �A@              �?      �?      @      =@              �?       @              6@              �?       @      @      6@      �?      �?       @              =@       @      �?      @       @      3@      @              @      @      2@      @      �?      �?      @      5@      @      �?      �?              :@      @      �?       @      @      5@       @              @       @      4@                                      0@       @               @      �?      ?@      @                              6@              �?      @      @      5@       @      �?      @      @      :@      �?      �?      @              1@              �?              @      2@      @                       @      4@      �?                      @      0@      �?              �?       @      8@      �?      �?       @       @      6@      @      �?              @      7@                      �?              4@      �?      �?      �?              2@      �?              @              ;@      �?              @              1@      @      �?      �?              1@      @      �?      �?      @      6@      @      �?      �?      @      ?@       @              @      @      5@              �?      @      �?      5@                       @      @      4@              �?      �?              2@      �?      �?      @              6@      @      �?      @      @      6@      @      �?       @      @      5@      @      �?      @      @      5@      @              @      @      2@      �?               @       @      5@              �?      �?      @      3@      �?      �?                      :@      �?      �?      @              7@       @      �?      @              9@       @              �?       @      7@      �?                              2@              �?      �?              :@       @      �?      @              1@      �?      �?      @       @      8@      �?      �?      @      @      8@      @      �?      �?       @      @@      @      �?      �?              ?@                      �?      @      5@      @              �?      @      8@      �?              @      @      4@      �?      �?                      8@       @      �?      @       @      6@              �?              @      9@       @      �?      @       @      2@      �?      �?      @              7@      �?      �?                      1@       @      �?       @              6@                      @       @      2@              �?      @      @      :@      @              @      �?      :@      @              @              1@              �?      �?      @      9@      @      �?      @      @      4@      �?              @      @      4@       @              @      @      5@      �?      �?       @      @      >@      �?              @              0@      �?      �?      �?      @      0@      �?               @              4@                                      5@      �?      �?              @      6@      @      �?      @      @      8@       @      �?              @      ?@      �?      �?      @              4@      �?              @              5@       @              @              7@              �?               @      4@       @              @      @      6@      �?      �?       @      @      5@      �?              @              6@      @      �?      �?      @      1@      @      �?      �?       @      2@      @                       @      1@      �?      �?      @      @      4@      �?              �?      @      8@              �?              @      7@       @      �?      @      @      2@      @              �?              7@                      @      @      >@      �?      �?      @      @      ?@      @      �?       @      @      2@       @      �?      @      @      0@                       @              3@      �?      �?      @      @      7@      �?              @      @      7@      �?      �?       @      @      6@                      @      @      2@      @      �?      �?              ;@       @      �?      @              5@       @              @      @      6@       @                      @      2@      �?                      �?      2@      �?              @              3@              �?      �?              :@      �?              �?      @      9@      �?                      @      7@       @      �?      @              5@                      @      @      :@      �?              @              5@      �?               @       @      9@       @      �?      @      @      <@      @              �?              3@      �?      �?      �?       @      6@      @      �?      �?      @      9@      �?      �?      @              2@      �?      �?      @      �?      4@      �?               @              3@      @              �?              4@      �?              @              8@              �?      �?       @      8@       @              @              0@              �?      @      @     �A@      @              @      @      :@      @      �?      �?      @      :@      �?      �?      �?              3@       @      �?      @       @      2@      �?      �?      @      @      1@      @      �?       @      @      4@       @      �?      @      @      7@       @      �?      @              <@              �?      �?      @      3@              �?       @              2@      �?      �?      �?      @      ?@      @              �?      �?      ;@      �?      �?              @     �@@      @      �?              @      ;@      �?      �?      �?      @      2@      @      �?      �?      @      ;@      �?              @              :@      �?      �?      �?      @      >@              �?      @      @      2@       @      �?       @      @      3@                              @      >@      @      �?      �?              8@      @              �?              7@      �?              @              0@              �?      �?      @      ?@      �?      �?      @              2@      �?              �?       @      4@      �?      �?      @              9@      @              �?      @      ;@      @      �?      �?      @      4@              �?      @      @      =@      �?      �?      �?              :@      �?      �?       @              =@              �?      �?              5@      @              �?      @      4@      @              �?      @      ?@                       @      @      9@       @      �?      @      @      1@                      @              2@                                      <@       @              �?              2@      �?      �?      @      @      9@      �?              @      @      1@      �?      �?              @      3@       @              @      @      4@      @      �?      �?      @      >@      @      �?              @      :@              �?      @      �?      5@      @              @      @      0@      @      �?      @              2@      @              �?      @      :@      @                      @      7@                      �?       @      1@                      @      @      4@       @      �?      @              4@                       @              ;@       @      �?      @      "@      2@      @              @       @      1@      �?      �?                      3@              �?      @      @      2@              �?              @      5@      @                              4@                      @      @      2@      @              �?              8@      @      �?      @              :@      �?              @      �?      6@      @      �?      @              2@      �?      �?                      =@      @               @      @      1@       @              @      @      :@      �?      �?      @      �?      3@      �?              @      �?      2@              �?      �?      @      3@              �?      @      @      0@              �?              @      4@       @               @              1@      �?              @              5@      �?      �?      @              :@                      �?              6@                              @      5@      �?      �?      @      @      0@      @                              1@      �?      �?       @       @      5@      @      �?      @      @      6@      �?      �?      @              1@       @      �?       @      @      1@      @      �?      �?              3@      �?              @              <@                      �?      @      1@      @              @      �?      0@       @      �?      @      @      <@      @      �?      @      @      5@       @      �?      @              9@       @      �?       @      @      9@              �?      �?      @      8@      @              @              2@      @      �?      �?      �?      5@                      @      @      6@      �?                      @      @@              �?      �?      @      4@       @      �?                      5@                      @      @      4@      @              �?              3@       @      �?      @      @      7@       @              @      @      0@      �?               @      �?      8@      �?      �?      @              :@                      @              6@      �?      �?      @              4@      �?              @              3@      @      �?      �?      @     �A@      �?      �?                      6@      @      �?              @      8@      @      �?      �?       @      :@      �?              @              1@      @              @       @      2@      �?      �?      @      @      8@       @              @       @      1@              �?      �?       @      9@       @      �?      @      @      1@              �?      �?      @      ;@      �?      �?      @      @      1@      �?      �?      @              1@       @      �?      @      @      3@      �?                              2@      �?      �?       @              5@      �?              @      @      1@       @      �?      @      @      5@       @              @              0@      @              @              9@      @      �?       @              9@      �?      �?              @      5@              �?      @      @      1@      �?              @              7@      @               @              2@              �?       @      @      2@              �?      @       @      0@      @                       @      5@       @              @      @      3@      �?              @              3@      �?              @      @      4@      �?      �?       @              1@       @              @              >@      @                              :@              �?       @      @      8@      �?              �?              5@      @                      @      5@                       @              3@      @      �?                      6@      @      �?      �?      @      B@              �?       @      @      2@      @      �?       @       @      =@      @      �?      �?      @      9@       @      �?      �?              3@      �?              @       @      8@      �?      �?      @      @      1@      @      �?      @              9@              �?                      9@              �?      @      @      5@       @              @              2@      �?      �?      @      @      =@      @      �?              @      2@      @              @              5@      @      �?      �?              5@      �?              �?      @      8@      @              @      @      6@              �?      @      �?      2@      @      �?      �?       @      9@      @      �?      @              1@      @      �?      �?      @      2@       @      �?      @      @      5@              �?       @      �?      :@              �?                      9@       @               @              :@      �?              �?              2@       @              @      @      1@      �?      �?      @      @      9@      �?      �?      �?              7@      �?      �?      �?      @      8@              �?       @       @      1@       @      �?      @      @      0@      @              @              2@                      �?      @      7@       @               @              9@      �?              �?       @      :@      @              �?      @     �A@              �?      �?      @      1@      �?              @      @      5@       @              �?              5@      �?      �?               @      9@              �?      @      @      7@                      �?       @      6@      �?      �?                      @@              �?      �?      @      ;@       @              @      @      0@       @              @              1@       @      �?      @      @      3@              �?              @      A@       @              @      @      6@       @      �?      �?              9@      �?              @              6@              �?      �?      @      <@      @      �?                      2@      @      �?      @      @      5@      @      �?              @      6@       @              @      @      ;@      @               @              7@      �?              @       @      <@      @      �?      �?      @      6@       @              @              9@                       @              ;@      @      �?              @     �A@       @               @      @      0@      @      �?      �?      @      3@      �?      �?      @      @      4@      @              �?      @      7@              �?              �?      6@      @      �?      @              7@       @      �?      �?              2@      @              @              5@              �?      �?              1@                      @              1@                      @              1@      �?      �?      @      @      0@      @      �?      @      @      8@      @              �?              6@              �?              @      4@                      @      @      0@       @      �?      @       @      3@      @              �?              :@                      �?      @      5@                       @      @      6@              �?      @       @      2@      �?      �?      @              1@      �?      �?      �?      @      5@      @      �?      �?              <@      @      �?      �?      @      1@      �?      �?      @      @      6@       @              @              3@      �?              @              2@                      �?              3@                      @       @      2@       @      �?      @      @      8@      @              �?              8@                      @      @      5@       @      �?      @              6@       @      �?      @       @      5@       @      �?      @              6@      �?              �?              1@       @      �?      @      @      4@              �?      @      @      2@      @      �?       @      @      0@      �?      �?                      5@      @      �?              @      9@       @               @      @      9@      @              @      @      4@      �?                      @      1@      �?              @      @      5@      @               @      @      :@      �?              �?      @      5@      @              �?      @      :@      �?      �?      @              1@              �?      @              1@      @                      @      @@       @              �?      @      >@                      @              0@      �?              @      @      1@      @      �?      �?              ;@       @               @              4@      @              @      @      5@      @              �?      @      :@              �?      @      @      <@      @      �?      @       @      4@                              @      9@       @              @              4@              �?      @      @      0@              �?      �?              =@      �?      �?      @      @      4@      �?              @              1@       @              @       @      1@       @              @      @      1@      @               @              :@      @      �?      �?      @      4@              �?      �?      @      A@      �?      �?      @      @      6@                      @      @      3@       @      �?      @      @      1@      �?              @              2@      �?      �?      �?              5@      @                      @      =@       @              @              1@      @               @      @      1@              �?      @              3@                      �?      @      9@      �?      �?      @      @      1@      @              �?       @      ;@              �?      @      @      6@                      �?              2@      @      �?       @      @      ;@       @      �?      @      @      >@      @              @              6@              �?       @              2@      �?              @      �?      <@      �?              @      @      :@      @              @              5@                      @              1@       @      �?      @      @      @@              �?      @      @      3@       @      �?      @      @      3@      �?      �?              @      7@      @      �?      �?      @      :@      @      �?      �?      @      2@      @      �?      �?              3@       @      �?      �?      @      3@              �?      �?      @      7@       @              @      @      8@                       @      @      5@      �?               @              1@              �?      @      @      <@              �?      �?      @      1@      @      �?       @              9@              �?              @      3@       @      �?      @              2@      �?      �?      @              1@              �?      @      @      5@              �?      @       @      6@      @                              2@      @                      @      6@      �?      �?      �?      @      2@      �?              @              1@      �?      �?              @      B@              �?       @              ;@      �?      �?      @              5@      �?      �?      @              1@      �?      �?              @      4@      @              @      @      4@      @      �?      �?              8@      �?      �?       @      @      7@       @      �?      @      @      8@      �?              @              3@      �?              @              1@                       @              4@              �?       @              0@       @      �?      @              5@      �?      �?      @              6@                      @              0@              �?       @      @      4@       @      �?      @      �?      6@              �?      �?      @      1@      �?              @              1@                      @              2@       @              @              2@      @              @      @      5@              �?       @      @      2@                       @              @@      �?              @      @      0@      �?      �?       @              9@      �?              @              1@              �?       @       @      8@      �?              @              2@      �?      �?      @              3@                      @      @      8@      �?      �?      @      @      3@                      @              4@      �?              @      "@      3@       @              @              0@      �?              @      @      :@      �?      �?      @      @     �@@      �?              @              5@      �?      �?      @      @      0@      �?              @              2@      @                              <@      @      �?      �?      @      >@      @              �?      @      7@       @      �?      �?      �?      6@       @      �?              @      1@       @      �?                      =@                      @      @      8@      @              @              <@       @      �?      @      @      0@      @              @      @      4@              �?       @      @      6@      �?                              0@       @      �?              @      4@      @      �?              @      ;@      @      �?      �?      �?      8@      �?              @              2@      �?      �?                      9@      �?              �?       @      ?@      @      �?      @      @      8@      �?      �?      @       @      5@      �?      �?      �?       @      ;@      @      �?      �?              7@      �?      �?      @      @      6@      @                      @      8@      �?      �?      @       @      2@      �?      �?      @              =@      �?              @       @      8@       @      �?      �?      @      4@       @      �?      @       @      >@      @              �?      @      2@       @      �?      @              8@      @      �?      �?      @      <@      �?      �?       @      �?      8@      �?               @              0@                      @      @      1@       @      �?      @      @      1@      @               @       @      5@      @      �?      @      @      7@       @      �?      @      @      :@      �?              @      @      0@              �?      @      @      1@                      @      @      1@      �?              @      @      6@                       @      @      5@      �?              @      @      1@      �?              @              7@      @              �?      @      ;@       @      �?       @      @      ?@      �?               @      �?      6@              �?              @      6@      �?      �?      @              1@      @      �?      �?      @      8@              �?      �?      @      9@       @              @      �?      8@      @      �?      �?       @      <@      @              �?              3@      �?      �?      �?       @      >@      @               @      @      5@      �?               @      @      0@      @              @      �?      5@      �?              @              2@      @      �?       @      @      5@      @      �?      @      @      ;@      @      �?      @              5@              �?      @      @      8@      @      �?                      ;@      @                      @      2@              �?      �?       @      6@              �?      @      @      5@              �?      �?      @      4@      @      �?      �?      �?      8@      �?      �?      �?      @      :@      @               @      @      2@      �?              @              0@      @      �?      �?      @      4@              �?              @      8@      �?      �?      �?      @     �@@      �?      �?       @      @      5@      �?      �?              @      9@      �?      �?      @      @      9@       @      �?       @       @      :@              �?              @      6@      �?      �?      @      @      1@      �?              @      @      1@              �?      �?       @      8@       @              @      @      2@       @      �?                      6@      @      �?      �?      @      9@              �?               @      2@                      �?       @      1@      �?      �?       @      @      2@       @              @      @      :@      @      �?       @      @      ;@       @      �?              @      8@       @      �?      @      @      <@              �?              @      5@              �?      �?              9@      @              �?              9@      �?      �?       @              2@      @      �?              @      5@      @                              2@              �?      @      @      3@                      @      @      2@      @      �?      �?      �?      4@      �?      �?      @      @      5@      @      �?       @      @      3@      @      �?      �?      @      9@      �?              @              1@      @              �?              2@                       @              0@      �?      �?      �?       @      <@              �?              �?     �A@                      @              3@                      @              4@              �?              @      6@      @              @              2@              �?      �?      @      3@      �?      �?      @       @      1@      @      �?      �?      @      1@                       @      @      4@      @      �?               @      1@      @              �?      @      0@      @      �?       @      @      2@                      �?       @      9@                      @       @      3@      �?      �?      @      @      2@      @      �?      �?      @      9@              �?      @      @      7@      @      �?      @              4@      �?      �?      �?      @      4@      @      �?                      ;@      �?              @      @      1@       @      �?      @      @      9@      �?              @              5@                       @              7@      �?              @              5@       @      �?      @      @      =@       @              @      @      :@      @              �?              2@      �?              @      �?      1@                              @      3@      @      �?      @      @      4@                      �?      @      :@      @                      �?      3@              �?      �?      @     �@@       @      �?      @      @      1@      @      �?      �?              4@              �?              @      7@              �?      �?      @      <@      @      �?      �?              8@                       @              2@       @      �?      @      �?      7@      @              �?      @      ;@      @      �?      �?      @      8@      @      �?      �?      @      8@       @              @              3@                      �?      @      9@       @              @      @      9@              �?       @      @      7@      �?      �?      @              2@      �?              @      @      2@       @              @      @      6@      @      �?      @      @      1@      @      �?      @              2@      @      �?       @      @      2@      @               @      @      @@                       @              8@       @      �?      @      @      6@              �?               @      4@      �?      �?      @              6@      @      �?      �?      @      8@              �?      �?              A@       @              @              1@       @      �?      @              1@       @      �?      @              2@                      @      @      0@      @      �?              @      1@              �?              @      :@                      @      @      0@              �?      @       @      >@       @              @      @      @@      @              @      �?      8@      @      �?      @      @      >@      �?      �?      @       @      2@      �?      �?      @      @      1@       @              �?      @      2@                                      :@      @      �?      �?      @      ;@      �?              @              4@       @              @      @      1@      �?               @      @      4@      @               @      @      8@       @              @      @      1@      �?              @      @      2@       @              @      @      6@      @      �?      �?      @      A@      @              @              7@      @      �?      @              0@       @      �?      @      @      3@      �?      �?      @      @      3@                      @              2@      @      �?               @      :@       @      �?       @              :@      �?              @      @      6@      @              �?      @      4@       @              @      @      :@      �?      �?      �?      @      3@      �?              @      @      3@      @      �?      @              4@      �?              �?      @      >@                       @      @      0@       @              @              6@      @      �?      @       @      7@      @               @       @      0@                      @      @      :@      @      �?      �?      @      7@      �?      �?      @              5@       @              @      @      2@      �?              @      @      4@       @      �?      @       @      5@       @      �?      @       @      2@      �?      �?      @       @      7@      �?              @      @      4@       @      �?      @      @      5@      �?      �?      @              1@      �?      �?      @              2@      @      �?                      8@      �?      �?      @      @      7@      @              @              2@      @      �?      �?      @      1@       @      �?      @       @      6@      �?      �?      @      @      5@       @      �?      @      @      9@      �?      �?      �?      @      7@              �?              @      3@       @              @              2@              �?      @      @      1@       @      �?               @      2@      @              �?              6@              �?      �?       @      <@      �?              @              0@       @              @      @      1@       @              @      @      8@      �?              @      @      0@      �?               @      @      8@      �?              @      @      1@       @              @              2@      �?              @              2@       @              @      �?      4@      @      �?       @      @      1@       @              �?      @      6@      �?               @              4@                      @      @      1@       @               @       @      ;@      @              �?      @      4@      �?              @      @      =@      �?              �?      @      4@      �?              @              5@      @              @      @      5@      @      �?       @      @      1@      �?              �?              3@      @               @      @      4@      �?              @      @      2@                      �?      @      4@       @      �?       @              3@      @      �?      �?      @      8@      @      �?      �?              9@      �?      �?      �?              =@       @      �?      @              1@       @              @      @      6@      �?              �?      @      7@      �?               @              1@                      @      @      7@      �?      �?              @      4@       @      �?      @      @      2@      @      �?      �?      �?      2@       @                              <@      @      �?      �?              9@      @      �?      �?              8@      @      �?       @              8@       @      �?      �?              3@      �?      �?      �?              @@              �?      @       @      1@      �?              @      @      0@      �?              @              9@                      @              2@      @              @              1@       @              @       @      3@                      @      @      5@      �?              @      @      6@      @      �?      �?      @     �B@       @              @              6@      �?              @      @      4@      @              @      @      2@              �?      �?              ;@       @      �?      @              2@      @      �?      �?              0@      �?              @      @      6@      @      �?      �?              6@      �?               @      @      2@              �?      @      @      6@      �?      �?      �?      @      2@      �?      �?              @      ;@              �?       @              4@      @               @       @      ?@       @      �?      @      @      4@      @              �?      @      1@                      �?              0@                       @      @      9@                      @      @      1@      �?      �?      @              1@                      @      @      7@                      @              6@              �?      �?       @      5@       @              @      @      8@              �?      @      �?      5@              �?      @      @      <@              �?      �?       @      1@      �?              @      @      6@      �?              @       @      8@              �?      �?      @      4@      @              @      @      6@      �?      �?      �?      @      1@                      @              6@      @      �?      �?      @      :@      @      �?      �?      �?      8@       @      �?      �?      �?      5@      @               @              7@      @      �?              @      3@       @              @              8@      @              @       @      1@      �?      �?       @      @      6@      �?      �?       @              3@      �?      �?              �?      4@              �?      �?      @      2@      @      �?              @      3@      @              @      @      3@      @               @              ?@      @              @              6@      @      �?       @              6@              �?       @       @      4@      @      �?      �?      �?      7@      @      �?      �?      �?      B@                      @      @      7@                      @              7@       @      �?       @              5@      �?              @       @      1@                      @              7@       @               @              1@      @              �?      "@      3@      �?              @      �?      5@      �?               @              4@       @      �?      @              4@              �?      @      @      4@      �?              �?      @      :@      @      �?      @      @      3@      �?      �?      �?              5@      �?               @      @      7@       @      �?      @       @      1@      �?      �?       @              2@                      @      @      7@      �?              @      @      9@      �?      �?      @              5@      �?      �?      @              A@      �?              @              1@      �?      �?      @      @      1@              �?      �?       @      3@              �?       @      @      0@      @      �?      @      @      8@      �?      �?       @      �?      7@       @      �?                      4@              �?      @       @      4@                      @              5@              �?              @      6@      �?              @              6@      �?              @       @      =@      �?      �?       @              9@      �?               @      @      6@       @              @      @      3@                      @      �?      8@      @              @      @      9@       @              @      @      8@              �?      �?      @      6@      �?      �?      @      @      1@      �?      �?      @              0@      �?              @       @      8@                      �?              5@      �?              @      @      3@      @      �?                      6@       @              @              1@      �?      �?       @      @      <@      @              �?              8@      @      �?       @      @      0@       @      �?      @      �?      4@      �?      �?       @              7@      @      �?      @              1@       @              @              0@                      @      @      2@              �?                      5@      �?              @              >@      @              �?      @      1@      @      �?               @      3@       @              @              0@      �?      �?      @              6@      @      �?       @      @      1@       @      �?      @       @      :@       @      �?      �?      @      >@                      �?      @      <@      @              �?      @      6@                      �?              4@      @              @              6@       @      �?      @       @      8@       @      �?      �?      @      6@      @              �?      �?      =@      �?      �?       @       @      9@      @              �?              3@      �?               @      @      9@              �?              @      7@      @              �?              6@              �?      @              4@      �?      �?      �?      @      8@              �?       @              4@       @              @              =@      �?      �?      @              5@      �?      �?      @      "@      4@       @      �?      @      @      4@                      @       @      4@                      @      @      1@      @      �?      @      @      1@      @      �?      �?              7@      @      �?      �?      @      7@      @      �?      �?              4@              �?      �?              0@                      @      @      1@      @              @              2@              �?              @      1@       @      �?      �?      @      7@      �?               @      @     �A@      @      �?      @       @      3@       @      �?      @      @      1@      @      �?      �?              6@      �?              @      @      1@                              @      3@      �?               @      @      :@       @              @       @      7@              �?       @      @      4@                      �?      @      5@      �?      �?      @      @      1@              �?      �?      @      4@      �?      �?              �?      5@      �?              @              3@      �?              @      "@      5@                       @              9@       @      �?      @              2@      @      �?      @              6@      �?      �?      @      @      4@      �?              @              8@      �?              @              0@              �?      @      @      5@      �?      �?      @              >@      @      �?       @       @      7@      �?      �?      @       @      :@      @              �?      @      8@                      @      �?      0@                       @              3@      @      �?      �?      �?      ;@      @              @              2@      �?      �?      �?      @      3@      @      �?      @      @      4@      @      �?              @      @@      �?              @              2@                      @      @      4@              �?      @      @      1@      �?               @       @      0@      @                              :@      �?      �?      @              0@      �?              �?              4@                      @      @      2@              �?      @              2@      �?               @              2@      @      �?      �?      �?      8@              �?      @              <@      �?               @              7@                      @       @      1@      �?      �?                      :@      @      �?      @      @      3@      @                              0@      @      �?      �?      @      ;@              �?               @      6@       @      �?      @      @      3@       @      �?      @      @      0@              �?      @       @      3@                      �?      @      ;@      @      �?      �?      �?      <@       @      �?      @      @      8@              �?      @              1@       @              @              0@      @              �?      @      5@      @              @      @      6@                      �?      @      4@                      @      @      6@      �?              @              5@       @              @      @      0@       @      �?      @      @      8@      @      �?      �?              1@      �?              @              6@       @              @              :@              �?              @      =@       @              @              4@      �?      �?       @      @      4@              �?       @      @      >@      �?              @              1@              �?       @      @      ;@      �?              �?      @      7@       @              @              9@      @      �?               @      0@              �?      �?      @      :@      �?              �?              2@       @      �?      @       @      1@       @              �?              3@      @      �?      @      @      :@                      �?      @      ;@      �?              @              7@      �?      �?       @      @      1@      �?              @              8@      @              �?              6@       @      �?       @      @      3@      �?              @              7@      �?      �?              @      4@      �?      �?      �?      �?      1@              �?      @              <@      @              @              1@       @      �?       @      @      7@              �?       @      @      1@      �?      �?      @      @      B@              �?              @      5@                      �?      @      4@                      @              5@      �?      �?      @       @      2@              �?      �?      @      4@              �?      �?      @      3@      �?      �?      @              3@      �?      �?      @      @      6@      @      �?              @      8@      @      �?      �?      @      <@      �?              @      @      6@                      @              4@      @      �?      @      @      8@      �?              @      @      >@              �?      �?       @      8@      @              @      @      7@              �?      @      @      6@              �?      �?      @      8@      @      �?      �?       @      <@              �?      @       @      4@      @      �?      @      @      5@      �?              �?              7@       @      �?      @      @      0@              �?       @      @      ;@       @              @              3@      �?      �?      @              4@       @              @      @      8@              �?               @      1@       @                       @      6@              �?              @      A@      �?      �?      �?      @      7@      @                       @      6@      @      �?       @              2@              �?      �?              1@      @      �?      �?      @      :@      �?      �?      @      @      ;@      �?              @              2@              �?      �?      @     �@@      @      �?      �?      @      7@      @              �?      @      4@              �?      �?      @      >@      �?      �?               @      =@                      @      @      1@      @      �?      �?      @      :@      �?      �?                      6@       @              @      @      4@                      @      @      2@       @      �?       @      @      9@      @              �?              1@      @      �?       @              1@      �?              @      @      3@       @              @              0@      �?      �?              @      9@       @      �?      �?              <@                                      1@      @      �?      @      @      5@                       @      @      0@      @      �?                      3@      @              @              6@      �?      �?      @              6@      �?              @              5@       @              @              5@      �?                      @      8@       @              @      @      8@      @      �?      �?              ;@      �?               @      @      >@              �?      @              1@                       @      @      2@      @      �?      �?      "@      7@      @      �?      @      @      6@      �?      �?              @      7@       @      �?      �?              4@       @              @      @      4@      �?      �?       @              5@      @      �?                      7@      @      �?      �?       @      5@      @      �?              @      8@       @      �?      @              0@              �?       @      @      :@              �?              �?      7@      @              �?      @      9@      �?      �?      @              1@      �?              �?              9@       @                              2@      @              �?              1@                      @      @      1@       @      �?      @      �?      7@       @              @       @      5@      �?      �?      �?              <@                      @              2@                       @              7@      @               @              2@       @      �?      @      @      3@      �?      �?                      8@      �?              @      @      5@      �?      �?              @      2@      �?              @       @      6@      �?               @              =@      �?      �?       @      @      3@              �?      @       @      9@       @      �?      �?       @      9@      @              @       @      3@       @      �?      @      @      7@                      @      @      4@      �?      �?      @              <@      @              �?      @      7@      @      �?      �?       @      3@      @      �?      �?      @      =@      @      �?      �?              2@                      @              2@      @      �?      �?      @      1@                      @      @      1@      �?      �?                      7@      �?      �?              @      4@       @      �?       @              2@      @      �?      �?      @      4@              �?      �?      @      :@      @      �?      �?      @      B@      �?      �?      @       @      7@       @              @      �?      4@                              @      5@      @              @       @      4@      @      �?      �?      @      6@      �?      �?      �?              5@      @      �?      �?      @      :@      @      �?              @      =@                       @      @      4@      @      �?      �?              9@      @      �?      �?      @      =@              �?      �?      @      5@      �?      �?       @      @      4@      @      �?      @      @      2@      �?      �?      @      @      3@      �?      �?      �?      @      3@      @               @      @      7@              �?              @      4@      @              �?      @      9@      @                      @      4@                      �?       @      6@                      @      @      7@      @      �?              @      =@      �?                              5@      �?              @      @      :@       @      �?      �?      @      @@              �?       @      @      6@              �?      �?       @      @@                      @              3@      @              �?      @      7@      @      �?                      4@      �?              �?      @      ?@      �?      �?      @              1@      �?               @              8@      @      �?      @      @      1@              �?       @       @      2@      �?               @      @      6@                       @              :@      �?      �?      @      @      5@      @      �?      @      @      9@      @              @      @      5@      �?      �?      @              4@                      @      @      1@                       @              5@      �?              �?              8@              �?              @      1@      �?              @       @      0@      �?      �?      @      @      1@              �?      �?      @     �A@                      @              0@       @      �?      @              4@              �?      @      @      4@              �?      �?      @      1@      �?      �?      @      @      A@              �?               @      :@      @                              8@       @              �?      @      7@      @              @      @      3@       @              @      @      4@      @      �?      �?              1@      �?                              1@                      @      @      3@      �?      �?      �?              <@      �?      �?      @      @      ;@      @      �?       @      @      ;@       @              @              0@      �?      �?      �?      @      9@              �?      �?      @      ?@      @              �?              8@      �?      �?      �?      @      4@      �?               @              2@      @              @      @      2@       @              @              2@       @      �?      �?      @      6@      �?              @      @      2@              �?      �?      @      0@      @      �?              @      =@      �?      �?      @      @      6@       @      �?      @              1@              �?       @      @      4@      �?      �?       @      �?      7@      �?              @      @      0@      @                      @      4@      �?      �?       @       @      2@      @      �?      �?      @      8@              �?      @      @      0@              �?      �?              5@                      @      @      2@              �?       @      @      1@      @              @              0@       @      �?      @              6@      �?      �?      @      @      6@              �?      @              0@                      �?      @      :@      �?              �?      @      <@      @      �?              @      :@      @               @              8@                      �?              7@       @              @      @      5@      @                      @      6@              �?      @      @      2@              �?       @              2@      �?              @       @      =@       @      �?      @      �?      8@      @      �?       @              8@              �?      �?      @      3@      @              @              3@      @              �?              4@      @               @              :@      @      �?      �?      @      6@                       @      @      :@              �?       @              1@      @              @              9@                      @      �?      2@       @      �?      @      �?      5@              �?       @      @      1@              �?      �?      @      3@              �?      @              1@       @              @      @      2@      �?              @              5@       @      �?      �?              2@       @      �?      �?      �?      9@       @      �?      @       @      3@                      @      @      7@      �?      �?      @      @      8@       @              @              =@      @      �?      �?              1@      @              �?      @     �A@      �?                              =@      @      �?      �?              8@      �?      �?      @      @      ;@              �?      @      �?      =@      �?      �?      @      @      4@       @              @              8@      @      �?      �?      @      ;@      @      �?      �?      �?      6@      �?              @      @      :@      @              �?       @      4@      �?      �?                      5@                              �?      6@       @      �?       @      @      5@      �?      �?      @      @      4@              �?      �?              2@      @              �?      @      1@              �?      �?              5@      @      �?      �?      @      >@      @              @              1@      @      �?      �?      @      4@              �?      �?       @      9@       @      �?      @      @      2@      @                      @      <@      �?              �?      @      <@                      @              3@      �?      �?       @      @      1@                      @              8@      �?      �?      �?       @      4@      @      �?      @      @      1@       @      �?       @       @      4@      @                              2@      @      �?      �?      @      4@                      �?      @      7@      �?              �?      @      0@              �?                      5@      �?              @              8@       @              @              9@      �?      �?       @       @      :@              �?      �?              <@                      @      @      3@      @      �?      @      @      7@      @      �?      �?      @      9@      @               @              1@       @      �?      @       @      0@      @      �?      �?      @      @@      @      �?      �?      @      5@      @              @      @      >@      @              �?              9@              �?      �?      @      8@      �?              @      @      8@      @      �?      �?              6@                       @       @      8@      �?      �?       @      @      8@       @              �?      @      1@              �?      @      @      8@       @              @      @      :@      �?      �?      @              1@      �?      �?      @      @      0@                      �?              3@      �?      �?      @              8@              �?                      1@              �?              @      4@      @      �?       @      @      ;@       @              @      @      9@                      @      �?      3@       @      �?              @     �@@                      @              0@                      @      @      7@      @      �?      @      @      6@              �?      �?              2@      �?      �?      �?              7@       @      �?              @      2@       @      �?      @              6@      �?      �?      @      @      1@              �?      @      @      2@      �?               @      @      6@      @      �?      �?      @      8@              �?      �?      @      @@      @               @      @      1@      @      �?      �?              6@      @              @      @      3@                       @      @      9@       @               @              7@       @      �?      @              7@      �?              �?      @      3@      @      �?      �?              :@      @      �?      �?      @      6@      �?      �?      @      @      9@      �?              �?              :@      @      �?      �?      @      8@      @              @      @      3@      �?      �?      �?       @      3@       @      �?      @      @      8@      @      �?      �?      @      ;@       @      �?      �?              @@      @      �?      �?              6@      @      �?      �?      @      3@       @      �?      �?              7@      �?              @              3@      @      �?      @      @      1@      @      �?      �?       @      5@      �?      �?                      2@       @              @      @      0@      �?                      @      2@                      �?       @      8@      �?      �?       @              4@              �?      �?      @      5@              �?      �?       @      8@      @                              4@      @              �?      @      1@      �?              �?      @      9@      @              @      @      1@      �?      �?      @      @      ?@                      �?      @      6@      �?              @              3@              �?      @       @      1@       @              @              ;@      �?              @              0@       @      �?                      <@              �?      @              2@      �?              �?       @      9@      @      �?      @              2@       @              @      @      6@      @               @      @      9@       @      �?      @       @      6@      @      �?      @      �?      <@      @      �?      �?      @      3@              �?       @      @      0@              �?      �?      @      A@      @      �?      �?              6@      �?              �?      @      3@      @      �?      �?             �@@       @      �?      @       @      6@       @      �?      @      �?      4@      @      �?      �?      @      6@      �?      �?      @      @      6@      @      �?       @              1@              �?      �?      @      ;@      �?      �?      �?      @     �B@              �?      �?      @      ?@       @              @      �?      :@      �?      �?                      3@                      @              2@      �?      �?      �?      @     �A@                      @      @      ?@       @      �?      @      @      7@      @      �?      �?      @      ?@              �?      �?       @      5@              �?      @      @      1@      �?              @              7@      �?              @      @      1@       @      �?      @              1@      �?              @      @      1@              �?       @      @      5@      @      �?      �?      @      7@      @      �?       @      @      5@      @      �?      �?      @      4@      �?              @      @      5@      @      �?               @      4@      �?              @      @      1@              �?      @      @      2@      �?      �?      @      @      7@      @      �?      �?      @      4@      @              �?              7@              �?      @      @      6@              �?       @      �?      1@                      @      @      0@      �?      �?      �?      @      4@      �?      �?      �?      @      <@      @      �?       @      �?      ;@      �?              @      @      ;@                              @      4@      �?              @      @      5@       @      �?      @      @      3@      @      �?      @              8@              �?      �?       @      <@       @              @              2@      �?              @              1@      @      �?      �?              :@       @      �?       @              ;@                      @       @      3@      �?              @      @      5@              �?       @      @      5@                                      >@      @              @              8@      �?               @      @      9@      �?      �?      @       @      :@              �?      �?      @      =@      @      �?      �?      @      0@              �?      �?      @      5@      �?      �?      �?              3@      �?      �?               @      7@      @              �?      @      1@      @              @              3@      @      �?              @      2@      �?      �?       @       @      1@      �?      �?      @      �?      9@      �?              �?      @      8@      �?      �?                      2@                      �?      @      1@              �?      �?              1@              �?                      2@       @      �?       @              >@      �?      �?      @              0@              �?      @       @      1@      �?      �?              @      4@      @      �?       @      @      4@       @              @              2@              �?      @      @      1@       @      �?      @      @      7@              �?      �?              8@      �?      �?      �?       @      5@       @      �?      �?      @      7@                      �?       @      8@              �?      @      @      7@       @      �?      @      �?      1@      @              �?      @      7@       @      �?      @              6@      @              �?      @      1@      @              �?              5@      �?              �?              9@                                      5@      @      �?              @      3@      �?                       @      5@              �?      �?      @      0@      �?      �?      �?      @      6@              �?               @      4@       @               @              9@              �?      @      @      3@       @      �?      @      @      ;@      �?              @       @      2@      @      �?                      1@       @      �?      @              2@      �?      �?              @      6@              �?      �?              9@       @               @              5@      �?              @      @      0@              �?              @      1@      @               @      �?      3@      @              �?      @      7@      �?                              2@      @      �?      �?      @      :@      @      �?                      5@      �?              �?      @      <@      �?              @      @      5@                      @              3@                      @      @      6@      �?              �?              5@              �?      �?              3@       @              @             �A@      �?              @      @      7@      �?      �?      @              1@      @      �?       @      @      7@                      @      @      7@      @      �?              @      4@      @              @              2@      �?      �?      @              7@      @      �?      �?              7@                       @              3@      @                      @      4@                      �?      @      5@      �?               @      @      :@      @                              2@      �?              @      @      9@                              @      8@       @      �?       @      @      9@       @      �?      �?      @      4@      �?                              ?@              �?      �?      @      :@       @                      @      3@              �?       @              4@       @      �?      @      @      6@      �?              @              5@                       @      @      3@              �?      �?      @      @@      �?      �?       @              <@      �?      �?      @      @      1@                      @              1@              �?      @              8@              �?              @      :@              �?                      4@                      @              1@      @              @      @      0@      �?              @       @      7@       @      �?      �?      @      5@       @              @      @      >@              �?      @      @      0@                      @       @      1@      �?              �?       @      <@      �?      �?      @      �?      3@      @              �?              8@      @              @      @      6@       @      �?              @      7@      �?      �?      @      @      6@                      @      @      2@              �?      �?      @      2@      �?      �?      �?             �@@              �?      �?      @      8@      @      �?      �?      @      3@      @      �?              @      4@                      @              7@      �?      �?      �?      @      :@      �?              @              3@      �?              �?      @      8@                      @      @      2@      �?      �?      @              1@      @                      @      5@      �?              @      @      5@       @      �?                      3@      @      �?      �?      @      9@       @      �?      @      @      2@      @              @      @      5@      �?                              9@      �?      �?               @      <@                       @      @      9@      �?      �?      @      @      5@      @               @      @      4@      �?                              3@      @      �?      @      @      8@      @      �?              @      6@      �?              �?      �?      3@       @              @              4@      �?      �?       @       @      7@      �?      �?      �?      @      7@      �?      �?      �?      @      4@      @              �?      @      =@                      �?      @      <@      @      �?      �?      �?      9@      �?              @              5@      @      �?      �?       @      3@              �?                      3@      @              @      @      9@              �?      @              1@      �?      �?      �?      �?      1@      @      �?      �?              <@              �?                      6@      @      �?                      4@      �?              @              4@      @               @      @      6@       @              @      @      4@      @      �?      �?      @      6@      @               @              3@              �?      @       @      6@       @      �?      @      @      1@      �?      �?      @              2@      �?      �?              @      :@      �?      �?      �?       @      <@      �?              @      @      2@                      �?      @      2@      @                              1@      �?      �?                      7@      �?      �?       @      @      ;@                      �?      @      9@      �?              @              :@                       @              5@                      @              =@      @      �?              @      1@      �?      �?       @      @      5@              �?      @      @      2@              �?      �?              ;@      @      �?      �?      @      9@      �?              @              2@       @      �?      @       @      2@      @               @      @      7@      @              �?      @      3@      �?               @       @      0@      @      �?              @      :@       @              @              5@       @              �?      @      =@       @              @      @      >@      �?              �?      @      2@                      �?              1@      @      �?      �?      �?      @@      @      �?      �?      @      :@       @      �?      @              4@      @               @      @      1@              �?      �?              1@      �?      �?      @              4@                                      4@      �?              @      @      1@      @      �?      �?      @      7@      @               @      @      1@       @      �?      @       @      1@              �?       @      @      B@      @      �?       @      @      2@      @      �?      �?      @     �@@      �?      �?       @      @      3@              �?      @       @      8@      �?              @       @      2@              �?      �?      @      ?@      �?      �?      @      @      6@       @      �?      @      @      6@       @              @      @      4@      �?      �?      @              5@      @              �?      @      8@      �?      �?      @              3@              �?      @              3@                              @      8@                      �?      @      8@                      @      @      3@                              @      5@       @              @      @      2@              �?       @      @      4@              �?      �?              A@      @              @      @      1@      @      �?                      1@       @      �?      @      @      9@                      @              8@                       @       @      9@      @      �?      �?              9@              �?      @      @      3@      �?                              0@      @               @              5@      @      �?      �?              8@              �?      @      @      ;@       @              @              ;@              �?      �?      @      9@      @      �?      @              0@       @              @              5@                       @       @      2@      �?      �?      �?      @      6@                      �?      @      :@      �?      �?      �?              5@      @              �?      @      2@       @              @      @      1@       @              @      @      0@      @              �?      "@      B@      �?      �?              @      7@       @      �?      @      @      >@              �?       @              1@      @              �?              1@                      @      @      2@      �?      �?      @       @      @@      �?      �?      @              2@                      @              1@      �?                      @      7@      �?               @       @      :@      @              @      @      8@      @              @              9@      �?              �?              6@      �?               @      @      4@      @      �?      �?       @      <@                      @      @      5@                      �?              8@      @               @              7@      �?      �?      @      �?      5@       @              @              ;@      �?      �?      @      �?      <@                      @       @      1@      �?      �?      @      @      3@       @      �?      @      @      >@      �?              @      @      :@       @               @      @      1@      @                      @      7@              �?              @      6@      @                              2@       @                      @      5@      �?               @      @      3@              �?       @      @      :@      �?      �?      @      "@      4@       @              �?              3@      �?              �?              9@              �?      @      @      6@      �?      �?      @       @      2@      @      �?      @      @      0@                       @              3@                      @      @      1@                      @      @      1@       @      �?      @      @      <@      �?      �?      @      @      7@      @      �?      @              6@                       @              <@      @              �?      @      4@       @      �?       @      @      4@      �?      �?      �?      @      6@       @              @              0@      @      �?      �?      @      9@      �?              �?      �?      :@      @      �?      @              1@                      �?      @      <@      @      �?              @      8@                      �?      �?      5@                      �?      @      <@      @              �?       @      4@       @              @      @      9@              �?      �?              7@                      �?              0@                      @              7@      �?      �?      @      @      2@              �?       @      @      :@      @              �?      �?      @@      �?              �?      @      =@                      �?              6@                      �?      @      5@                      @      @      9@      @              �?       @     �@@      �?      �?      @              6@       @      �?              @      1@      �?              @       @      9@              �?       @       @      4@      @      �?      �?      @     �A@      �?              �?       @      ;@      �?      �?      @      @      7@      �?               @      @      6@      �?      �?      @       @      8@              �?       @      @      ?@              �?                      1@              �?      @      @      ;@      @              �?              7@       @      �?              @      2@      �?      �?       @       @      B@      @               @      @      2@      �?      �?      @      @      1@       @                              :@                      @              3@      @              @              ;@       @      �?      @              4@              �?      �?      �?      3@              �?      @      �?      4@      @              �?              6@                       @      @      6@      @              �?              2@      �?      �?      �?      @      :@       @      �?      @              0@      @               @      @      7@      @      �?      �?              :@      @      �?      @      @      9@                       @              3@      @              �?      @      6@                      @              9@       @      �?              @      <@       @      �?      @              8@      @      �?      �?      @      ;@       @      �?      @              1@                      @              0@      @      �?      @              3@      �?              @              7@      �?              @              4@      �?              @       @      2@      �?      �?      �?       @      4@       @              @              7@       @      �?      @              4@      @              @              4@       @      �?      @      @      0@      �?      �?      @              0@      @      �?      @              5@      �?              @      @      1@      �?              @      @      2@      �?              @              1@      �?      �?              @      4@      @              �?      @      3@                      @              5@      �?      �?                      7@      �?              @      @      :@       @      �?      @      @      5@              �?      @      @      4@       @              @      @      7@                       @      @      0@      @      �?       @              6@      �?      �?       @      @      2@      @      �?      �?      �?     �@@       @      �?      @      @      2@              �?      @      @      1@      �?              @      @      6@      @      �?      �?              3@      �?      �?      @      @      1@      �?              @              0@       @      �?      @              8@                      @      @      8@              �?               @      4@      @              @       @      2@      @               @              3@      �?                      @      5@      @      �?              �?      7@      �?              @              2@       @      �?      @      @      0@      �?                      @      1@      �?      �?                      8@       @              �?       @      9@              �?      �?      @      3@      �?              �?      @      5@       @              @      @     �@@       @      �?      @      @      5@      @      �?      �?      @      3@              �?      �?      @      <@      �?                              =@      @      �?              @      2@      @      �?       @      @      1@      @              @      @      @@       @      �?      @       @      4@              �?       @      @      5@                      @              3@      �?      �?      �?      @      5@      @                      @      6@              �?      �?      �?      1@      @      �?      �?              5@      �?      �?      �?      �?      4@                      �?      @      B@                      �?      @      8@      �?      �?      �?              ?@      @              �?       @      3@              �?      @      @      4@       @              @              1@                              @      ;@                              @      4@                      �?       @     �A@      �?      �?      �?      @      ;@      @              @       @      2@      @      �?      @       @      1@      @      �?      �?       @      7@       @              @      @      3@      @                      �?      3@      �?               @      @      2@      @      �?      �?      @      5@      @      �?      �?              1@      @      �?      �?      �?      @@       @      �?       @       @      4@      @              @      @      7@       @      �?       @      @      5@      @      �?      @      @      4@      �?      �?      �?              9@       @      �?      �?      �?      8@      �?      �?       @       @     �@@      �?                              <@              �?      @      @      3@      �?      �?                      4@      @      �?              �?      6@       @      �?      @      @      3@      �?      �?              �?      :@                      @      @      8@      �?      �?      @      @      4@       @              @              2@      @              @      @      2@      @      �?      �?      @      @@      �?      �?      @       @      >@      �?              @      @      4@      �?              @              0@                       @      @      0@      @      �?       @      @      1@       @              @      @      9@      @      �?       @      �?      A@      @              �?      @      5@       @      �?      @      @      6@      @      �?      �?      @     �@@              �?                      2@              �?               @      2@      �?      �?       @      @      4@              �?      @       @      6@       @              @              3@      @      �?                      4@      @      �?      �?       @      9@      �?      �?                      =@      �?      �?      �?       @     �A@       @              @              >@              �?      �?      @      2@              �?      @              0@      �?      �?               @      <@              �?      �?      �?      6@      @      �?      @              1@                      @      @      7@      @               @      @      7@                      @              2@              �?      �?              :@      @                      @      4@       @      �?      @      @      0@      @      �?              @     �@@                      @      @      2@      �?      �?      @      @      1@       @      �?      @      �?      1@       @      �?       @      @      2@      �?              @       @      3@      @      �?      �?       @      8@       @              @      @      >@              �?      @       @      2@       @      �?      �?      @      ?@              �?      @      @      6@       @               @      @      1@      @      �?       @       @      2@      �?              @              1@      �?               @      @      2@      �?      �?      �?      @     �@@       @      �?               @      7@       @      �?      @      �?      5@      �?      �?      @      @      4@                              @      7@      @      �?      @              7@      @              �?      @      B@                      �?              7@      @      �?       @      @      3@      �?              @              2@       @      �?      @      @      >@                      @      @      8@       @              @              3@       @      �?      @      @      >@       @      �?      @              0@      @      �?      �?      @      >@      �?      �?      @      @      5@      �?      �?      @      @      1@      @                              3@      @      �?      �?              1@      @      �?       @              4@                       @      @      4@      @      �?               @      3@      �?      �?      @       @      1@      �?               @              5@      @      �?      @      @      1@                      @      @      3@      �?      �?      @              3@      �?              @              7@       @      �?      @      @      7@      @      �?      �?              2@                      @      @      7@      �?              @              5@      @      �?      �?      @      5@      @              @              2@              �?      @       @      4@      @      �?      @      @      1@                      �?              4@              �?       @              =@                      @      @      7@       @      �?      @              4@                      �?             �@@      @      �?      �?       @      6@      @      �?      @              2@                       @      @      7@       @              @              9@              �?      @      @      8@      �?              @              5@                      @              ;@      �?      �?      @              0@      �?      �?              @      4@      �?                      �?      :@      @      �?       @      @      9@      @      �?                      5@              �?      @              2@       @      �?      @      @      4@      @              �?              1@       @                              7@      @      �?      @              2@              �?              @      1@                       @      @      2@      @      �?      �?       @      8@      @      �?       @              6@                       @      @      A@                      @      @      5@      @      �?       @       @      1@      �?                       @      0@                      @              5@      @      �?              @      2@       @              �?              3@      @      �?      �?      @      :@              �?      @      @      :@      @               @      @      <@      �?      �?       @              3@      @      �?                      5@      �?      �?      @      @      6@                      �?              ?@              �?      @              2@      �?                      @      5@      �?      �?      @      @      ;@      �?      �?      @      @      1@                       @              7@                      @      @      5@      @              @              :@      �?      �?              @      4@                              @      4@      @      �?      �?      @      3@              �?      @      @      6@      �?      �?      @      @      4@                      @      @      6@      �?              �?      @      2@      �?              @       @      1@                       @              =@      @      �?      �?      @      0@      �?      �?      @      @      1@      �?              @              0@      �?      �?      �?      @      1@              �?       @              9@                      �?              4@      �?              @      @      1@       @      �?       @      �?      0@      �?      �?      @      @      4@                       @       @      8@                       @      @     �@@      @               @      @      1@      �?      �?      @       @      8@              �?      �?              <@       @              @      @      <@                      @              4@      @               @              2@                              @      :@              �?              @      7@      @      �?      @       @      8@              �?      �?      @      ;@       @              @      @      9@      �?               @              5@      @      �?      @       @      6@              �?      @      @      7@      @              @      @      5@      @      �?      �?              4@      �?      �?       @      @      7@              �?       @       @      7@      �?      �?       @      �?      B@      �?      �?      �?      @      7@      @                      @      3@      @              �?              @@      �?                       @      ?@      @      �?       @      @      2@      @              �?              0@              �?              @      3@      �?              @              0@              �?      @       @      2@       @      �?      @              1@       @      �?      @      @      5@      @              @              4@              �?              @      2@      @      �?              @      =@       @      �?      @      @      A@      �?              �?      @      @@      @      �?      @      �?      2@      @              @      @      :@       @              @              6@      @              @      @      6@              �?      @      @      6@       @              @      @      ?@      �?              @              2@      �?              @      @      4@              �?       @              4@      @              �?      @      1@                      @              2@                      @      @      6@      �?      �?       @       @      0@      @      �?      �?              9@      �?      �?      @              8@      �?                              3@      @      �?       @      @      :@      @      �?       @      @      2@       @      �?      �?      @      5@              �?      �?              4@                      @              7@      @      �?              @      ;@      @      �?      @      @      3@       @              @              5@      �?      �?              �?      @@       @              �?      @      :@      �?      �?      �?              8@      @      �?      �?              1@       @      �?      @      @      1@                      @      @      1@              �?      @      @      9@      @      �?               @      6@      �?              @      @      5@       @      �?              @      2@                              @      <@      �?               @      @      4@      @              �?      @      2@                      �?      @      1@      @              @      @      5@      @      �?      �?       @      4@      @      �?      �?       @      6@      @                              5@              �?      �?      @      ?@              �?      �?              3@       @              @      @      8@      �?               @              8@       @              @              3@      �?      �?              �?      >@      �?      �?      �?      �?      3@              �?      �?      @      >@      �?              @      @      @@              �?                      4@                      @              1@                      �?      @      4@              �?                      @@                                      7@              �?      @              9@      �?      �?      @      @      :@                      @      @      2@      @      �?      �?      @      ;@       @              @      @      6@              �?      �?      @      2@      �?              @      @      5@      �?      �?      �?      @      9@                       @      @      5@      @              �?      @      7@              �?              @      3@      @               @      @      8@      �?      �?      @       @      1@       @      �?      @      @      4@       @      �?      @       @      2@                                      7@       @                      �?      0@      @              �?       @      6@                       @              4@      �?              @      @      2@      @      �?      @      @      5@      �?               @              1@       @              @      @      1@       @              @              7@      �?              @              0@                                      1@      �?              �?              ?@       @              @      @      4@      �?              @      @      ;@                      �?      @      7@      �?      �?              �?      6@                      @      @      4@      �?      �?      @              2@              �?      @       @      1@       @      �?      @      @      ?@      �?              @      @      4@      �?              @              5@      �?              @      @      0@       @              @      @      2@       @      �?       @      @      7@      @      �?      @      @      1@      �?              @      @      1@              �?      �?      @      2@      @              �?      @      ;@       @      �?      @              2@      �?      �?      @      @      0@      @               @              8@                      @      @      :@              �?              @      <@                      @      @      3@                      �?              5@       @               @      @      8@       @                              5@       @              �?      @      1@      �?      �?      @              5@              �?                      0@      @      �?      @      �?      7@      �?              @              2@      �?              @      @      3@       @              @      @      4@      @              �?              ?@      @      �?      �?      �?      6@      @      �?      �?              6@       @      �?              @      2@      @              @       @      4@      @      �?      �?             �@@              �?      �?      @      0@      @      �?              @      8@              �?              @      9@      @      �?      �?      @      @@      @      �?      @              0@      �?              @              1@                      @      @      1@      �?      �?      @      @      6@      @      �?       @      @      2@                       @              =@      @      �?      �?      @      8@                      @              0@      @      �?      @      �?      4@                      @              5@      @      �?       @              8@                      @      @      9@       @      �?      �?              :@      @      �?              @      <@              �?      �?      @      7@              �?      @              5@              �?      �?      @      :@      @      �?      @      @      1@      �?      �?      @       @      4@                              @      1@       @      �?      @      @      :@      �?                      @      0@      @      �?      �?              3@      �?                              4@      �?      �?              @      6@      �?      �?              @      5@      @      �?      �?      @      5@       @      �?      @      @      3@              �?      �?      @      =@              �?      �?              6@       @      �?       @      @      4@       @      �?      @       @      6@                       @              4@      @      �?      @              0@      @      �?      �?      @      6@      �?                      @      8@       @              @      @      8@      @      �?      @      @      :@       @                      @      :@      @      �?      �?      @      4@      �?      �?       @              3@       @      �?      @      @      7@      @      �?      �?              0@       @      �?      @      @      3@      @              @      @      3@                              @      8@              �?      @      @      2@      �?              @      @      1@      @      �?      �?      @      0@      �?      �?      @              7@      @      �?      �?      @      7@              �?      �?      @      2@              �?       @              9@      @              @              0@      �?      �?      @      @      1@      @      �?      �?      @      5@      @              �?      @      7@      �?      �?      @      @      2@       @                              1@      �?      �?       @      @      >@              �?      �?              3@      @      �?      �?              5@                      �?      "@      ;@      @              @      @      2@                      �?      @      6@      �?      �?      @              2@              �?      �?      @      :@                      @              ;@       @      �?      �?              <@      @               @      @      1@       @              @      @      8@              �?      �?              3@      @      �?      @              2@              �?      �?       @      9@       @      �?      �?      @      5@      �?      �?      @              2@      �?              �?       @      3@      �?      �?      @      @      7@      �?      �?       @      @      8@       @               @      @      2@                      �?       @      @@       @              @      @      6@      �?              @       @      3@                       @      @      8@      �?              @      @      9@      @              @      @      1@      @      �?      �?      @      5@              �?       @      @      7@      �?      �?      @      @      7@      @      �?      @      �?      2@      @              @              1@              �?      �?      @      2@      @      �?              @      ;@       @      �?      @      @      >@      �?      �?      �?      @      <@       @      �?      @              0@      �?              @      @      2@       @              �?      @     �A@      �?              @      @      2@              �?      �?      @      4@      @      �?      �?      @      2@                      �?              8@      �?               @      @      :@      �?              @      @      5@      �?      �?      �?      �?      6@      �?              �?      @      <@              �?      @      @      4@      @      �?      @      @      3@      �?              �?      @      2@                      �?      @      5@      @      �?      �?      @      :@              �?       @              4@      @                              9@                      @              2@              �?      @      @      3@       @              @      @      6@              �?      @      @      0@                                      6@       @      �?      @              0@       @              @              6@      @      �?      �?      @      :@      @      �?      �?      @      1@              �?      @              5@              �?       @      @      4@      �?                       @      >@       @              @      @      4@      �?              �?       @      A@      @              �?              2@      @              @      @      4@      �?      �?      @      @      3@                              @      ?@      �?              @      @      3@      �?              @              3@      �?      �?      @      �?      :@      �?              @              ;@      �?      �?      @      @      5@      @              @      @      0@      �?      �?                      @@                      @      @      4@                       @              4@              �?              @      3@      @               @      @      ;@       @      �?      @              4@              �?              @      3@      �?      �?      @      @      2@      �?              @      @      ;@      �?      �?      @      @      1@      @      �?       @      @      2@       @              @              1@      �?              @      @      :@      @      �?      @      @      4@              �?      @      @      8@      @      �?      @              3@       @      �?              @      @@      �?      �?      @              5@       @      �?      �?      @      9@      �?               @              0@      �?      �?      �?      @      7@       @                      @      9@      @              �?      @      B@      @              @      @      ;@      @      �?      @      @      4@       @      �?      @       @      1@      @      �?              @      5@              �?      �?       @      =@      @      �?      �?      @      :@      @      �?      �?       @      <@      @              �?      @      <@      @              �?              1@      �?              @              <@      �?              @       @      2@                      �?      @      9@      @      �?      @      @      ;@      @      �?      �?       @      4@       @              @      �?      4@       @              �?      @      =@              �?       @      @      1@      @              @      @      5@      �?      �?              �?      5@       @      �?               @      >@      @      �?              @      2@              �?      @              3@      @      �?      �?              1@              �?      �?              >@      �?              @              2@      �?      �?       @              8@      @      �?       @              1@                      �?      @      1@       @                      @      <@              �?      �?      @      9@      @              @       @      0@              �?      @              2@      �?              �?              5@       @      �?       @      @      =@      �?      �?       @              7@      �?              �?      @      6@              �?      �?      @      6@              �?                      6@      @              �?      @      7@      @      �?              @      1@      @      �?              @      :@      �?              �?      @      3@      @      �?              @      9@      �?              @      �?      5@       @      �?      @       @      2@      @      �?      �?      @      9@              �?       @      @      8@      �?              �?              =@              �?      �?      @      <@              �?      @      @      7@      @      �?      �?      @      1@      @      �?                      4@      @              @      @      5@      @      �?      �?              ;@       @              @              1@      �?              @      @      7@       @      �?      @      @      >@                      @      @      0@      @              @      @      3@                      @      @      1@      @      �?      �?              5@                              @      3@      �?      �?      �?       @      4@              �?      �?              <@              �?      �?      @      6@      �?      �?      �?      @      5@      @      �?      �?              2@      �?      �?              @      <@       @                      @      :@      �?              �?      @      7@       @      �?      @      @      2@                      @      @      9@              �?      �?      @      9@      �?              @      @      2@                       @              :@              �?      @      @      8@      @      �?      �?      @      ;@              �?      �?      @      1@      �?              �?              ;@              �?      @              4@              �?      �?              4@      @               @      @      7@      �?      �?               @      :@      �?              �?       @      @@              �?      �?      @      5@      �?      �?      @      @      0@      @      �?      �?      @      7@       @                      @      1@      �?              @      @      0@       @              @      @      4@       @              �?       @      7@       @               @              0@       @              @              5@      @      �?      �?      @      5@      �?              @      @      3@      @      �?              @      8@                      @      @      2@              �?      �?      @      ?@      �?      �?      @      �?      1@       @      �?              @      5@       @      �?       @      @      7@      @      �?               @      6@      �?              @              7@      @      �?       @              1@              �?       @      @      6@              �?      @      @      5@       @              @              3@       @      �?      @      @      7@      �?      �?              @      :@      �?      �?      �?              8@       @              @      @      >@      �?      �?      �?              7@              �?      �?      @      :@      �?      �?      @      @      6@      �?      �?      @      �?      5@                               @      ;@      �?      �?      �?      @      ?@              �?       @      @      3@      @                       @      6@       @              @              ;@      �?      �?      �?              6@      @      �?      �?       @      9@              �?      @      @      9@              �?      �?              0@      @      �?      @      @      1@              �?      @      �?      4@      @              �?       @      8@      �?      �?      @      @      4@      @              �?              ;@       @      �?       @              :@      �?      �?      �?      @      3@              �?      �?      @      8@      @              @      @      0@      @              �?      @      4@      �?      �?              �?      8@      @                      @      :@              �?      @      @      4@      �?      �?      �?              3@      @      �?      �?      @      3@      @                      @      1@       @      �?       @              ?@       @      �?              @      4@                      @              4@       @              @      @      1@       @      �?      @      @      6@       @      �?      @      @      7@      @      �?                      0@       @              @      @      1@      @      �?      �?       @      :@      @                      @      B@      �?              @              1@      �?              �?              =@                              @      8@       @      �?              @     �@@      �?      �?               @      4@      �?      �?      @       @      8@      �?      �?              @      6@                      @              2@      @              @      @      4@                       @      �?      2@       @      �?      @      @      >@      @      �?      @       @      1@      �?                              2@       @      �?       @       @      4@                       @              4@      @      �?              @      4@      @      �?      �?      @      1@      �?      �?      �?              0@      �?      �?                      6@       @      �?      �?      �?      :@      �?      �?      @      @      5@       @              @              8@       @              @      @      4@      @              @              8@       @      �?      @              ?@                       @      @      2@       @      �?       @              ;@      �?              @      @      6@      @              �?      @      2@      �?              @              1@      @              @      @      :@      �?               @              8@      @      �?      �?      �?      8@              �?                      7@       @      �?      @              3@      �?      �?      @      @      3@                      @      @      9@      �?              @              2@      @               @              4@       @      �?      @              0@       @      �?                      2@       @      �?              @      5@              �?       @      @      5@              �?      �?      @      A@      �?              �?              7@      @              �?      @      2@      �?      �?       @              3@              �?      @      @      2@                      @              7@       @      �?      @      @      8@                      @              0@      @      �?      �?       @      6@      �?      �?                      =@      @      �?      �?              7@       @              @              2@                      �?              3@      @                       @      9@      �?      �?      @       @      1@                       @      @      1@      �?      �?      �?      @      2@       @      �?      @      @      7@      �?      �?      �?      @      2@      @      �?       @      @      7@       @      �?      @      @      0@              �?      �?      @      7@      @      �?      @      @      3@                      @       @      @@       @                      @      4@      @      �?      @      @      3@       @      �?      @              2@       @               @      @      0@                      @      �?      6@      �?              �?             �A@      �?              @       @      2@      @                              :@      @               @      @      1@      �?               @      @      6@              �?       @              8@       @      �?       @              4@      �?      �?      @      @      >@      �?      �?              @      7@      �?      �?      @      @      5@      �?      �?      �?              :@      �?      �?      �?      @      ?@      �?      �?      @              1@      @              �?              6@      @      �?      �?              A@                               @      <@                       @              8@      @      �?              @      4@              �?      @       @      4@      �?      �?       @      @      2@       @              @              1@      �?              @              :@      @              �?      @      >@      �?      �?      @              3@                       @              4@              �?      @      @      1@      �?      �?       @              8@      @      �?      �?      @      7@      @              �?       @      2@      @      �?      �?      @      7@      �?      �?      �?      @      ;@      �?      �?      �?              ;@      @      �?      �?              7@      @      �?      �?      @      >@      �?                              8@              �?      @              5@      @              @              2@              �?      �?       @      6@      �?      �?      �?      @      9@      @              �?              ;@      @              �?              8@      �?      �?              @      8@      �?              �?              ;@              �?      �?              ;@      @              �?              4@      @              �?      @      0@              �?      �?       @      7@       @              @              1@      @      �?      @      @      7@      @              �?      @      ;@      @      �?       @      @      7@      �?      �?      �?      @      =@      �?      �?      @      @      <@      �?      �?      @      �?      4@                      �?      @      4@      �?              @      �?      8@       @      �?      @      @      8@                      �?      @      3@      �?              @      @      <@      �?      �?      �?             �A@      @              �?      @      5@              �?      @       @      1@              �?      �?      @      =@              �?      @      @      6@                      @      @      9@      �?      �?      @              2@                      @       @      5@              �?      �?              A@      @               @      @      9@              �?      @       @      3@      @      �?      @      @      5@      �?              �?              9@              �?      @      @      1@      �?      �?      �?              =@      �?      �?      @      @      7@      @      �?      �?      @      ;@      @      �?      �?              2@      @              �?       @      0@                                      0@      @                      @      4@       @              @              2@      �?      �?      �?      @      8@      �?              @              :@              �?              "@      :@       @              @              3@      �?              @      @      3@      @      �?      �?              :@      @               @              ?@              �?      �?       @      8@              �?      �?              5@      �?               @      @      1@                      �?      @      :@      �?      �?       @      @      4@                      @      @      8@      @      �?      �?              ;@      �?      �?      @      @      3@              �?      �?             �@@      @              �?      @      1@      �?      �?      @              6@      �?              @              2@              �?      �?      @      7@       @      �?      @      �?      9@      �?      �?      �?       @      6@       @              @              6@              �?              @      8@              �?      @      @      8@       @              @      @      7@      �?              @              5@      @      �?      �?              2@      �?      �?      @              5@       @      �?      @      @      4@      @              �?      �?      3@      @              �?              4@              �?       @      @      4@                      @      @      7@              �?      @      @      1@      @      �?      �?              9@              �?      �?              :@              �?      �?      @      5@      @      �?      �?              :@       @               @      @      5@      �?               @              8@                      @      @      2@      @                              ;@      @      �?       @              :@      �?               @      @      6@      @                              2@      �?      �?                      0@              �?      �?      @      6@      �?              @              8@      @      �?      �?      @      8@                      @      @      :@      @      �?      �?      @      3@       @              @      @      6@              �?       @      @      4@                      @              1@      �?              @       @      6@      �?              @       @      4@      @      �?               @      2@       @              @      @      6@      @      �?      @       @      :@      �?      �?       @              6@      @              �?              2@      �?              �?              7@      �?              @      @      B@                      @      @      7@              �?              @      2@       @      �?      �?       @      ?@                      @       @      8@       @              @      @      9@                      @      @      6@      @              @       @      7@      @      �?      �?      @      @@      @      �?       @      @      4@      @      �?      @              :@       @      �?      @              3@      �?              @              1@      �?      �?              @      2@      @      �?      @              2@      @      �?      �?       @      3@      @      �?      �?      @      1@      @      �?      �?      @      6@      @               @      @      6@              �?      @      @      @@       @      �?      @      @      9@      �?      �?      @      @     �@@      @                      @      9@      @      �?      @      @      1@                      �?      @     �@@                      @      @      4@       @      �?      @      @      8@      �?               @      @      4@      �?      �?      @              7@      �?      �?      �?      @      :@      @              �?      @      >@      �?      �?       @       @      4@      @              @      @      3@      �?      �?      �?              6@      @              @              0@                      @      @      1@      @      �?      �?              7@                      @      @      6@      @              �?              4@      @      �?       @      @      3@       @              @              4@                      @              1@      �?              @      @      8@       @              @       @      3@                       @       @      1@       @              @      @      2@                      @      @      =@      �?      �?      @      @      7@      @              �?      @      9@       @              @      @      4@       @      �?      @      @      9@      �?               @              1@      �?      �?       @      @      5@      �?              @              5@      �?      �?      @      @      <@              �?              @      3@              �?      @      �?      3@      �?                              6@       @      �?      @              1@      @      �?      �?      @      6@      �?      �?       @              3@       @              �?      @      8@      �?               @              =@      �?              @       @      :@      @      �?       @      @      <@       @      �?      @              4@      �?              @      @      3@       @      �?       @      @      3@      @      �?      @      @      =@       @               @      @      9@      �?      �?       @       @      4@                                      5@              �?      �?      @      5@      @              �?      @      ;@      �?      �?                      <@              �?      @      @      5@      �?      �?      @      @      ;@      @      �?      �?      @      9@      @               @      @      5@      �?      �?      @      @      =@                      @       @      7@      �?      �?      @      @      2@                      �?      @      8@      @      �?      �?      @      5@      @              @              :@                       @      @      A@      �?      �?      @              1@       @               @              2@              �?              @      4@                              @      5@              �?      �?      �?      :@      @      �?      @      @      2@       @               @      @      3@      @      �?      �?             �B@       @      �?      @              7@              �?      �?      @      @@      �?              @      @      =@      @              @              6@      @              @              ?@      �?              @              9@       @      �?      @       @      6@      @      �?      @      @      5@      @      �?      �?      @      ?@      �?              @              7@      �?      �?       @      @      1@      @      �?      @       @      1@       @      �?              �?      <@      �?              @              1@      @              �?      @      8@              �?                      3@      �?      �?       @       @      2@      �?                              6@              �?      �?      �?      5@      @      �?       @      @      1@      �?      �?              @      8@              �?                      6@      @               @      @      0@       @      �?      @              3@      @              @      @      8@      �?      �?      @              2@      @      �?      �?      @      8@      �?      �?       @      @      2@      �?              @              3@       @                      @      1@       @      �?      @      @      2@      @      �?              @      7@      �?      �?       @      @      4@       @      �?      @      @      3@                      �?      @      1@                       @      @     �@@       @      �?       @      @      4@       @      �?       @              2@              �?      �?      @      5@      �?      �?       @      @      2@      @      �?      @      @      3@                      @              2@      �?      �?      @      @      9@      @      �?       @      @      ;@                              @      5@      �?               @      @      7@      @      �?      �?      @      8@      �?              @      �?      4@       @              �?              8@      @      �?              @      ;@      �?      �?      �?      @      8@              �?      �?      @      :@       @      �?       @      @      >@              �?      �?              6@              �?      @              4@              �?              @      :@      @      �?      �?       @      9@      �?      �?      @      @      6@              �?      @              6@       @              @      @      =@      @      �?       @       @      9@                       @      @      :@      @              @      @      7@      @      �?      �?      @      2@      @      �?      �?              <@                      @      @      6@              �?       @              3@      @      �?      �?      �?     �B@      @      �?       @      @      3@      �?              @      @      2@      @                              7@      �?      �?       @              3@                      @       @      3@                                      3@      �?      �?      @       @      3@                      @      @      4@      @      �?      @              9@      �?      �?      @      @      7@      @      �?      @      @      2@      @              @              5@              �?       @      @      0@      @      �?               @      9@      @               @      @      7@      �?              @      @      ;@       @      �?       @      @      6@      �?              @       @      <@      @      �?       @              5@      �?               @      @      9@                      @      @      1@      �?      �?      @              1@              �?       @              6@                       @       @      6@      �?      �?      �?      �?      4@                      @      @      ;@      @              �?      @      5@      @               @      @      4@                      @      @      A@       @      �?      @              0@      �?      �?      @      @      3@              �?      �?      @      <@      �?              @      @      1@                      �?      @      7@              �?       @              2@      �?               @       @      4@       @      �?      @       @      9@      �?      �?      @      @      1@      @      �?      @      @      0@       @      �?      @      @      4@       @               @      @      4@      �?              @              2@      �?               @       @      >@      @      �?              @      :@       @              @              4@              �?      �?              3@      @      �?      �?      @      <@      @               @      @      7@              �?      @      @      6@      �?      �?              @      :@      @                      @      :@       @              @       @      5@      @      �?      �?       @      5@      �?              @      @      1@              �?      @      @      2@              �?      �?      @      2@      @      �?      �?       @      8@      @               @      @      6@      �?              @      @      2@              �?      @      @      6@                      �?      @      9@       @      �?       @      @     �@@      @      �?      �?      @     �@@      �?              �?      @     �@@      @              �?      @      2@              �?      @      @      4@      �?      �?      @      @      9@              �?      @      @      5@      �?      �?      @              0@      @      �?      �?              =@                                      1@      @              @              5@      �?      �?      @      @      3@                                      4@      �?      �?      @              9@      @      �?      �?              ;@      �?      �?       @              2@      �?      �?      @              2@                      �?              4@                      @      @      8@              �?      @      @      1@       @      �?      @       @      7@      @              @      �?      2@       @      �?       @      @      5@      �?      �?       @      @      1@      @      �?      �?      @      @@              �?      �?              5@      @                       @      5@                      @      @      1@      �?      �?      @      @      5@      @              @              =@              �?              @      :@                      �?      @      4@      @              �?      @      2@      @      �?              @      :@      @                              4@      �?      �?      �?              2@      @              @              0@      @               @              :@      @      �?      �?              1@              �?      �?      @      1@      �?              @              3@              �?                      5@      �?      �?              @      5@                      �?      @      A@                      @      @      1@              �?      @      @      5@       @              @      @      1@              �?      @      @      2@              �?       @      @      ;@      �?      �?      @      �?      8@              �?               @      4@      �?      �?      @       @      :@                      @      @      7@      @      �?      �?              3@              �?      @      @      2@      @              �?      @      8@      �?              @              1@      @                              2@       @              @              1@      �?              @      @      5@      @              �?              3@              �?      @              1@       @              @              5@              �?      �?              8@              �?              @      ;@              �?       @      @      7@      �?      �?       @              4@                      @      �?      2@      @      �?              @      <@      @              �?      @      5@       @      �?      @              5@      @      �?      @       @      1@      �?               @      @      6@              �?      �?      @      5@      �?      �?      �?      @      :@      @               @              1@       @      �?      @      �?      6@       @              �?              2@      �?      �?      �?      @      =@      @              �?      @      :@              �?      @              8@      @      �?                      6@      �?      �?      @      @      1@      @               @      @      2@                      �?      @      2@      @      �?      �?              :@      �?              �?      @      9@      @      �?      �?      @      3@       @              @      @      0@                              @      5@      @              @      @      7@       @              @              5@      �?      �?              @      9@                       @              8@              �?      @       @      =@      �?              @              5@              �?      @       @      :@      @              �?              =@                      @      @      1@      @      �?      �?      @      >@      �?      �?      @              0@      �?      �?       @              =@      @              �?      @      3@      �?      �?      �?      @      ;@                       @       @      9@      @      �?      �?      @      2@       @               @              =@       @              @              4@              �?      �?      @      3@      �?              @      @      5@      �?              @      @      5@      �?              @      @      1@              �?       @      @      0@      �?                       @      <@      �?      �?              @      6@      @              @              6@      @      �?      �?      �?      =@       @              @      @      2@       @               @              ;@                      @              4@      �?      �?                      6@      �?              @      @      5@      �?      �?      �?      @      4@      @      �?      �?              5@      @              @      @      2@       @              @              5@       @               @      @      8@                      @       @      1@              �?      �?      @      1@              �?              @      1@                                      1@       @                      @      8@                      @       @      6@       @      �?       @              8@      �?      �?      @              4@      �?              @      @      2@      @      �?                      6@              �?      �?      @      9@      @      �?      �?      �?      @@      �?               @      @      6@       @      �?      �?              <@      �?      �?      @      @      4@                      @      @      2@                                      5@      @              �?      @     �@@                      �?      @      >@      @      �?      �?      �?      1@      @      �?      �?      @      8@      @               @              =@       @      �?      @      @      1@              �?       @      @      3@      �?              @      @      2@      @               @              1@                      �?      @      8@       @              @       @      4@      @      �?      @      @      0@       @              @              2@      @              @              5@      �?              @      @      8@      @                       @      2@              �?      @              1@      �?              �?      @      5@      @      �?      �?              3@      @               @              2@       @      �?              @      ;@              �?       @              1@      @      �?              @      2@       @      �?      @      @      8@      �?      �?              @      3@      �?                      @      2@      @      �?      �?      @      8@              �?      @              7@      �?      �?      @              5@              �?      @      @      7@      �?      �?              @      3@              �?      �?              :@                      @              5@                              �?      <@      @      �?      �?      @      6@      �?      �?      �?      �?      ;@      @      �?      �?      @      6@      �?                             �@@      @      �?      �?      @      2@                      �?      �?      :@      @      �?      �?      @      ;@      �?      �?                      7@              �?              @      >@       @              @      @      <@      �?      �?       @              7@      �?      �?      @      @      2@              �?       @      @      9@      �?              �?              ?@       @              @      �?      1@      �?      �?      @              4@      @      �?      �?              1@      @              �?      @      5@      @      �?      �?      @      8@                      @      @      3@       @      �?      @      @      5@              �?      @      @      4@      �?      �?      @              3@      �?              @              4@      @                      @      5@              �?      �?      @      7@      �?      �?               @      :@      @              @              2@      �?      �?      @      @      5@      �?              @              1@      �?      �?      @      @      0@      �?      �?       @              3@      @      �?      �?      @      0@      @              @      @      8@      �?               @              4@       @      �?                      8@      �?               @      �?      A@      �?      �?       @              4@                      �?              0@       @              @       @      2@      �?      �?      @       @      1@       @               @       @      =@      @      �?       @              7@      @      �?       @              3@       @      �?      @              4@      �?      �?       @      @      3@      �?                              0@                      @      @      8@      �?      �?      @      @      5@       @      �?      @      �?      8@              �?      �?      @      1@       @      �?       @       @      4@                      �?       @      <@      �?                      @      3@      �?      �?      @       @      4@      @      �?      �?      @      1@       @              @      @      3@      @      �?      �?              9@      �?                              1@      @      �?      �?      @      9@              �?       @      @      4@                      @      @      :@              �?       @      @      4@      @      �?      @      @      0@      �?      �?      @      @      2@      �?              @      @      4@                      �?      @      1@      @      �?      @      @      1@      �?      �?       @      @      <@      @      �?      �?              3@      �?      �?      �?      @      3@       @      �?      @              3@      @              �?              3@              �?      �?      @      6@      �?      �?      �?              ;@      �?              @              3@      @      �?      �?      @      6@      @      �?      @      @      5@       @      �?      �?      @      2@       @              @      @      6@      �?      �?      @      @      6@              �?      @              ;@              �?      @              7@       @              @      @      1@      @      �?      �?      @      8@              �?      @              2@      �?              @              2@       @      �?      @      @      9@                       @      �?      ;@      �?              @              0@      @              �?      @      >@      @      �?       @      @      3@              �?      �?      @      6@      �?      �?      @      @      =@      �?              �?              5@              �?      �?      @      :@      @                      @      3@      @      �?      �?      �?      >@      @               @      @      6@                      �?       @      >@      @              �?      @      1@       @      �?      @       @      ;@      @      �?                      :@      @      �?              @      3@      �?      �?      @       @      0@              �?      @              3@      @      �?      �?      @      6@              �?      @      @      1@      @      �?      �?      @      1@      @      �?      �?      @      8@      @                      @      :@                                      7@                              @      :@      �?      �?      @      �?      5@              �?                      8@      �?              @      @      A@      �?      �?      @      @      ;@      �?      �?       @      @      1@      �?                              2@              �?      @      @      2@              �?      �?      @      8@      �?              @              2@                                      6@       @              @      @      6@              �?      �?      @      =@       @               @      @      =@      @      �?      �?              4@      �?      �?       @      @      :@      @      �?      @      @      4@      @                      @      6@       @      �?      @      @      8@       @              @              3@              �?      @      @      8@       @              @      �?      6@      �?      �?       @      @      2@      �?      �?      �?       @      4@      @              @      @      8@              �?       @              3@      �?      �?      �?       @      0@       @      �?       @              3@      �?      �?       @              :@       @      �?      @      @      9@      @              �?      @      4@      �?      �?      @      @      ;@      �?      �?              @      8@      @              @      @      2@      @              @              6@              �?               @      7@              �?      @              0@      �?              @              ?@      �?                              5@              �?      �?      @      <@      @      �?      �?              1@       @      �?                      ;@              �?      @      @      6@      @      �?      �?              @@              �?      �?              5@      �?              �?              :@      �?      �?              @      3@      @      �?      �?      @      3@      @      �?      @      @      1@      �?              @      @      1@      �?              @              2@              �?      @              0@      @      �?      �?      @      7@      �?      �?              @      7@      @      �?      �?      @      3@                      �?              <@      @              �?              >@      �?              @      @      4@       @              @       @      1@      @      �?      �?       @      5@       @      �?      @      �?      4@      @      �?      �?      �?      2@      @      �?      �?      @      7@       @              @              7@      @      �?       @      @      2@       @              �?       @      5@       @      �?      @      @      2@      @      �?      �?      @      4@              �?      @      @      5@      �?              @      @      1@                      @      @      1@      �?              @              1@      @      �?       @      @      4@      @      �?      @              0@      �?              @      @      4@              �?      �?      �?      4@      @      �?              �?      =@      @              @              2@       @              @      @      0@       @              @      @      1@       @      �?       @      �?      :@                              @      2@      �?      �?              @      <@      �?      �?                      2@      �?              @       @      3@              �?      @       @      3@              �?      �?      @      3@      @      �?       @      @      7@                      @              1@              �?       @      @      0@      �?              @      @      1@       @              @      @      1@      @              @      @      3@      �?                              6@                       @              ;@       @              @      @      5@       @              @              6@                      �?              4@      @      �?       @      @      5@      �?      �?              �?      7@      @               @      @      3@      �?      �?      @      @      1@      �?      �?       @      @      9@      �?              @      @      4@      �?      �?      @      @      2@       @      �?       @              ?@      @              �?              3@              �?       @      �?      3@      @      �?      @      @      7@       @              �?       @      5@      �?      �?      @       @      1@      @      �?      �?      @      7@      �?      �?      @       @      3@      @              �?       @      ;@      @              @              4@      @      �?      �?      @      7@      @      �?      �?              5@      �?      �?              @      8@      �?               @              8@      �?      �?      @      @      5@      @              �?              2@              �?       @              1@       @              @      @      5@      @      �?      �?      @      <@              �?                      0@       @      �?      �?      @      6@                      @      @      1@       @              �?              6@      @              @              9@      �?      �?      �?              9@      �?      �?              @      5@       @      �?       @      @      3@      �?              @      @      4@              �?       @              =@      �?      �?       @      @      1@                      @              6@              �?      �?      �?      ;@      @      �?       @       @      =@      �?      �?      �?       @      ;@      �?              @      @      7@              �?              @      2@      �?      �?      @              1@      @              @      �?      6@      �?      �?      @       @      ;@      �?              �?              5@      @              �?      @      4@      @      �?      @              6@       @      �?      @      @      9@              �?                      ;@      �?      �?       @      @      3@      @              �?              6@       @                       @      4@      �?              �?      @      0@              �?      @              1@                       @              ;@              �?       @      @      2@      @      �?      �?      �?      8@      �?      �?      @      @      0@              �?              @      3@      �?      �?      @       @      5@      @      �?      �?      �?     �@@      �?              �?              <@       @      �?       @              4@      @              @      @      2@      @                              3@      �?      �?      @      @      3@              �?       @      @      1@              �?      �?      @      4@                       @              :@                              @      1@                      �?      @      3@      @      �?      �?      @      6@      @               @      @      8@      @      �?      @       @      8@              �?      �?       @      =@      @              �?              6@              �?       @      @      3@       @              @              2@      @      �?      �?      @      1@              �?              @      6@              �?      �?              5@              �?       @              0@              �?      @              1@              �?                      7@       @      �?       @      @      5@      @      �?      �?      @      8@              �?                      3@      �?      �?      �?              3@                      @      @      ;@       @      �?      �?              4@      �?              @       @      0@      �?      �?      �?              3@       @      �?       @      @      3@      @                      @      6@       @               @              :@       @      �?      @      @      4@       @              @              1@       @      �?      @              2@      @      �?      �?      @      <@              �?               @      5@      @      �?      �?      @      4@                      @      @      7@      @              �?      @      B@       @              @              2@       @              @              9@      @      �?      �?              :@      @              �?      @      4@              �?      �?      @      7@      �?      �?      @      �?      9@      �?      �?       @      @      1@      �?      �?      @              7@      �?      �?              @      >@              �?      @      @      9@                      @      @      0@              �?      @      @      2@              �?      �?      @      <@      �?              @      @      2@                      �?      @      6@      @      �?      �?              9@              �?      �?      @      :@      �?              @              3@      �?               @              6@      �?      �?                      A@      @      �?       @              2@       @              @      @      4@              �?      @      �?      <@      �?      �?      �?       @      =@      �?      �?      �?      @      9@                              @      0@      �?      �?      �?      @      ;@       @      �?              @      1@      @              �?              2@      @      �?              @      2@      @      �?      �?              ?@      @      �?      �?              6@                       @              2@      �?      �?              @      2@              �?      @       @      <@                       @              8@      �?              @              4@      @               @              0@      �?              �?              <@      @      �?      @       @      5@      @      �?      �?              6@              �?      �?      @      4@      @              @       @      2@      �?              @      "@      5@       @      �?      @       @      6@      @              �?              4@                      @      @      <@              �?              @     �A@      @              @       @      :@      @                      @      0@      �?      �?       @       @      ;@      @              �?              3@      �?              @              5@              �?       @      @      0@                      �?              4@       @              @      @      2@      @      �?      �?      @      8@      @               @      @      =@      �?      �?      �?              8@      @               @      �?      5@      @      �?      @      @      3@      �?      �?       @      @      3@       @      �?              @      4@       @              �?      @      @@      @      �?              @      3@      �?              @              :@              �?      �?      @      7@      @      �?      �?      �?      1@                      @      @      :@              �?      �?      @      8@      @      �?              @      3@       @      �?      �?      @      7@                      @      @      1@              �?      @              3@      �?      �?      @      @      :@      �?      �?       @      "@      1@              �?       @      @      4@      �?      �?      @      @      A@      @      �?              @      3@       @              @              2@              �?      @      @      0@       @      �?       @      @      7@       @      �?               @      1@      �?              @              :@      �?      �?       @              3@              �?      @              4@      @               @      @      :@      @              @      @      0@                      �?      @      8@       @      �?      @              8@      �?              @              9@       @      �?      @       @      1@                       @              7@              �?       @              :@      @      �?              @      3@       @      �?      @       @      4@      @      �?      �?              9@              �?      @      @      <@      @      �?      �?      @      2@              �?      @      @      1@      �?               @              2@      @      �?      �?       @      7@      @      �?              @      6@                      @      @      9@                      @      @      2@              �?      @      �?      :@      �?              @      @      6@      �?                      @      @@                      �?              8@      �?              @              >@              �?       @              1@      @      �?      @      @      7@              �?      @       @      9@              �?      @       @      3@              �?      @      @      6@      @      �?      �?      @      6@       @              @      @      1@      �?              �?       @      =@       @      �?       @      @      6@      @              @              1@      �?      �?      @      @      6@      @      �?      �?      @      5@      @              �?      @      3@       @      �?       @      @      9@                      �?      @      7@       @      �?      @              7@       @              �?      @      4@      �?              �?      @      5@              �?      �?      @      2@      �?               @      @      ;@              �?       @       @      1@              �?               @      8@       @      �?      @      @      7@                      �?              4@              �?      @      @      8@      @      �?                      2@              �?      @      @      <@                      @      @      6@      �?      �?               @      7@              �?      @       @      9@              �?              @      5@      �?      �?      @      @      5@              �?      �?              >@      @                      @      6@      �?      �?      @      @      3@       @              @      @      :@      @      �?                      0@       @      �?       @      @      ?@      @              �?      �?      1@      @      �?              @      9@      �?                              2@              �?      @      @      >@      �?      �?       @       @      >@              �?      @      @      1@      @              @              0@      @              �?      @      4@      �?               @              0@       @              @              8@      �?              @              2@              �?      @      @      3@       @      �?      @      @      6@      @                      @      2@       @              @      @      8@      �?              @              A@      �?      �?       @      @      2@      @      �?      �?              3@       @      �?      @      @      7@      �?              @      @      3@      �?      �?      @              0@      @                       @      1@              �?       @              3@      @      �?                      8@       @                              6@      @      �?      �?              0@              �?      @      @      2@              �?      �?      @      5@      �?      �?                      >@      @      �?      �?      @      :@      @      �?              @      1@       @      �?      @      @      9@                       @       @      2@      @                              0@              �?       @              6@      �?      �?      �?      @      8@      �?      �?       @      @      6@       @              @              0@                      @      @      2@      �?      �?      @              2@      �?              @      @      =@      �?               @              6@       @      �?      @              4@      @      �?      @       @      2@      @      �?      @              1@      @               @      �?      5@       @              @              5@���      �t�bhhK ��h��R�(KMI��h#�BHz  �      8            �       �       &      �      s      �       !            ;      �       ~             �       W      �      '       �             )      �       )      �             �      	      7      @      `      �      �      �      �      n      s      �      �      f      �	      	      �      7      �      x      +      �      G      �      �      �
      �                          H            F      �      M      �      �      �      <       7            �      [      �      h      :	      H
      �
      �
      q      p      K       �      �            .      X      �      �      �      Y      �      �      �      �      �      �      {	      �      �      �      �
      �      �      U      �      P      4      �      :      :      ]            ~      �      �      u      �       �      �       �      �      �      �      �      >      �
      �      X      y      v	      �             �      �      ;      f      5      �                  Y      �             (       S      �      �            �      a      �	      �      �      /      �       R      �      E      U      �      R      Z      x      �            �                  q      8      �            �      
      �                  �       X             �      p       �       �            p      �      �      %      %      �      �      �      �      "             �      J      w      	      �      �      �      (            �      6      �
      `      �       s       �      =      �             �      �      �      	      #	      I	      �	      +
      T
      b
      f
      �
      �
      F      v      �      �      �      �      +      1      <      [      �      �      3      �      �      �      �            3      F      �      i             �       �       k      }            �      5                  �      �      �      �      |      �      �      p      �      �      w            �      �       R      �      �      �            8      E      u      �      l      =	      a	      '      a      �      u      ;      �      ;      �             M      �      �      '            V      �      �      �      �            4      �      O      �      	      A	      Y	      �	      �	      �
            �      �                  �      !       	       �             �       �       #      E      �            �      �            :      B      M      �      �      N      �      �      x	      d      m      
      J       t      �
      ^      0      �	      �       �      ]      7
      
      B      &      �            Z      6	      	      �      �      �      �      �	      �	            ^	      7      �
      �
      �            4      `      �      L      /      �      �      R      5             v      �      �      �      �                  �      %      U      }      �            �      �      >      _      N      U	      ^      �      
      o      S      �      �      �      �      g      �      	      �      _      �      D      K      /      �      �	      �      Y
      �      �      V      �       �      �      6      �      �       �      i      �      P      �      0      c      �              G            �	            �      V      �      �      �      _      �      �      �      ;      j      m      p      v      �      �      �      �      �            +      ]      �      t      �      ~      �      �      �      %                   c      �      �      x      z             v      �      �
            �                        g      �      �      �      �      b	      �      �      �      �      �      �	      �            9      h      s      �      q      Q       �            �      �      �             *      y      �      j      )            C      �      �      c      d      Y            �      �            H      a       3      �      �       �      1            �      ^      �            �            )      H      �      �      �      y      ~      �      �	      �      t            "
      �            �            �	      0      �
            N
            #      8      �      y      �       �      U      '	      �      �      Y      F      	      �      �      �      �       �      
      y      >      8      >      &      �      �      �      �      6      Y       �             �      .      y      �      �      q       �      s      d      �      �      �      �      $      �      �      �      �      �      �      �      n      �      G      �      �      Z      V      r      �      �      =      p      r      �                  ,      G      S            w      �      �      �      	      %	      ~	      �	            �      �      T      !      "       �      c      �      �       �
      �      �      r	                  �      l      �
      �
      6            %      q      �      �      �      �      +      �      �      �      �      �      �      �      T      s      z      �      R      �      �      �      �      e      y      �      @
      �
             
      �      �      �      [                  �      ?      �      �             �            �      a      �	      �      =      �      �      �      �            #      �      j
      Y      A                  �      �      �      �      C      �                  J      �      �      �	      �	      
      A      _      k      A            �      %       �       J      �      s      �      b                  �      �      �      �      �      �	      �	      �
      �      )      �      �       �      y       N      �       K      �      �      f       �            V
            �      �      �      �      b      �      Z
      �      5      w      �             w      �       5      k      �      �      �      �      )	      �      .	      �	      �      B            �      \      �      �      H      �      �      �      \	      �	      :
      �
      N      �      /      f      �            �      �      �      �            Z      x
      �                  �      �            �      �            �      �            �       q      �
      �            ;      �      d
      9      g      �      k
      m      8	      r             ]      �	      4	      �      &	      j      �            )      �      �      �      �      �	      0
      a
      �      `      �      �      �      �      _      a      �            �      �            X            t      �
      �      �             <      L      �      �      �      �      u      L      	      "      �
      +      l      1      '      �	      �      �      �      �      r      �      z      t	            
      �      $      A      E      N       _      j      �      �      D
      ~      �      �      4      a      �            +      n      N      |      �      <      q      �                  �      �	      �      -      D      j      b            �            G      �      Z      �      �      -      )      �      3      �      0      �       	      �      w       �      ;      D            �      �       �            �	            {      :      �      �       S	      �      O            }      �      �      
       �       e      �            �      H      �            d      B            $      �      "      �      m      �      _      
      �      =      ?      B      �	      �      �      *	      G      �      �      �      j       �              	      �       =       g      (      .      k      Q      �      g      �      �      �      �      ~      �      s      I      �      �      x      �      y      �      7	      �	      �	      %
      s
      ~
      �
      �
      �      5      �	            �      �      E      �      �      �      O	            �            6       �      �            �
      �      $      �      �       8      {      �	      P      '      ?	      W      z      ]      �      �      8      �      �      �            �      $	      p	      8
      ;
      �            1       g       �       0      e      o      �      �      .      
      �      �      O      e      �      �      ?      �      >      c	      `      c      �      b      �            `      e      �      �      e      �      �      '
      ;      �
      }            �      �      �      �      �      �             7      �      �
      8            A      G      �      �      �      	      �                  �      e      %      �      <      �      �      �            +      8      W      �      �      �      6      �	            �      �      �
             �      �      �      &      (      !      %      �      �      �      w      y      x      �      ,      �      �      y      !      [      �      �      `      �             �       �	      �                  B       �      �      ]      �      �      (      z      �      W      �      <      �      H      k	      �	      �       �             (            0            b      *      �      �      �	      
      �      �      �      P       �       �       v      �      �      6      d             
      h      �      _      r      F      �      	      �	      "	      
      �      �	      `
      D       3      c       �       b      �      �      �      ~      �      n       M      �      �      �      a            �      �      }            �      v       ;       �      �      I      �      �      g      v      �      }      ?      K      �      �      Q	      F                   �            \       �             �      '      Q      =      �            �      �      -      B      �      �      	      �      �      g
      �      �
            x      5      �      R       \
      d      �      	      =      �      �            �      \      �                  h      �      �      �
      �      �       �      "      3      �      A      S      �      �      �      2       �       �       [      0      h      K      v      �      R	      ?
      �
      -      W      w      �      +      �      m      W      �      �      ?      O      �      �             Y      u
      �
      �
      �            �      �       x      �      
      �      �      �      	      �      �      �      �      �      �      O      �      /      �      P            �	      �
            �      >      �      Z                    P            �      �      7      g      |      �      �
      �
      ;      �      \      �      �      �      �      �                  L      �      �      �      �       �      �      �      �      �      �      ^      a      �      �            K	            �      �             Z      �      �      �      �      �      �      �      A      �      �      	      m      �      �      �      4      D      �      �      �      �      �      �      �	      �
      �
                   I       �       �      �                  �      �      �      �      .      �            �      �      {      �      a      �      �      �             �      
      �      �      �      �      
      l      �      �      �      �      �             Q      V      �      �      7      �      �      �      �      �      �            0      �      �       �      n      Q      �      �      �       �      �      �
      �      �            �      ,
      �                  h      �      �      z      U      &      �      �      �      �      !      �      E      t      3      a      #       �      #      �      �       �      �      �      /      +      -      �      h	      �	      �
      �
      C      �      �            �      �      �            �      �      �      �            �      �      �       �       "      �	      |      =             |	      �      �            
      j      �      i            ,      s      �            �	      �	      
      �
      �
      �      �      S      o      �      @      O      �      .      &      2      6      �      �      �      "      �      q      �	      ]      �      k      |      �	      �      �	      2             �	      a      �      �      �       B
      )
      %      �
      N      �      �
      �      �
      �      �      �            �      ?      6            �      {      F      
      2      s	      M      2      �      �      Z      �      a            @            �      r      �      �      �      �      q      k      �       �            �      ^      �            V      y	      �	      <
      f            �      �      �      ^      4      �       �      �      �      �      
      #            �       T      c            �
            �      t      ?      �      �      �      A      `      �      �      �      A      �      �       �             
      4
      �      �      �      d       *      �      n      R      �      0      J	      �	      �
      �      �            �      �      �      �      W      �      C      1      
            �      �      �      �      >      �      �      �	      *      �      �            �              {      k      x       �      V      �	      `      �      �	      q      �      /
      �      -
      �      o      !      �      �             :      �      �      4      |       �      �            /      �      v      �       �      �	      �      p      �      e       u      T      �      �      �	            V      �      �             �      �      K      ]      D	      f      <      %      @                  &      6      �      �      ~      C       6
      @      !      %      �
      �      �      z      v      V       M
      T      �      �	            �      �
      \      	      �	      [      X      �      	      	      �	      �	      
      >
      �
      �
            �      �      �      �      �                   9                        '      r      #      �
      �      �	      "      ^      �      9      ?      �      �      �      W       -      �      �
      �      �	      5	      	      �            �      �      ~      c      �      �            �	      l
      �            �      �      �       9      �      �      D      1      J      �      �      �	      !
      q
      �
      �
      �      �      )      -      M            9       �       ,      t      x      �            Y      u      �      _      H	            �      <      #      u	      �      �      L      �      A      �      �      �            3      e	      
      �
      �      �
      b      �             (      R      �      �      �      �      �      �            K      o      r      �      �      S      �                  _      �	      �      �      T      �
            ^
      
      *                        (      q      x      :      �      1      B      �      �      c      f      �      �      O      �      �      �                   /       ]       �       �      �      K      S      l      �      �      �      �       Z      -       !            �      \      �	            �      7      �
      �	      J      /      A      �      �      �	      �      W	      r      -            �            	      |      X      �      I            5      �      O      \      �      �      �      �            J      �      ^      �      �      n      �      �      �                  u      �      �      �            �      R      H      n      :      Q      j      �      �      2      �       �      4      !      W      h      m      C            �       8      3      �	      �      [       >       \      �       �      $            �      �      �      �      M	      V	      w	      �
      �
      �
      �
      T      �      �      8       (      �       �      �      �      �      �                  K      �      �      t       Q              �      +      �      �      &
      �      '      z       �       �	      �      1      �      �            �       [	      <	      	      @      �       P      �      �      e
      n
            /      :      D      �      �      �      r      �      D      E      U      1      �      �      �      �      <      C      �      E       4      �       s      ,      �      �      %      �            Q      ~      �      	      =      _       �
      .      Z      �      p      :       �      G      �      �      �      n      �      �      k            �      �      u      M      �      �	      �	      �      )      �      �      C      N      u      w                        �      �      M      h      �            �      �      �             �      ?      �      	      0	      �	                  g      �            �      #      I      �	      H      �
      �
      �      �
      7      �      &      U       �      d      �      6      F            �      �      �      C             I      �      w                  B	      �       &      �            �      �            �      �	      �	            M      R      �      I      �      B      �      �      i            �      l            -      ^       o      )      V      ,      e      �      
                  �      ^      �      	      �      �	      �	      F
      �      2      }	      �      �      ?      �       �      �             7      T                  X       o       �      r      #
      �
      L      �      E	      @      �      �      �      �      �      !      �      �      �            6      �      �            �      �       �       �      [      w
      �
      a      �      |      �      �      	      /      �            [      �            �      �            ?      =      D      �            �       
      �	      b                  n	      :      �      F      `      �      �      �	      �	      p
      �
      �
      1      �      �      �      �      K      �      �      �      	      	      �	      I
      �
      }      d      �             U            0      �
      C      +      �      Q      ,      �      �            *      /            -      J      2      �	      c            �
            �      v      f      �      �       �      |      �             �      f      �      �      �      �      :      �      �      O      Q      �      �      M            �      �      �      �      �            f      w      �      �      �	      r
      �
      E      G      7      �      !      �      G      �      �	      �
      �      2      F      �            ,      ]      �      t      �      �      $      `      l            ?       �             �      "      �
      �
            �      �      �                    G      j      �      �      �      9      g      #      �      �      �      >      �      �	      o
      �
      2      S      �             �       �      �      �      o	      q	      �	      �	      �	      n      �	      O
      R            G      �
            �      *      �      �      �      &      >      �       �      �      X      c      �            �       �      V      9            �	            		      �      �      n      �      �      �            5      �      �      �      �      	      {      �            C      \      �      .      �      8      �      �      �      �      �      1      �      M      �      
      L            @	            �	                        �	             I      �      K      �       �	      �	      Q      	      �      -      �      �      �            �      _      �      �      z
      �      �	            �      �             p      �      �      �      �      .      E      N      �      �      '      (	      �	      �	      �
      �
      �
            �      �      _      s      �                   1	      T	      �
      Z      p      �            0      j      �      �      l                  �      9      �      .      m      1      �      �      �      C
      }
      �      �            �      �      �      �      F      z      �      �      �            �       �      �            �      �      .      �	      
      �
      �
      �
      d      F      �      �       A            {      b       3      �      
      j	      A       @      5      O       &      �	      �      �      
      b      �
      '      d                  �      
      �       �
            �      �      e      �      �      �      �      �      {      �      �
      l	      �      E      N	      �      �      �
      �
                  $      �      >      T       {       m      �      �            �      �      G       	      �            �	      �      �      �      ]
            #      �	      �      }      �      \      l      z	      �      J             g      >      �      3      �      �      �      �      �      Y      �      9	      2	      h      �      �      i            �      ,            �      �      �      
      3
      t      �            7      g      2      �      �      (      k      �            D      W      �            ,      �	            �      �      �       �
      �      �      ^            Z	      H      �      �      
      9            V      �      �      *       �      �      �      N      $       4            b      �
      g      B      �      �       3      �      �      *      �             �      �       '            h      S      W      %      q      �      H      �      <      �      �      o      �            P      �      3      8            i            s      �      �	      �
      �
      e      .       @       `       �       i      �      �            �            4       H       l       �             b      
      `      �      /      O      p      �            �      E      �      *      P      �      �      �            ;	      �	      
      �
      �
      ,      �      �      �      �            B      �      �
      �      �      1      �
      �       2      �      �      �      �      �      �      �      �      "      �
      i      �      �      =      �      �      �            M      �      �      c      &      �      �
            �      �       �      �	      �      	            �      �             n      �      �      f      �                    Z      �      2
      �      �      �      (      2      >      �      �            o      �      �      �      �
      �            }      {      �      �      }      �      �      ,      T      �      �      �      J      �      �      �      F      #      '      �      �      �      \      �	      ?      |      �      d      l            �            �      I      �      �      �      �
      h      w      �      }       �       �       �       ;      <      �      �      �            L      
      �      �      �      �      �      �      �      �      �      f	      1
      �      �            �      �      �      ;      �      �      �      �      �      �      �      5      "      9      �            �      V      �       �
      ,       �	      	      >      �	      <      i
      �       5      �      �
             W
      �      T            Y      m	      �
      P      �      �      �      �	      J
      �       r      |      �      �            x      E      �      U      �      c      i      p            
      �      �      �	      �      i	      �      �
      �
      Q
      �      �      y      |      �      <      P      �      �      �      �      �      [      �      i      �      	      �	      �	      	      �      �      }      �      �       O      K      (      �      �      G	      G
      �
      �       �      �            X      l      �      �      '      0      �            $      X      �      0            �      C	      
      t
      �      P      �            y
      v
      i      $
      �      "      �      z      �	      �      �      7      L	            
      �      �      n            !      4      9
      �      9      L                        &       0       �       �      y      �      "      �      �      �      v      �      �      �      >	      �	      �
      j      o      A
      �      �            S      U      2      �            W      5      =             W      �      �      �      =      �      )             �      	      �      H      9      =
       
      �      /	      �      (      �      �      r      �      �	      +      �      �      �
            �      �      (      N      �       �      L
      �      B      �             �       �      �      �      :      R      �      �      �      �      $      �      g	      �	      �      �      	      �            �      �      X
      �	      �      �      �      �      j      �      �      �      !      �      	      4      .      �      �      �      �      J      U      D      ]      \      O            U      �
      j      �      �      {
      �
            I      T      s            
      L      �      �      q      $      I                        :             �      �	      �      �      f      �      Q      �       �      �       $      X      �      �      �            %      �            �      �      C      E      \      i      �      �      �      �
      �      �      �	            �            f      �                         �      �      -      t      �            @      D      U      �      �       �       �      �      J            e             �      �      �      �      	      �      ^      m      �      �      �      �      �      �      x      J      �      �      �      U
      m      h
      �      �      D      �	      �      �      �       �      u             h       �
      +	      H      @      �      h      =      |
      ]             
      p      �	      �      k      A      �       �      �      �            �      �      �      �      �            P	      �	      

      S
      [
      [            I      �      �            �      �                  �      C      �            P
      R
      9      {      �      �             Q      �      �      ,      B      �      �      �      �      m
      t      �      6      �             C      �      �      �            +             �      L      �      �      S      k      �      �      �       Y      �      *      w      �      �      m       �            �      	             �                  	      u      �      �      B      ^      v      T      7       o      d      �      �      &            �      ]	      _	      (
      6      /      �      �            R      �      !	      X	      �	      �	      .
      �      ;      �            �      '      Y      o      �      b       	      F	      d	      �	      5
      E
      3       D      �      �
      �      �       �      k       �      +      P      �       X      ]      �      �      N      �      �      �      ~      z      �	      #      
      *
      �      c
            �
      �      
      �
      ?      �            �            }      �      �      �      �            )      �
      �       1      �      u      �      �      �            X      �      $      �      �      �      �      �
      $      #      {      [      �      8      �      Y      i      L       �      m      �                  [            K
      �      o      e      *      	      �      )      �
      S      �      I      �      -      �      5      _
      �      �      �      �      �      H      �      M       �      �       �      �            �      .      �            t      -	      �	      �      �      :      ~      *      <      �            4      S       �      �       u       �      �       @      "      N      �
      �      �      |      {            ~      �      �      �      �      �            �      @      K      �      �      �                   �      �            �      �      �      �      *      �      �      �      )      �      F      z      �      �      
	      �	      ;      L      �            �      �      G      �      3	      �      �      �      x      �      �      z            �      l      �      k      @            �	            �      `	      �
      �      �      �      Z      ,	      	
      �
      �
      �t�bhhK ��h��R�(KK���h �V32�����R�(K�|�N(�	idx_start��idx_end��is_leaf��radius�t�}�(hah#K ��hbh#K��hch#K��hdhOK��uK KKt�b�B�          I              �:r�(@        �              ��S°@�      I              g��U�#@        �              @���I@�      �              ��6ҭ�@�      v              F�\��i@v      I              /Y˿�!@        �              ��v �@�      �              ���/�@�      �              �/7�R@�      �              .!	��@�      �	              ���!Ȍ@�	      v              �/_ee@v      _              F�\��i@_      I              �NO���@        �               9�c��T@�       �              �;f��@�      �              ����R@�      �              ��Z���@�      �              S[�:XL	@�      �                    @�      �              htN�=@�      �              �.�!hp@�      �              �;f��@�      �	              ��v �@�	      �
              ۞[E~�@�
      v              ����w�@v      j              ���!Ȍ@j      _              �/_ee@_      T              ��b�n�@T      I              ȭ��~@        z               �٨�h�@z       �               �9B.��@�       n              �Md4�o@n      �              �9B.��@�      c              �9B.��@c      �              �Md4�o@�      W              �;f��@W      �              .!	��@�      L              .!	��@L      �              �Md4�o@�      @              `�*�:
@@      �              �LX�z�@�      5              ��ci3�
@5      �              S[�:XL	@�      )              	Ў���@)      �                    @�                    �9B.��@      �              .!	��@�      	              9�c��T@	      �	              �;f��@�	      
              �9B.��@
      �
              ��Z���@�
      �
              ��v �@�
      v              ��v �@v      �              �;f��@�      j              ��v �@j      �              I?h��@�      _              ����w�@_      �              �l��v�@�      T              @���I@T      �              wIs �@�      I                    @        =               ���T@=       z               �Md4�o@z       �               �Md4�o@�       �               �f~ @�       1              4o��r��?1      n              I?h���?n      �              I?h���?�      �              �VTY��@�      &              �Md4�o@&      c              �VTY��@c      �              4o��r��?�      �              I?h���?�                    .!	��@      W              �9B.��@W      �                     @�      �              �Md4�o@�                    �Md4�o@      L                     @L      �              4o��r��?�      �              I?h���?�                    �VTY��@      @              �VTY��@@      }              �;f��@}      �              �VTY��@�      �              ���T@�      5              �٨�h�@5      r              �Md4�o@r      �              .!	��@�      �              `�*�:
@�      )              ��v �@)      f              S[�:XL	@f      �              �LX�z�@�      �              �l��v� @�                    �9B.��@      [              �NO����?[      �              .!	��@�      �              �9B.��@�      	              �٨�h�@	      O	              .!	��@O	      �	              �9B.��@�	      �	              �VTY��@�	      
              �Md4�o@
      D
              .!	��@D
      �
              �;f��@�
      �
              �;f��@�
      �
              9�c��T@�
      8              �;f��@8      v              �;f��@v      �              �9B.��@�      �              .!	��@�      -              .!	��@-      j              4o��r�
@j      �              .!	��@�      �              �٨�h�@�      !              ��v �@!      _              ��v �@_      �              �Md4�o@�      �              ۞[E~�@�                    ��ci3�
@      T              ����w�@T      �              	Ў���@�      �              �/_ee@�                    �.�!hp@      I              ST����@                      �LX�z��?       =              ���T@=       [              4o��r��?[       z              4o��r��?z       �              I?h���?�       �              4o��r��?�       �              �f~ @�       �              S[�:XL�?�                    ��ҩ*�?      1             4o��r��?1      O             4o��r��?O      n             4o��r��?n      �             I?h���?�      �             S[�:XL�?�      �             �YaD+��?�      �             �VTY��@�                   4o��r��?      &             I?h���?&      D             I?h���?D      c             �f~ @c      �             ��ҩ*�?�      �             4o��r��?�      �             4o��r��?�      �             4o��r��?�      �                    @�                   �Md4�o@      8             �Md4�o@8      W             �VTY��@W      u             �;f���?u      �             4o��r��?�      �             4o��r��?�      �             I?h���?�      �             I?h���?�                   4o��r��?      -             �;f���?-      L             4o��r��?L      j             �;f���?j      �             �;f���?�      �             I?h���?�      �             S[�:XL�?�      �             S[�:XL�?�                   �f~ @      !             4o��r��?!      @             �f~ @@      ^             �Md4�o@^      }             �9B.��@}      �             �f~ @�      �             I?h���?�      �             �YaD+��?�      �             4o��r��?�                   ���T@      5             .!	��@5      S             S[�:XL�?S      r             I?h���?r      �                    @�      �             �Md4�o@�      �             �VTY��@�      �             �9B.��@�      
             �;f��@
      )             9�c��T@)      G             �Md4�o@G      f             �Md4�o@f      �             �VTY��@�      �             �;f��@�      �             �YaD+��?�      �             ��ҩ*�?�      �             �VTY��@�                   �Md4�o@      <             S[�:XL�?<      [             ��ҩ*�?[      y             I?h���?y      �                    @�      �             �l��v� @�      �             �9B.��@�      �             ���T@�      	             .!	��@	      0	             �LX�z��?0	      O	             .!	��@O	      n	             �l��v� @n	      �	             �9B.��@�	      �	             �f~ @�	      �	             4o��r��?�	      �	             I?h���?�	      
             4o��r��?
      %
                    @%
      D
             �Md4�o@D
      b
             �Md4�o@b
      �
             �9B.��@�
      �
             �9B.��@�
      �
             .!	��@�
      �
             .!	��@�
      �
             �;f��@�
                   .!	��@      8             �VTY��@8      W             �Md4�o@W      v             �9B.��@v      �             �YaD+��?�      �             �9B.��@�      �             S[�:XL�?�      �             .!	��@�                          @      -                    @-      K             4o��r�
@K      j             wu�.@j      �                    @�      �             �Md4�o@�      �             .!	��@�      �             4o��r��?�                   9�c��T@      !             �;f��@!      @             �;f��@@      _             9�c��T@_      }             4o��r��?}      �             I?h���?�      �             �Md4�o@�      �             �LX�z�@�      �             �٨�h�@�                   .!	��@      5             �LX�z�@5      T             �C-�Ґ@T      r             .!	��@r      �             ��ci3�
@�      �             I?h��@�      �             �)�0+@�      �             ��hdE@�                   �YaD+�@      *             �6��?@*      I             �m�ܩ@�t�bhhK ��h��R�(KKK�K��hO�B�O                                        0@                                      0@                                      5@                                      0@                              @      0@                                      5@                                      8@                                      0@                      @              0@                              @      0@                       @      @      0@                                      5@                              @      5@                                      8@                                      ;@                                      0@                                      3@                      @              0@                      @              2@                              @      0@                              @      0@                       @      @      0@                       @      @      0@                                      5@                       @              5@                              @      5@                       @      @      5@                                      8@                              @      8@                                      ;@                                      >@                                      0@      �?                              0@                                      3@      �?                              3@                      @              0@                      @              0@                      @              2@                      @              2@                              @      0@                              @      3@                              @      0@                              @      0@                       @      @      0@                      @      @      0@                       @      @      0@                      @      @      0@                                      5@       @                              5@                       @              5@                      @              5@                              @      5@                              @      5@                       @      @      5@                       @      @      5@                                      8@                       @              8@                              @      8@                      �?      @      8@                                      ;@                              @      ;@                                      >@                              @      >@                                      0@                      �?              0@      �?                              0@      �?              �?              0@                                      3@                      �?              3@      �?                              3@      �?              �?              3@                      @              0@      �?              @              0@                      @              0@      �?              @              0@                      @              2@      �?              @              2@                      @              2@      �?              @              2@                              @      0@       @                      @      0@                              @      3@      �?                      @      3@                              @      0@                              @      3@                              @      0@                              @      3@                       @      @      0@                       @      @      2@                      @      @      0@                      @      @      2@                      @      @      0@                       @      @      0@                      @      @      0@                      @      @      0@                                      5@                                      5@       @                              5@       @                              5@                       @              5@       @               @              5@                      @              5@      �?              @              5@                              @      5@       @                      @      5@                              @      5@                              @      5@                       @      @      5@                      @      @      5@                       @      @      5@                      @      @      5@                                      8@       @                              8@                       @              9@                      @              8@                              @      9@                              @      8@                      �?      @      8@                      @      @      8@                                      ;@                      �?              ;@                              @      ;@                      �?      @      ;@                                      >@                      �?              >@                              @      >@                      �?      @      >@                                      0@                                      0@                      �?              0@                       @              1@      �?                              0@      �?                              2@      �?              �?              0@      @              �?              0@                                      3@                                      3@                      �?              3@                       @              3@      �?                              3@      @                              3@      �?              �?              3@      �?              �?              3@                      @              0@                      @              0@      �?              @              0@      �?              @              0@                      @              0@                      @              0@      �?              @              0@       @              @              0@                      @              2@                      @              2@      �?              @              2@      �?              @              2@                      @              2@                      @              3@      �?              @              2@      �?              @              3@                              @      0@                              @      2@       @                      @      0@       @                      @      1@                              @      3@                      �?      @      3@      �?                      @      3@      @                      @      3@                              @      0@      �?                      @      0@                              @      3@      �?                      @      3@                              @      0@      �?                      @      0@                              @      3@       @                      @      3@                       @      @      0@      �?              @      @      0@                       @      @      2@      �?               @      @      2@                      @      @      0@      �?              @      @      0@                      @      @      2@      �?              @      @      2@                      @      @      0@                      @      @      2@                       @      @      0@                       @      @      2@                      @      @      0@                      @      @      3@                      @      @      0@                      @      @      2@                                      5@                                      7@                                      5@                               @      5@       @                              5@       @                              7@       @                              6@       @                       @      5@                       @              5@                       @              5@       @               @              5@       @              @              5@                      @              5@                      @              5@      �?              @              5@      �?              @              5@                              @      5@                              @      7@       @                      @      5@       @                      @      7@                              @      5@      �?                      @      5@                              @      5@      �?                      @      5@                       @      @      5@       @               @      @      5@                      @      @      5@      �?              @      @      5@                       @      @      5@      �?               @      @      5@                      @      @      5@      �?              @      @      5@                                      9@                                      8@       @                              9@       @                              8@                       @              9@       @               @              9@                      @              8@                      @              8@                              @      9@      �?                      @      9@                              @      8@       @                      @      9@                      �?      @      8@                      �?      @      8@                      @      @      8@                      @      @      8@                                      ;@      �?                              ;@                      �?              ;@                       @              ;@                              @      ;@                              @      ;@                      �?      @      ;@                      @      @      ;@                                      >@                                      @@                      �?              >@                      �?              ?@                              @      >@                              @     �@@                      �?      @      >@                      @      @      >@      @      �?      @      "@     �B@      @      �?      @      "@      5@      @      �?      @      "@     �B@      @      �?      @      @      5@      @      �?      @      "@      5@      @      �?      @      "@      8@      @      �?      @      "@     �B@      @      �?      @      @      5@      @      �?      @       @      5@      @      �?       @      "@      5@      @      �?      @      "@      5@      @      �?      @      @      8@      @      �?      @      "@      8@      @      �?      @      "@      ;@      @      �?      @      "@     �B@      @      �?      @      @      3@      @      �?      @      @      5@      @      �?      @       @      2@      @      �?      @       @      5@      @      �?       @      @      5@      @      �?       @      "@      5@      @      �?      @      @      5@      @      �?      @      "@      5@      @      �?       @      @      8@      @      �?      @      @      8@      @      �?       @      "@      8@      @      �?      @      "@      8@      @      �?      @      @      ;@      @      �?      @      "@      ;@      @      �?      @       @      >@      @      �?      @      "@     �B@      �?      �?      @      @      3@      @      �?      @       @      3@      �?      �?      @       @      5@      @      �?      @      @      5@      @      �?      @       @      2@      @      �?      @       @      2@      @      �?      @       @      5@      @      �?      @       @      5@      @      �?       @      @      3@      @      �?       @      @      5@      @      �?       @      @      5@      @      �?       @      "@      5@      @      �?      @      @      5@      @      �?      @      @      5@      @      �?      @      "@      5@      @      �?      @      "@      5@       @      �?       @      @      8@      @      �?       @      @      8@      @      �?      @      @      8@      @      �?      @      @      8@      @      �?       @      @      8@      @      �?       @      "@      8@      @      �?      @      @      8@      @      �?      @      "@      8@      @      �?       @      @      ;@      @      �?      @      @      ;@      @      �?      �?      "@      ;@      @      �?      @       @      ;@      @      �?      @       @      >@      @      �?      @       @      >@      @      �?      @      @     �B@      @      �?      @      "@     �B@      �?      �?      �?      @      3@      �?      �?      @       @      3@      @      �?      �?       @      3@      @      �?      @       @      2@      �?      �?      �?       @      5@      �?      �?      @       @      5@      @      �?      �?       @      5@      @      �?      @      @      5@      �?      �?      @       @      2@      @      �?      @       @      2@      �?      �?      @       @      2@      @      �?      @       @      2@      �?      �?      @       @      5@      @      �?      @       @      5@      �?      �?      @       @      5@      @      �?      @       @      5@       @      �?       @      @      3@      @      �?       @      @      3@      �?      �?       @      @      5@      @      �?       @      @      5@      @      �?       @      @      2@      @      �?       @      @      5@      @      �?       @      "@      3@      @      �?       @       @      5@      @      �?      @      @      1@      @      �?      @      @      5@      @      �?      @      @      2@      @      �?      @      @      5@      @      �?      @      @      5@      @      �?      @      "@      5@      @      �?      @      @      5@      @      �?      @      "@      5@       @      �?       @              8@       @      �?       @      @      8@      @      �?       @              8@      @      �?       @      @      8@       @      �?      @      @      8@      @      �?      @      @      8@      �?      �?      @      @      8@      @      �?      @      @      8@       @      �?       @      @      8@      @      �?       @      @      8@      @      �?       @      @      8@      @      �?       @      "@      8@      @      �?      @      @      8@      @      �?      @      @      8@      @      �?      @      "@      8@      @      �?      @       @      8@       @      �?       @      @      ;@      @      �?       @      @      ;@      @      �?      @      @      ;@      @      �?      @      @      ;@      @      �?      �?      @      ;@      @      �?      �?      "@      ;@      @      �?      @       @      ;@      @      �?      @       @      ;@      @      �?      �?       @      =@      @      �?      @       @      >@      @      �?      �?       @      >@      @      �?      @       @      >@      @      �?      �?      @     �B@      @      �?      @      @     �B@      @      �?      �?      "@     �B@      @      �?      @      @      B@      �?      �?      �?              3@      �?      �?      �?      @      3@      �?      �?      @       @      1@      �?      �?      @       @      3@      @      �?      �?       @      2@      @      �?      �?       @      3@      @      �?      @       @      2@      @      �?       @       @      2@      �?      �?      �?              5@      �?      �?      �?       @      5@      �?      �?       @       @      5@      �?      �?      @       @      5@      @      �?      �?       @      5@      @      �?      �?       @      5@      @      �?      @              5@      @      �?      @      @      5@      �?      �?      @       @      2@      �?      �?      @       @      2@      @      �?      @       @      2@      @      �?      @       @      2@      �?      �?      @              2@      �?      �?      @       @      2@       @      �?      @       @      2@      @      �?      @       @      2@      �?      �?      @       @      5@      �?      �?      @       @      5@      @      �?      @       @      5@      @      �?      @       @      5@      �?      �?      @       @      3@      �?      �?      @       @      5@      @      �?      @       @      3@      @      �?      @       @      5@       @      �?       @      @      2@       @      �?       @      @      3@      @      �?       @      @      1@      @      �?       @      @      3@      �?      �?      �?      @      5@      �?      �?       @      @      5@      @      �?       @      @      5@      @      �?       @      @      5@      �?      �?       @      @      2@      @      �?       @      @      2@      �?      �?       @      @      5@      @      �?       @      @      5@      �?      �?       @       @      3@      @      �?       @      "@      3@       @      �?       @       @      5@      @      �?       @       @      5@      �?      �?      @      @      1@      @      �?      @      @      1@      �?      �?      @      @      5@      @      �?      @      @      5@              �?      @      @      2@      @      �?      @      @      2@      �?      �?      @      @      5@      @      �?      @      @      5@      @      �?      @      @      2@      @      �?      @      @      5@      @      �?      @      "@      2@      @      �?      @      "@      5@      @      �?      @      @      2@      @      �?      @      @      5@      @      �?      @       @      2@      @      �?      @      "@      5@       @      �?       @              7@      �?      �?       @              8@       @      �?       @       @      8@       @      �?       @      @      8@      @      �?       @              7@      @      �?       @              8@      @      �?       @       @      8@      @      �?       @      @      8@       @      �?      @              8@       @      �?      @      @      8@      @      �?      @      @      8@      @      �?      @      @      8@      �?      �?      @              8@      �?      �?      @      @      8@      @      �?      @              8@      @      �?      @      @      8@       @      �?       @      @      7@      �?      �?       @      @      8@      @      �?       @      @      7@      @      �?       @      @      8@      �?      �?       @      @      8@      @      �?       @      @      8@      �?      �?       @       @      8@      @      �?       @      "@      8@       @      �?      @      @      8@      @      �?      @      @      8@      �?      �?      @      @      8@      @      �?      @      @      8@      �?      �?      @      "@      8@      @      �?      @       @      8@      �?      �?      @       @      8@      @      �?      @       @      8@       @      �?       @              ;@       @      �?       @      @      ;@      @      �?       @              ;@      @      �?       @      @      ;@      �?      �?      @      @      ;@      @      �?      @      @      ;@      @      �?      @      @      ;@      @      �?      @       @      ;@      �?      �?      �?      @      ;@      @      �?      �?      @      ;@       @      �?      �?      "@      ;@      @      �?      �?       @      ;@      @      �?      @      @      ;@      @      �?      @       @      ;@      @      �?      @      @      ;@      @      �?      @       @      ;@      �?      �?      �?       @      =@      @      �?      �?       @      =@      @      �?       @       @      =@      @      �?      @       @      >@      @      �?      �?      @      >@      @      �?      �?       @      >@      @      �?      @       @      >@      @      �?      @      @      >@      @      �?      �?      @      @@      @      �?      �?      @     �B@      @      �?      @      @      ?@      @      �?      @      @     �B@      @      �?      �?       @      @@      @      �?      �?      "@     �B@      @      �?      @      @      B@      @      �?      @      @      B@�t�bKKK�M8=M?:M^rJ�� �sklearn.metrics._dist_metrics��newObj���ht�EuclideanDistance�����R�G@       hhK ��h��R�(KK��h �f8�����R�(Kh$NNNJ����J����K t�b�C        �t�bhhK ��h��R�(KKK��h��C        �t�b��bNt�b�_sklearn_version��1.1.3�ub.