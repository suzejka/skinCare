��rR      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K
�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�Ch                                                                	       
                     �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K	�
node_count�K}�nodes�hhK ��h��R�(KK}��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�BX         *                    �?�9�y���?�             c@                          �5@      �?0             H@                           �?�g��s��?             9@                           �?0�����?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @	                            �?h/�����?             2@
                           �?r�q��?             (@������������������������       ��q�q�?             @                           3@r�q��?             @������������������������       �                     @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                           3@9��8���?             @                          �1@VUUUUU�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                           �?�q�q�?             @������������������������       �      �?              @������������������������       �                     �?       %                     @|�!*�?             7@       $                   �@@VUUUUU�?             .@                          �6@VUUUUU�?             (@                           �?�q�q�?             @������������������������       �                     @������������������������       �                      @        #                   �8@r�q��?             @!       "                   �7@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @&       )                    �?      �?              @'       (                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @+       f                    @�'�sS�?i            @Z@,       Q                    @�ލL�t�?Q            @T@-       D                    @8�Z$��?4             J@.       ;                    @+	����?             >@/       6                    �?9��8���?             (@0       5                      @B{	�%��?	             "@1       4                     �?؇���X�?             @2       3                    6@z�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �                      @������������������������       �      �?              @7       8                     �?VUUUUU�?             @������������������������       �                     �?9       :                      @      �?              @������������������������       �                     �?������������������������       �                     �?<       A                   �2@��[��"�?             2@=       @                      @���(\��?
             $@>       ?                    �?      �?              @������������������������       �      �?             @������������������������       �      �?             @������������������������       �                      @B       C                    �?      �?              @������������������������       �      �?             @������������������������       �      �?             @E       F                     @�GN�z�?             6@������������������������       �                     @G       P                   �5@�t����?             1@H       O                   �3@      �?             0@I       L                    �?������?             .@J       K                     @�q�q�?	             "@������������������������       �����X�?             @������������������������       �      �?              @M       N                     @r�q��?             @������������������������       �z�G�z�?             @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?R       e                    !@T�<q,��?             =@S       Z                    �? �P|��?             ;@T       U                    @�z�G��?
             $@������������������������       �                     @V       W                    1@      �?             @������������������������       �                     �?X       Y                   �7@���Q��?             @������������������������       �                      @������������������������       ��q�q�?             @[       b                    @���I��?             1@\       a                    <@t�E]t�?             &@]       `                     �?p=
ףp�?
             $@^       _                    @�$I�$I�?             @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?c       d                    4@�8��8��?             @������������������������       �      �?             @������������������������       �                      @������������������������       �                      @g       l                     �?9��8���?             8@h       k                    9@{�G�z�?             @i       j                   �4@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @m       x                    7@�W�3��?             3@n       o                   �2@N贁N�?             .@������������������������       �                     �?p       s                   �4@�m۶m��?             ,@q       r                    �?�q�q�?             @������������������������       �                     �?������������������������       ����Q��?             @t       u                    @      �?              @������������������������       �                     @v       w                    �?z�G�z�?             @������������������������       �                     �?������������������������       �      �?             @y       z                    9@      �?             @������������������������       �                     �?{       |                    <@�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�b�values�hhK ��h��R�(KK}KK��hV�B�2        �?      ,@      7@       @      @      @      @      J@      "@      <@      @      �?      �?      �?       @               @      @      @               @      @      *@      @              �?      �?      @              �?                               @              (@      �?              �?              @                                                              �?                      �?                                                                              �?                      �?                                                                                                      �?                                                                              �?                                      @                                                                                              �?       @              �?                               @              &@      �?                              �?                                               @              "@                                                                                       @              @                                      �?                                                              @                                                                                                      @                                      �?                                                               @                                      �?                                                                                                                                                                       @                              �?      �?              �?                                               @      �?                      �?      �?                                                                      �?                              �?                                                                      �?                                                                                                      �?                              �?                                                                                              �?                                                                                                                              �?                                               @                                                      �?                                              �?                                                                                                      �?                                      �?              �?      @      @                      @      �?      @                              �?                      @                              @              @                              �?                      @                              @                                                                      @                               @                                                                      @                                                                                                                                       @                                              �?                                                      @                                              �?                                                      �?                                                                                                      �?                                              �?                                                                                                                                                              @                                                                                                                      @                                              �?              @                              �?                                                      �?                                              �?                                                      �?                                                                                                                                                      �?                                                                      @                                                                      @      7@                      �?      @      I@       @      .@      �?      �?                      @      (@                              @     �F@              (@      �?      �?                      @       @                              �?     �@@              "@              �?                      @       @                              �?      0@              @              �?                              �?                              �?       @              �?              �?                              �?                                      @              �?                                              �?                                      @                                                              �?                                      @                                                              �?                                       @                                                                                                       @                                                                                                       @                                                                                                      �?              �?                                                                              �?      �?                              �?                                                              �?                                                                                                              �?                              �?                                                                                                      �?                                                                      �?                                                      @      �?                                       @              @                                       @      �?                                      @              �?                                       @      �?                                      @              �?                                      �?                                               @              �?                                      �?      �?                                       @                                                                                                       @                                                      @                                               @               @                                       @                                               @                                                       @                                                               @                                                                                      1@              @                                                                                      @                                                                                                      (@              @                                                                                      (@              @                                                                                      &@              @                                                                                      @              @                                                                                      @               @                                                                                      �?              �?                                                                                      @              �?                                                                                      @              �?                                                                                      �?                                                                                                      �?                                                                                                                      �?                                              $@                              @      (@              @      �?                                      $@                              �?      (@              @      �?                                      @                                      @                                                              @                                                                                                      @                                      @                                                              �?                                                                                                       @                                      @                                                                                                       @                                                               @                                      �?                                                              @                              �?      "@              @      �?                                       @                              �?      @                      �?                                       @                              �?      @                                                               @                              �?      @                                                               @                                      @                                                                                              �?                                                                                                              @                                                                                                                              �?                                      �?                                       @              @                                              �?                                                      @                                                                                       @                                                                                               @                                                                      &@                      �?       @      @       @      @                                                                               @      �?       @                                                                                       @      �?                                                                                                      �?                                                                                               @                                                                                                                       @                                                      &@                      �?              @              @                                              &@                                       @               @                                                                                                      �?                                              &@                                       @              �?                                              @                                       @                                                              �?                                                                                                      @                                       @                                                              @                                                      �?                                              @                                                                                                      @                                                      �?                                              �?                                                                                                      @                                                      �?                                                                      �?               @              �?                                                                                                      �?                                                                      �?               @                                                                                                       @                                                                                      �?                                                        �t�bub�_sklearn_version��1.1.0�ub.