���"      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K
�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK	��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�CH                                                         	       �t�b�
n_classes_�h�scalar���h%C	       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C	       �t�bK��R�}�(h	K�
node_count�K=�nodes�hhK ��h��R�(KK=��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�BX                               @�����V@s            �\@                            �?����@Q            @T@                           �?���W��?             3@                           @�1H����?              @������������������������       �      �?              @������������������������       �                     @������������������������       �                     &@                           �?P�k��@>             O@	                           @�������?"             A@
                          �4@���'���?             @������������������������       �                     @������������������������       �                     @                          �1@* ����?             ;@                            �?z&F�Y�?             @������������������������       �|%��b�?             @������������������������       �                      @                          �4@.a�� �?             6@������������������������       �                     3@                          �5@|%��b�?             @������������������������       �                      @������������������������       �                     �?                          �0@�l���?             <@������������������������       �                     @                           �?�ݎ���?             6@                           @b#���?             .@                           @�9>����?             ,@������������������������       �|%��b�?             @������������������������       �                      @������������������������       �                     �?                           @�9>����?             @������������������������       �                     @������������������������       �                     �?!       (                    �?��-� @"             A@"       '                    4@_�z|�X�?             @#       $                    �?�c�����?             @������������������������       �                      @%       &                   �1@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @)       :                   �4@���W�e�?             <@*       3                    @p��I�?             8@+       2                    �?�TS�~�?             *@,       -                   �1@��&��?
             $@������������������������       �                     �?.       1                    �?|%��b�?	             "@/       0                    3@�Z���?             @������������������������       ��c�����?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     @4       7                    �?bo-���?             &@5       6                    3@|%��b�?             @������������������������       �                     �?������������������������       �                      @8       9                   �3@�c�����?              @������������������������       �                     @������������������������       �      �?             @;       <                     @      �?             @������������������������       �                      @������������������������       �                      @�t�b�values�hhK ��h��R�(KK=KK	��hV�B(        9@      @      @      @      0@      @      (@      3@      5@      (@      @      �?      @      ,@              �?      3@      5@                      �?      @                      �?      &@                              �?      @                      �?                                      �?                              �?                                              @                                                                                                      &@              (@      @                      ,@                       @      5@      @      @                      �?                       @      4@      @      @                                                              @                                                                              @                                                                      @                      �?                       @      4@               @                      �?                       @                       @                      �?                                                                                               @                       @                                                      4@                                                                      3@               @                                                      �?               @                                                                                                                              �?       @                              *@                      @      �?                                                              @               @                              *@                              �?       @                              (@                              �?       @                              (@                                       @                              @                                                                       @                                                                                                      �?      @                              �?                                      @                                                                                                      �?                                      *@               @      �?       @      @      &@                                       @      �?              @                                                      �?              @                                                                       @                                                      �?              �?                                                                      �?                                                      �?                                                               @                                                      *@                               @       @      &@                      &@                                       @      &@                      @                                              "@                      @                                              @                      �?                                                                      @                                              @                      �?                                              @                      �?                                              @                                                                      �?                       @                                               @                                                                      @                      @                                       @       @                      �?                                       @                              �?                                                                                                               @                              @                                               @                      @                                                                       @                                               @                       @                               @                                       @                                                                                                       @                                �t�bub�_sklearn_version��1.1.0�ub.