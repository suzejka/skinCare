��u.      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C`                                                                	       
              �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K�
node_count�KG�nodes�hhK ��h��R�(KKG��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B�         *                   �5@�큺s@�             c@                           @vD,͒�@g            �Y@                            @�����@X             V@                          �4@���J�l@:             M@                            �?ݾ�*y_�?1            �H@                           3@��Tx�?$             B@������������������������       ���Y���?             6@������������������������       �J��MY.�?             ,@	       
                    �?׻����?             *@������������������������       ��c�����?             @������������������������       �M�)9��?	             "@                           �?hJN�@	             "@                           @z&F�Y�?             @������������������������       �|%��b�?             @������������������������       �                      @                            �?      �?             @������������������������       �                      @������������������������       �      �?              @                           �?��XF��?             >@                          �1@hJN��?             @������������������������       �                     �?                           4@�Z���?             @������������������������       �                     @������������������������       �      �?              @                           @6� 7�?             8@                            @M�)9��?             2@������������������������       ��c�����?             @������������������������       ����;E��?             ,@                           �?V�T����?             @������������������������       �                     @������������������������       �      �?              @        !                     �?�{���?             .@������������������������       �                     �?"       %                    �?�X�Ą�?             ,@#       $                    @      �?              @������������������������       �                     �?������������������������       �                     �?&       '                   �2@�c�����?             (@������������������������       �                     �?(       )                     �?r�Mh�?             &@������������������������       �|%��b�?             @������������������������       ��Z���?             @+       4                    �?� æ���?2             I@,       1                    @�,�4�?             @-       0                    �?z&F�Y�?             @.       /                     �?      �?             @������������������������       �      �?              @������������������������       �      �?              @������������������������       �                     �?2       3                    �?      �?              @������������������������       �                     �?������������������������       �                     �?5       >                   �6@��� O�?+            �E@6       =                    @^�z|�X�?             (@7       :                     @q-�"�?
             $@8       9                    �?�c�����?              @������������������������       �                     @������������������������       �      �?             @;       <                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @?       F                   �8@��OD�P�?             ?@@       C                     �?p�h8/�?             1@A       B                    �?       @             @������������������������       �      �?              @������������������������       �      �?              @D       E                    @�%�`I��?             *@������������������������       �                      @������������������������       �>���i��?             @������������������������       �                     ,@�t�b�values�hhK ��h��R�(KKGKK��hV�B�        "@      �?       @      �?      :@       @      �?     �C@      @@      :@       @      (@      @                              6@       @      �?      @      ?@      8@              &@      @                              3@       @      �?      @      ?@      8@              �?      @                              *@       @      �?       @      "@      8@              �?      @                              (@                              "@      6@                      @                              $@                              "@      &@                                                      @                              @      &@                      @                              @                               @                                                               @                                      &@                                                      �?                                      @                                                      �?                                       @                                                      �?       @      �?       @               @              �?                                      �?       @               @                                                                      �?                       @                                                                               @                                                                                                      �?                       @              �?                                                                               @                                                                      �?                                      �?      �?                              @                      �?      6@                              �?                              @                              �?                                                                                              �?                              �?                              @                                                                                              @                                                              �?                              �?                                                                                               @                      �?      5@                                                               @                              0@                                                              �?                              @                                                              �?                              *@                                                                                      �?      @                                                                                              @                                                                                      �?      �?                                                              @                       @                              $@                                                              �?                                                                      @                      �?                              $@                                                              �?                              �?                                                              �?                                                                                                                              �?                                      @                                                      "@                                                                                              �?                                      @                                                       @                                       @                                                      @                                      �?                                                      @       @      �?       @      �?      @                      A@      �?       @       @      �?       @                               @                       @                              �?       @                               @                      �?                                       @                              �?                      �?                                      �?                              �?                                                              �?                                                      �?                                                                      �?                                                                                                                      �?                              �?                                                              �?                                                                                                                              �?              �?       @      �?       @                      @@      �?       @       @                               @              �?                      @      �?               @                               @              �?                      @      �?                                               @                                      @                                                                                              @                                                       @                                       @                                                                      �?                              �?                                                                                              �?                                                              �?                                                                                                                                               @                      �?              �?      �?                      :@               @                              �?              �?      �?                      (@               @                              �?              �?                              �?              �?                                                                              �?              �?                              �?              �?                                                                                                      �?                      &@              �?                                                                               @                                                                      �?                      @              �?                                                                              ,@                                �t�bub�_sklearn_version��1.1.0�ub.