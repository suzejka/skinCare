���J      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C`                                                         	       
                     �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K
�
node_count�Kw�nodes�hhK ��h��R�(KKw��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B         >                     �?W�XYv�?�             c@       +                   �5@M n�r�?K            �R@                           �?������?4             J@������������������������       �r�q��?             @       *                    !@Fp�u=q�?.             G@                            �?���|���?,             F@                           �?Er���&�?             1@������������������������       �                     @	                           @��X��?             ,@
                           �?pƵHP�?             *@                           �?      �?             @                           3@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?                           @x�5?,�?	             "@                           3@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       ��8��8��?             @������������������������       �                     �?       #                    �?�dIG���?             ;@       "                   �4@����[��?             2@                           �?     @�?             0@                           @      �?              @������������������������       �                     �?                          �1@������?             @������������������������       �      �?             @������������������������       �VUUUUU�?             @       !                    @      �?              @                            @����X�?             @������������������������       �      �?             @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                      @$       )                    @|	�%���?	             "@%       (                    @      �?              @&       '                    @      �?             @������������������������       �                      @������������������������       �      �?              @������������������������       �      �?             @������������������������       �                     �?������������������������       �                      @,       =                    A@\X��t�?             7@-       2                    �?b>���?             5@.       /                   �7@�8��8��?             (@������������������������       �                     @0       1                   �8@z�G�z�?             @������������������������       �                     �?������������������������       �                     @3       6                    7@h/�����?	             "@4       5                     �?�q�q�?             @������������������������       �                      @������������������������       �                     �?7       <                    @�q�q�?             @8       9                    �?z�G�z�?             @������������������������       �                      @:       ;                    :@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @?       v                   �8@>���>�?N            �S@@       O                    �?�"e����?H             R@A       N                    7@J�w�"w�?             3@B       K                   �3@�θ�?             *@C       H                    �?:/����?             @D       G                    �?      �?             @E       F                   �1@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?I       J                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?L       M                   �5@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @P       e                     @��h�7�?5            �J@Q       \                   �4@<�.����?             ?@R       U                    @>
ףp=�?             4@S       T                    �?      �?              @������������������������       �      �?             @������������������������       �                     @V       W                    �?      �?             (@������������������������       �                      @X       [                   �2@�z�G��?
             $@Y       Z                   �0@z�G�z�?             @������������������������       �      �?             @������������������������       �                     �?������������������������       ����Q��?             @]       `                    @*L�9��?             &@^       _                    �?�Q����?             @������������������������       �VUUUUU�?             @������������������������       �                      @a       d                     @      �?             @b       c                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @f       k                    �?�ˠT��?             6@g       h                    @�X�C�?             ,@������������������������       �                      @i       j                    �?��8��8�?             (@������������������������       �����X�?             @������������������������       �{�G�z�?             @l       o                    @      �?              @m       n                    @VUUUUU�?             @������������������������       �                     �?������������������������       �      �?              @p       s                   �3@�Q����?             @q       r                    �?�q�q�?             @������������������������       �      �?              @������������������������       �                     �?t       u                   �5@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�t�b�values�hhK ��h��R�(KKwKK��hV�B�,         @      @      :@      6@      *@      �?      0@       @       @       @      2@      G@       @      �?       @      $@       @      �?      @       @       @               @      C@                       @      $@              �?      @       @                       @      6@                              �?                                                      @                               @      "@              �?      @       @                      @      6@                       @      "@              �?      @                              @      6@                              @                      @                                      @                                                                                              @                              @                      @                                      @                              @                      @                                      @                                                       @                                       @                                                       @                                      �?                                                       @                                                                                                                                      �?                                                                                              �?                              @                      @                                      �?                              �?                       @                                                                                              �?                                                                      �?                      �?                                                                       @                      @                                      �?                                                                                              �?                       @      @              �?                                      @      .@                      �?      @                                                       @      "@                      �?      @                                                       @      "@                      �?       @                                                       @      @                                                                                              �?                      �?       @                                                       @       @                      �?      �?                                                      �?      �?                              �?                                                      �?      �?                               @                                                              @                               @                                                              @                              �?                                                              @                              �?                                                               @                                                                                              �?                               @                                                                                      �?                      �?                                      �?      @                      �?                                                              �?      @                                                                                      �?      @                                                                                               @                                                                                      �?      �?                      �?                                                                      @                                              �?                                                                                                               @                                       @      �?                       @                               @                      0@       @      �?                                                       @                      0@              �?                                                                              &@                                                                                              @              �?                                                                              @              �?                                                                                                                                                                              @       @                                                               @                      @       @                                                                                      �?       @                                                                                                                                                                                      �?                                                                       @                      @                                                                      �?                      @                                                                                               @                                                                      �?                       @                                                                      �?                                                                                                                       @                                                                      �?                                                               @                                                                       @      8@      (@      &@              "@                       @      $@       @               @      8@      (@      @              "@                       @      $@       @               @              @                                               @      @      @               @              @                                               @      @                       @              @                                               @                                               @                                               @                                              �?                                               @                                              �?                                                                                                                                               @                                              �?                                                                               @              �?                                                                               @                                                                                                              �?                                                                                               @                                                      @                                                                                              @                                       @                                                                                                                                                              @                      8@      @      @              "@                              @       @                      2@      @      @               @                              @      �?                      .@      �?                      �?                              @                              @      �?                      �?                                                               @      �?                      �?                                                              @                                                                                              "@                                                              @                               @                                                                                              @                                                              @                              @                                                              �?                              @                                                              �?                              �?                                                                                              @                                                               @                              @       @      @              �?                                      �?                      @      �?                                                              �?                      �?      �?                                                              �?                       @                                                                                                      �?      @              �?                                                                      �?                      �?                                                                      �?                                                                                                                      �?                                                                              @                                                                              @      @      �?              @                              @      �?                      @       @                      @                                                               @                                                                                              @       @                      @                                                               @                              @                                                              �?       @                       @                                                              �?       @      �?                                              @      �?                              �?      �?                                                      �?                                      �?                                                                                      �?                                                              �?                      �?      �?                                                      @                              �?                                                               @                              �?                                                              �?                                                                                              �?                                      �?                                                      �?                                      �?                                                                                                                                                      �?                                              @                                                        �t�bub�_sklearn_version��1.1.0�ub.