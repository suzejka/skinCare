���d      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K
�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C�                                                                	       
                                                        �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K
�
node_count�K{�nodes�hhK ��h��R�(KK{��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B�         l                    @�~Q$���?�             c@       S                    @��YEd��?�             `@       H                    @�r���?\             W@       +                   �5@����[�?H             R@                           @g�x�P��?*             E@                           �?�9����?             6@                          �1@�ˠT�?             &@������������������������       �                     �?	                           3@
ףp=
�?
             $@
                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                            �?      �?              @������������������������       ��q�q�?             @                             @
ףp=
�?             @������������������������       �      �?              @������������������������       �VUUUUU�?             @                          �4@b���i��?             &@                           �?��Q��?
             $@                            �?h/�����?	             "@������������������������       ��8��8��?             @                           �?�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                     �?������������������������       �                     �?       &                      @p=
ףp�?             4@       %                    @.k��\�?             1@       "                    @     ��?             0@       !                    �?�q�q�?             @                            3@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     @#       $                    �?ףp=
�?
             $@������������������������       �                     @������������������������       �r�q��?             @������������������������       �                     �?'       *                    �?VUUUUU�?             @(       )                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?,       9                    @[�[��?             >@-       2                    �?��]�`��?             *@.       /                    �?���Q��?             @������������������������       �                     �?0       1                     �?      �?             @������������������������       �      �?              @������������������������       �      �?              @3       4                     @      �?              @������������������������       �                     @5       6                    �?�Q����?             @������������������������       �                     �?7       8                     @      �?             @������������������������       ��q�q�?             @������������������������       �                     �?:       ;                    �?J,�ѳ�?             1@������������������������       �                     @<       ?                   �6@�T�x?r�?             &@=       >                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @@       G                     �?      �?              @A       D                    @�8��8��?             @B       C                    @�q�q�?             @������������������������       �      �?              @������������������������       �                     �?E       F                    <@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �      �?              @I       R                   �4@��(\���?             4@J       Q                     @�����H�?             2@K       N                   �2@      �?             0@L       M                    �?      �?              @������������������������       �                     @������������������������       �      �?             @O       P                    �?      �?              @������������������������       �      �?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @T       c                     @���z�?%            �B@U       X                     �?ffffff�?             4@V       W                    @      �?             @������������������������       ��q�q�?             @������������������������       �                     �?Y       \                   �7@     @�?             0@Z       [                    �?      �?              @������������������������       �                     @������������������������       �      �?             @]       b                    @      �?              @^       a                    <@�8��8��?             @_       `                    �?���Q��?             @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @d       i                   �3@�"�O�|�?             1@e       h                    �?��S�ۿ?             .@f       g                     @�����H�?	             "@������������������������       �؇���X�?             @������������������������       �                      @������������������������       �                     @j       k                   �5@      �?              @������������������������       �                     �?������������������������       �                     �?m       n                     �?��8��8�?             8@������������������������       �                     @o       z                    @��uJ���?             3@p       q                    �?     ��?             0@������������������������       �                     @r       u                     �?�θ�?             *@s       t                    @�q�q�?             @������������������������       �      �?              @������������������������       �      �?             @v       w                   �2@؇���X�?             @������������������������       �                     �?x       y                    6@r�q��?             @������������������������       �z�G�z�?             @������������������������       �                     �?������������������������       �                     @�t�b�values�hhK ��h��R�(KK{KK��hV�B0E        0@      @      �?      ,@      �?      9@      "@       @      5@      �?      �?      @      $@      @      .@      @      2@      �?      0@      @      �?      ,@      �?      6@      "@       @      5@      �?      �?      @      $@      @       @      @      *@      �?       @      @              ,@      �?      .@      @       @      5@      �?      �?      @      �?      @       @       @      (@      �?       @      @              ,@      �?      *@      @       @      @      �?      �?      @      �?      @       @       @      $@      �?       @                      ,@              $@      @              @              �?              �?       @       @              �?              �?                      �?              @      @              @                                       @       @              �?              �?                                      @      @                                                      �?      �?              �?                                                                                                                      �?                                      �?                                      @      @                                                              �?              �?                                                              �?                                                                              �?                                                              �?                                                                                                                                                                                                                              �?              �?                                      @      @                                                              �?                                                                      �?       @                                                                                              �?                                       @      �?                                                              �?                                                                      �?                                                                      �?                              �?                                      �?      �?                                                                                                                      �?              @                      @                                      �?      �?                                                      �?              @                      @                                      �?                                                                              @                      @                                      �?                                                                               @                      @                                      �?                                                                               @                      �?                                                                                                                      �?                                                                                                                                              �?                      �?                                                                                                      �?                                                                                                                                                                                                                                      �?                              �?                      *@              @                      �?              �?              �?                                                                      *@              @                                      �?                                                                                      *@              @                                                                                                                              @               @                                                                                                                              �?               @                                                                                                                              �?              �?                                                                                                                                              �?                                                                                                                              @                                                                                                                                              "@              �?                                                                                                                              @                                                                                                                                              @              �?                                                                                                                                                                                      �?                                                              �?                                                              �?                              �?                                              �?                                                              �?                                                                                                                                              �?                                                                              �?                                                                                                                                                                                                                                              �?                                                      @                      �?      @       @       @              �?              @              �?               @      "@      �?              @                              @       @                                      @              �?              �?                                                              @       @                                                                                                                                      �?                                                                                                                                               @       @                                                                                                                                      �?      �?                                                                                                                                      �?      �?                                                                                                      @                                                                              @              �?              �?                              @                                                                                                                                                                                                                              @              �?              �?                                                                                                                              �?                                                                                                                              @                              �?                                                                                                               @                              �?                                                                                                              �?                                                               @                      �?                       @              �?                                              �?      "@      �?                                                                                                                                      @                       @                      �?                       @              �?                                              �?      @      �?                                                               @              �?                                                                                                                                              �?                                                                                                                               @                                                                                               @                      �?                                                                                      �?      @      �?               @                      �?                                                                                              @                                              �?                                                                                               @                                              �?                                                                                              �?                                                                                                                                              �?                       @                                                                                                                      �?                      �?                                                                                                                                              �?                                                                                                                      �?                                                                                                                                      �?              �?                                               @                      0@                                                               @                                                       @                      0@                                                                                                                       @                      ,@                                                                                                                      �?                      @                                                                                                                                              @                                                                                                                      �?                      @                                                                                                                      �?                      @                                                                                                                      �?                      @                                                                                                                                              @                                                                                                                                               @                                                                                                                                                                                                               @              ,@              �?                      @      @                                              "@                       @      �?                                                      @      @                                              "@                       @      �?                                                      �?      @                                                                                                                                      �?       @                                                                                                                                              �?                                                                                                                                      @                                                      "@                       @      �?                                                      �?                                                      @                                                                                                                                              @                                                                                      �?                                                      @                                                                                      @                                                       @                       @      �?                                                      @                                                       @                              �?                                                      @                                                       @                                                                                      �?                                                       @                                                                                       @                                                                                                                                                                                                                                      �?                                                                                                                                       @                      ,@              �?                       @                                                                                                      ,@                                      �?                                                                                                       @                                      �?                                                                                                      @                                      �?                                                                                                       @                                                                                                                                              @                                                                                                                                                              �?                      �?                                                                                                                      �?                                                                                                                                                                      �?                                                                                                                                              @                                                                      *@      @      @                                                                                                                                              @                                                      @                                                                      *@      @                                                              @                                                                      *@                                                                                                                                              @                                                                      @                                                                      $@                                                                       @                                                                      @                                                                      �?                                                                      �?                                                                      �?                                                                      @                                                                      �?                                                                      @                                                                                                                                              �?                                                                      �?                                                                      @                                                                      �?                                                                      @                                                                                                                                              �?                                                                                                                                                      @                �t�bub�_sklearn_version��1.1.0�ub.