��e1      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK
��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�CP                                                                	       �t�b�
n_classes_�h�scalar���h%C
       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C
       �t�bK��R�}�(h	K�
node_count�KU�nodes�hhK ��h��R�(KKU��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B�         @                    @[ZM�@s            �\@       !                     @&�����@S            �T@                           �?]���f@1            �H@                            �? ۉ����?             &@                           �?��'4���?              @������������������������       �      �?              @                           �?|%��b�?             @������������������������       �                     @	       
                    3@|%��b�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                     @                          �2@��q�u�?&             C@                           @���G�?             ,@                           �?M�)9��?	             "@������������������������       �                     @������������������������       �V�T����?             @                           �?�Z���?             @������������������������       �                      @������������������������       �|%��b�?             @                            �?�+���7�?             8@                           6@V�T����?             @������������������������       �|%��b�?             @������������������������       �                     @                            �?V�T����?             2@                           �?�c�����?              @                           @V�T����?             @������������������������       �                      @������������������������       ��c�����?             @������������������������       �      �?              @                            �?���?
             $@������������������������       �V�T����?             @������������������������       �                     @"       3                   �2@׮m@"             A@#       $                    �?���dK��?             3@������������������������       �                     @%       ,                    �?n>�v�9�?             0@&       '                    �?���?
             $@������������������������       �                     @(       +                    �?V�T����?             @)       *                   �1@�Z���?             @������������������������       �                     �?������������������������       ��c�����?             @������������������������       �                     �?-       .                    @_�z|�X�?             @������������������������       �      �?              @/       0                    @�c�����?             @������������������������       �                      @1       2                    �?      �?              @������������������������       �                     �?������������������������       �                     �?4       =                    @�)T��@             .@5       :                   �4@4�q��?             (@6       7                     @��b}�?              @������������������������       �                      @8       9                    �?^�z|�X�?             @������������������������       �      �?              @������������������������       �      �?             @;       <                    �?      �?             @������������������������       �      �?              @������������������������       �      �?              @>       ?                   �5@|%��b�?             @������������������������       �                      @������������������������       �                     �?A       J                    @WA�M�} @              @@B       E                    �?��F���?             2@C       D                    @M�)9��?	             "@������������������������       ��Z���?             @������������������������       �                     @F       G                   �2@�t�I�|�?	             "@������������������������       �                     �?H       I                     �?��b}�?              @������������������������       �      �?              @������������������������       �|%��b�?             @K       T                    @�bN�� @             ,@L       O                    1@4S����?             &@M       N                    �?V�T����?             @������������������������       �                      @������������������������       ��c�����?             @P       S                    �?z&F�Y�?             @Q       R                    @|%��b�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�t�b�values�hhK ��h��R�(KKUKK
��hV�B�         @      5@      4@       @      "@      @      5@      3@      @      @      @      0@      4@              "@              @      3@      @      @      @       @      4@               @              @      @                      @       @      �?                                      @                               @      �?                                      @                                      �?                                      �?                               @                                              @                                                                              @                               @                                              �?                              �?                                                                              �?                                              �?                      @                                                                                      @      3@               @              @                                       @      @               @                                                      �?                       @                                                                              @                                                      �?                      @                                                      �?      @                                                                               @                                                                      �?       @                                                                      @      .@                              @                                      �?                                      @                                      �?                                       @                                                                              @                                      @      .@                                                                       @      @                                                                      �?      @                                                                               @                                                                      �?      @                                                                      �?      �?                                                                      �?      "@                                                                      �?      @                                                                              @                                                                       @                      �?               @      ,@      @      @              @                      �?                      (@      @                                                                              @                      @                      �?                      (@                              �?                                              "@                                                                              @                              �?                                              @                              �?                                              @                                                                              �?                              �?                                              @                                                                              �?                               @                      �?                      @                              �?                      �?                                                      �?                                              @                                                                               @                              �?                                              �?                                                                              �?                              �?                                                                              @                                       @       @       @      @              @                                       @      �?              @              @                                              �?              @                                                                               @              @                                              �?               @              �?                                                              �?               @                                              �?              �?               @                                       @                                      �?                                      �?                                      �?                                      �?                                                                                      �?       @                                                                               @                                                                      �?                      @      @               @              @      ,@                               @      @                                      (@                                      �?                                       @                                      �?                                      @                                                                              @                               @      @                                      @                              �?                                                                              �?      @                                      @                              �?      �?                                                                               @                                      @                              @      �?               @              @       @                                      �?               @              @       @                                      �?                              @                                                                               @                                              �?                              @                                                               @              �?       @                                                                      �?       @                                                                      �?      �?                                                                              �?                                                       @                                                      @                                                                        �t�bub�_sklearn_version��1.1.0�ub.