��2K      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K
�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C�                                                                	       
                                                               �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K
�
node_count�KW�nodes�hhK ��h��R�(KKW��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B         &                    �?�(W��?�             e@                            �?>z��.�?D             Q@                           >@r�q��?             8@                          �5@>F?�!��?             5@������������������������       �                     &@                           �?ףp=
��?
             $@������������������������       �                     @       	                   �6@�8��8��?             @������������������������       �                      @
                          �7@      �?             @������������������������       �                     @������������������������       �                     �?                          �@@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           7@}��7�?,             F@                           @�
t�F��?             1@                             @9��8���?             (@������������������������       �                     @                           �?��"e���?	             "@                          �5@�8��8��?             @                           �?���Q��?             @������������������������       �                      @                           3@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     @       %                     @�+$�jP�?             ;@       "                    �?F]t�E�?             &@        !                    �?���Q��?             @������������������������       �                     @������������������������       �                      @#       $                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     0@'       .                    @I.�!���?d             Y@(       -                    @�x?r���?             6@)       *                      @���N8�?             5@������������������������       �                     2@+       ,                     @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?/       H                    @|1z�?�?N            �S@0       E                     @��Y��?5            �J@1       2                    @*D>��?'            �C@������������������������       �                     2@3       D                    !@4և����?             5@4       =                    �?Dy�5��?             3@5       8                    @      �?              @6       7                   �5@      �?              @������������������������       �                     �?������������������������       �                     �?9       <                    @r�q��?             @:       ;                   �3@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @>       ?                   �1@}��7�?             &@������������������������       �      �?             @@       A                    6@�$I�$I�?             @������������������������       �                      @B       C                    ;@{�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �                      @F       G                     @����X�?             ,@������������������������       �        
             $@������������������������       �                     @I       N                    8@.n���?             9@J       M                     �?0�����?             2@K       L                   �4@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     0@O       P                    @������?             @������������������������       �                     @Q       R                   �:@      �?             @������������������������       �                     �?S       T                   �;@VUUUUU�?             @������������������������       �                     �?U       V                   �<@      �?              @������������������������       �                     �?������������������������       �                     �?�t�b�values�hhK ��h��R�(KKWKK��hV�B�3        3@      @      .@      �?      @      �?      @      =@      9@      @      @      @      4@      0@       @      @      @      @      @      @      @      @              @      �?      @                       @      @      @      2@      0@              @                      @                                              �?                               @      @       @      0@                                                                                                                               @      @              0@                                                                                                                                                      &@                                                                                                                               @      @              @                                                                                                                                                      @                                                                                                                               @      @              �?                                                                                                                               @                                                                                                                                                              @              �?                                                                                                                                      @                                                                                                                                                                      �?                                                                                              �?                                               @                                                                                                      �?                                                                                                                                                                                                       @                                                              @      @      @              @              @                                       @       @      0@              @                      @      @              @              @                                                               @                      @                      �?      @                              @                                                               @                      @                      �?      @                                                                                                                                                                                      @                                                               @                      @                      �?                                                                                                       @                      @                      �?                                                                                                       @                      @                                                                                                                                                       @                                                                                                                               @                      �?                                                                                                                              �?                                                                                                                                                      �?                      �?                                                                                                                                                                              �?                                      @                                                                                                                                      @                                                                                                                                              @                                      @                                       @              0@                                       @              @                                      @                                       @                                                       @              @                                                                                                                                       @              @                                                                                                                                                                                                                                                                                               @                                                      @                                       @                                                                                                              @                                                                                                                                                                                               @                                                                                                                                                                      0@                                              0@      �?      $@      �?                              =@      9@       @      �?       @       @               @              @      @                      �?                                                      4@              �?                                                                              �?                                                      4@                                                                                                                                                      2@                                                                                              �?                                                       @                                                                                                                                                       @                                                                                              �?                                                                                                                                                                                                                              �?                                                                      0@              $@      �?                              =@      @       @               @       @               @              @      @                              $@                                      =@      @       @              �?                       @                      @                                                                      9@      @       @              �?                       @                      @                                                                      2@                                                                                                                                                      @      @       @              �?                       @                      @                                                                      @      @                      �?                       @                      @                                                                      @                              �?                      �?                      �?                                                                                                      �?                      �?                                                                                                                              �?                                                                                                                                                                              �?                                                                                              @                                                                              �?                                                                      �?                                                                              �?                                                                      �?                                                                                                                                                                                                                                      �?                                                                      @                                                                                                                                                       @      @                                              �?                      @                                                                       @       @                                                                                                                                                       @                                              �?                      @                                                                                                                                                       @                                                                               @                                              �?                       @                                                                               @                                              �?                                                                                                                                                                               @                                                                                       @                                                                                              $@                                      @                                                                                                              $@                                                                                                                                                                                              @                                                                                              0@                      �?                                      �?                      �?       @                              @      �?              0@                      �?                                                                      �?                                                                              �?                                                                      �?                                                                                                                                                      �?                                                                              �?                                                                                                                              0@                                                                                                                                                                                                                      �?                      �?      �?                              @      �?                                                                                                                                              @                                                                                      �?                      �?      �?                                      �?                                                                                                      �?                                                                                                                              �?                              �?                                      �?                                                                                                              �?                                                                                                                      �?                                                                      �?                                                                              �?                                                                                                                                                                                                                              �?        �t�bub�_sklearn_version��1.1.0�ub.