���3      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK
��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�CP                                                                	       �t�b�
n_classes_�h�scalar���h%C
       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C
       �t�bK��R�}�(h	K
�
node_count�KY�nodes�hhK ��h��R�(KKY��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�Bx         (                    �?���@�             c@                          �7@2�xx�S@0             H@                           @�&,�@�@"             A@                           �?K���?             :@                            �?	o���8�?             ,@������������������������       �                     @                           4@��'4���?              @       	                    �?�c�����?             @������������������������       �                      @
                          �1@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?      �?             @                          �5@|%��b�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     �?                             @η:�?             (@������������������������       �                      @                           �?�c�����?             @������������������������       �                     �?                           �?|%��b�?             @������������������������       �      �?              @������������������������       �                     �?                           �?      �?              @������������������������       �                     @                           �?      �?             @������������������������       �                     �?                          �6@|%��b�?             @������������������������       �                      @������������������������       �                     �?        '                    >@5�ڣX�?             ,@!       &                     �?��Yo��?
             $@"       #                    �?      �?             @������������������������       �                      @$       %                   �8@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @)       L                   �7@A����m @i            @Z@*       ?                     @�:
K�D�?U            @U@+       >                     �?o�gv��?A            @P@,       9                    @2ߗ2�$�?)            �D@-       0                     �?�\`���?             6@.       /                    �?      �?             @������������������������       �                     @������������������������       �                     @1       8                    @>s_X��?             0@2       7                    �?��0r��?             &@3       6                   �2@�Q$��?	             "@4       5                    �?      �?              @������������������������       ��c�����?             @������������������������       ��c�����?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @:       ;                    @cB���?             3@������������������������       �                     .@<       =                    !@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     8@@       C                    @x��s�?             4@A       B                    @|%��b�?             @������������������������       �                     �?������������������������       �                      @D       E                     @W�oθ�?             1@������������������������       �                     (@F       K                   �5@��&��?             @G       J                   �3@�c�����?             @H       I                    �?|%��b�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?M       V                   �8@Pu�x�{@             4@N       Q                    @��h/%^�?             *@O       P                    �?|%��b�?             @������������������������       �                     @������������������������       �                      @R       S                    �?������?             @������������������������       �                     @T       U                    @      �?             @������������������������       �                      @������������������������       �                      @W       X                    @������?             @������������������������       �                      @������������������������       �                     @�t�b�values�hhK ��h��R�(KKYKK
��hV�B�        *@      H@      ;@       @      "@      $@      @     �@@       @      @      &@              ,@       @      @       @      @       @              @      $@              *@       @                      @       @              @      "@              *@                              @      �?                       @              @                                      �?                      @                                                                               @              @                                      �?                                      @                                      �?                                       @                                                                              �?                                      �?                                      �?                                                                                                                      �?                       @               @                                                               @              �?                                                              �?              �?                                                              �?                                                                                              �?                                                              �?               @                              @                                               @                                                              �?                                              @                                                                              �?                              �?                                               @                              �?                                              �?                                                                              �?                              �?                       @                              �?              @                                                                              @      �?                       @                              �?                      �?                                                                                                       @                              �?                                               @                                                                                                              �?                      �?              �?              @       @                                      �?              �?                       @                                      �?              �?                       @                                                                               @                                      �?              �?                                                              �?                                                                                              �?                                                                                                      @                                                                      @                                               @      H@      *@              @       @              ?@       @       @       @     �E@      @                                      ?@               @              E@      @                                      0@               @              2@      @                                      0@               @              @      @                                      ,@                              @                                              @                              @                                                                                                                              @                                      @                                      &@                                      @                                      @                                      @                                      @                                      @                                      @                                      �?                                      @                                      @                                      �?                                      �?                                                                                                                       @                                                                              @                              .@                                               @               @              .@                                                                                                                               @               @                                                               @                                                                                               @              8@                                                                       @      �?       @                                      .@                       @      �?                                                                              �?                                                                       @                                                                                               @                                      .@                                                                              (@                                       @                                      @                                      �?                                      @                                      �?                                       @                                      �?                                      �?                                                                              �?                                                                              �?                                      �?                                                                      @      @              @       @                       @                      @      @                                               @                              @                                               @                              @                                                                                                                               @                      @       @                                                                      @                                                                               @       @                                                                       @                                                                                       @                                                                                              @       @                                                                               @                                                                      @                                        �t�bub�_sklearn_version��1.1.0�ub.