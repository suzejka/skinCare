���      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C@                                                         �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K�
node_count�K�nodes�hhK ��h��R�(KK��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B�                             @�`��@s            �\@                           �?���@0             H@                           �?T'�Ȭ@             ;@                             @n���?             @������������������������       �                     @                           �?      �?             @������������������������       �                      @������������������������       �                      @	       
                     �?>pF�`�?             4@������������������������       �                      @                           �?���V��?             (@                          �3@      �?             @                          �1@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �?              @������������������������       �                      @������������������������       �                     5@                           @��'�lm�?C            �P@                            @�;[R/��?3            �I@                           @1@� h�?#            �A@������������������������       �                     8@                           �?"S,f�B�?             &@������������������������       �                     @                           4@|%��b�?             @������������������������       �      �?             @������������������������       �                      @                           �?���l��?             0@������������������������       �        	             "@������������������������       �                     @������������������������       �                     0@�t�b�values�hhK ��h��R�(KKKK��hV�B�        3@      1@       @      C@      9@      �?      $@      @      @       @       @              5@      �?      $@      @      @       @       @                      �?      $@      @      @               @                                       @      @                                                                               @                                       @                                                               @                       @                                                       @                              �?      $@      �?                                                       @                       @                              �?       @      �?                                              �?       @      �?                                              �?      �?                                                              �?                                                      �?                                                                      �?      �?               @                                                                                      5@                              0@      "@              C@      @                                      "@              C@      @                                                      ?@      @                                                      8@                                                              @      @                                                      @                                                               @      @                                                       @       @                                                               @                                      "@              @                                              "@                                                                              @                                      0@                                                        �t�bub�_sklearn_version��1.1.0�ub.