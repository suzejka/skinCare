���      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C�                                                                	       
                                                                                                  �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K�
node_count�K�nodes�hhK ��h��R�(KK��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B�                            �0@�E�_��?�             e@������������������������       �        
             $@       8                    �?��<����?�            �c@       !                   �7@��ӭ�a�?H             R@                           �6@�,b+���?%            �B@                           @�ѳ�wY�?"             A@                           @��S�r
�?             <@                           �?�"w����?             3@	       
                      @>
ףp=�?
             $@������������������������       �                     @                          �3@����X�?             @                          �1@      �?             @������������������������       �      �?              @������������������������       �                      @                          �4@VUUUUU�?             @������������������������       �                     �?                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                           3@h/�����?	             "@������������������������       �                     �?                            �?      �?              @������������������������       ��q�q�?             @������������������������       �                      @                            �?�<ݚ�?	             "@������������������������       �                     @������������������������       �                      @                           �?      �?             @������������������������       �                     @                            �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @"       1                      @0J5y��?#            �A@#       &                    �?�a�2�t�?             2@$       %                    �?և���X�?             @������������������������       �                     @������������������������       �                     @'       0                   �@@�T�x?r�?             &@(       )                    �?      �?              @������������������������       �                      @*       /                     �?9��8���?             @+       ,                    <@VUUUUU�?             @������������������������       �                     �?-       .                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                     @2       3                    �?�t����?             1@������������������������       �                     @4       7                    @�n_Y�K�?             *@5       6                     @�q�q�?             (@������������������������       �և���X�?             @������������������������       ����Q��?             @������������������������       �                     �?9       T                    @}8�IL��?V            �U@:       M                     @�W�!l��?+            �E@;       J                     �?In�.P��?             ?@<       C                     �?P7�Z�?             3@=       >                    �?      �?              @������������������������       �                     @?       @                    7@VUUUUU�?             @������������������������       �                     �?A       B                    :@      �?              @������������������������       �                     �?������������������������       �                     �?D       E                    @}��7�?             &@������������������������       �                     @F       I                   �3@�$I�$I�?             @G       H                   �1@{�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �                      @K       L                    6@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?N       Q                    �?      �?             (@O       P                    5@z�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @R       S                    �?����X�?             @������������������������       ��q�q�?             @������������������������       �                     �?U       p                   �8@��&!�?+            �E@V       o                     @n�1�^�?"             A@W       `                     �?      �?              @@X       [                   �5@�
t�F��?             1@Y       Z                   �2@@4և���?             ,@������������������������       �z�G�z�?             @������������������������       �        	             "@\       _                    @VUUUUU�?             @]       ^                     �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?a       d                   �4@l�l��?             .@b       c                    @r�q��?             @������������������������       �                     @������������������������       �                     �?e       l                    �?�n���?	             "@f       g                   �5@0�����?             @������������������������       �                     �?h       i                    @r�q��?             @������������������������       �                     @j       k                   �6@      �?              @������������������������       �                     �?������������������������       �                     �?m       n                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @q       t                    @������?	             "@r       s                     �?�q�q�?             @������������������������       �                     �?������������������������       �                      @u       x                    �?�������?             @v       w                   �;@      �?              @������������������������       �                     �?������������������������       �                     �?y       |                    @      �?             @z       {                   �?@      �?              @������������������������       �                     �?������������������������       �                     �?}       ~                   �;@      �?              @������������������������       �                     �?������������������������       �                     �?�t�b�values�hhK ��h��R�(KKKK��hV�B@_         @      4@      �?       @      @      @      $@      @      �?       @       @      @      @      3@      �?      (@      @      @       @      &@       @      @      4@      ,@                                                                                                                                                                                      $@               @      4@      �?       @      @      @      $@      @      �?       @       @      @      @      3@      �?      (@      @      @       @      &@       @      @      $@      ,@              @              @      @      @      "@      @              �?      �?      @      @              �?      (@      @       @      �?      @      @      @      �?                      @              @      @      @      "@      �?                              @                      �?              @                      @                      �?                      @              @              @      "@      �?                              @                      �?              @                      @                      �?                      @              @              @      "@      �?                                                                       @                      @                      �?                      �?              @              @       @      �?                                                                       @                      @                      �?                      �?              @                      �?      �?                                                                       @                      �?                      �?                                      @                                                                                                                                                                              �?                                      �?      �?                                                                       @                      �?                      �?                      �?                                                                                                                       @                                              �?                      �?                                                                                                                                                                      �?                                                                                                                                               @                                                                                                              �?      �?                                                                                              �?                                                                                                                                                                                              �?                                                                                      �?      �?                                                                                                                                                                                              �?                                                                                                                                                                                      �?                                                                                                                                                                                      @      �?                                                                                                      @                                                                                      �?                                                                                                                                                                                      @                                                                                                              @                                                                               @                                                                                                              @                                                                               @                                                                                                                                                               @                                      @                                                                                                                                                                                              @                                                                                                                                                       @                                                                                                                                                                                                                                                                              @                      �?              �?                                                                                                                                                      @                                                                                                                                                                                                                      �?              �?                                                                                                                                                                              �?                                                                                                                                                                                                              �?                                                                                              @                                                                                                                                                                                                                      @              �?      �?              @                      (@      �?       @      �?              @      @                                                                              @              �?      �?              @                              �?       @      �?               @      @                                                                                                                      @                                                                      @                                                                                                                                                                                              @                                                                                                                      @                                                                                                                                                      @              �?      �?                                              �?       @      �?               @                                                                                                      �?      �?                                              �?       @      �?               @                                                                                                                                                                                               @                                                                                                      �?      �?                                              �?       @      �?                                                                                                                      �?      �?                                              �?                                                                                                                                                                                              �?                                                                                                                                      �?      �?                                                                                                                                                                                      �?                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                       @      �?                                                                                                      @                                                                                                                                                                                                                                                              (@                                      @                                                                                                                                                      @                                                                                                                                                                                               @                                      @                                                                                                                                                      @                                      @                                                                                                                                                      @                                      @                                                                                                                                                      @                                       @                                                                                                                                                      �?                                                                       @      1@      �?      @       @              �?       @      �?      �?      �?      �?              3@                              �?      �?      @      �?      �?      "@      ,@      �?      $@              @                                                                              �?                                      �?      @                      @      *@      �?      @              @                                                                              �?                                      �?                              @      *@      �?      @              @                                                                              �?                                      �?                              @       @      �?                                                                                                                                              �?                              @                                                                                                                                                                                              @              �?                                                                                                                                              �?                              �?              �?                                                                                                                                                                                                                                                                                                                                              �?                              �?                                                                                                                                                              �?                                                                                                                                                                                                                              �?                      @              @                                                                              �?                                                                               @              @                                                                                                                                                                                                              @                                                                              �?                                                                               @                               @                                                                              �?                                                                               @                               @                                                                              �?                                                                                                                                                                                                                                                                               @                               @                                                                                                                                                                                                                                                                                                                                                      �?      &@                                                                                                                                                                                              &@                                                                                                                                                                                      �?                      @                                                                                                                                              @                                              @                                                                                                                                              �?                                               @                                                                                                                                              �?                                               @                                                                                                                                                                                               @                                                                                                                                              @                                               @                                                                                                                                              @                                                                                                                                                                                              �?                                      �?      @      �?      �?       @              �?       @      �?      �?      �?      �?              2@                              �?                      �?      �?       @      �?      �?      @              �?       @              �?                                                      2@                              �?                              �?      �?      �?      �?      @              �?                      �?                                                      2@                              �?                              �?      �?      �?      �?      �?                                                                                              *@                              �?                              �?                              �?                                                                                              *@                                                                                              �?                                                                                              @                                                                                                                                                                                              "@                                                                                      �?                                                                                                                                      �?                              �?                      �?                                                                                                                                                                      �?                      �?                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                              �?                                                              @              �?                      �?                                                      @                                                                      �?      �?              @                                      �?                                                                                                                                                      @                                                                                                                                                                                                                                      �?                                                                                                                                                      �?              �?                                                                              @                                                                      �?      �?                              �?                                                                              @                                                                      �?                                                                                                                                                                                              �?                                      �?                                                                              @                                                                                                                                                                                              @                                                                                                              �?                                                                              �?                                                                                                                                                                                              �?                                                                                                              �?                                                                                                                                                                              �?                                                                                                                                                                              �?              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                       @                                                                                                                                                                              �?                                       @      �?      �?      �?      �?                                                                      �?              �?                                                                       @                                                                                                                      �?                                                                                                                                                                                              �?                                                                       @                                                                                                                                                      �?                                              �?      �?      �?      �?                                                                      �?                                                                                                      �?      �?                                                                                                                                                                                              �?                                                                                                                                                                                      �?                                                                                                                                      �?                                              �?                      �?                                                                      �?                                                                                              �?                      �?                                                                                                                                                                      �?                                                                                                                                                                                                                      �?                                                                                                                      �?                                                                                                                                              �?                                              �?                                                                                                                                                                                                                                                                                                                                              �?                        �t�bub�_sklearn_version��1.1.0�ub.