���     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.1.3�ub�n_estimators�M,�estimator_params�(�	criterion��	max_depth��min_samples_split��min_samples_leaf��min_weight_fraction_leaf��max_features��max_leaf_nodes��min_impurity_decrease��random_state��	ccp_alpha�t��	bootstrap���	oob_score���n_jobs�NhN�verbose�K �
warm_start��hN�max_samples�NhhhKhKhKhG        h�sqrt�hNhG        hG        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h5�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C�                                                                	       
                                          �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhKhKhKhG        hh.hNhJ�q�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��h>�f8�����R�(KhBNNNJ����J����K t�b�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFh2�scalar���h>�i8�����R�(KhBNNNJ����J����K t�bC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hK�
node_count�K�nodes�h4h7K ��h9��R�(KK��h>�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hwhZK ��hxhZK��hyhZK��hzh>�f8�����R�(KhBNNNJ����J����K t�bK��h{h�K ��h|hZK(��h}h�K0��uK8KKt�b�B�                             @8xl^]�?�	           ��@       	                     @��_��?           P�@                          �4@��-/�?I           D�@                           �?��4ɖ�?"           @�@������������������������       ���S�r��?H             \@������������������������       �0-C�&�?�           ��@                           �?�пɣ��?'           H�@������������������������       ��FQʱ��?�            pv@������������������������       ��J��1��?;           �@
                           �?L�Zi���?�           ��@                          �5@�Jä��?�             u@������������������������       ����.��?r            �f@������������������������       �qR�X���?_            `c@                           �?8�ȷ��?�            Px@������������������������       �m	�B�{�?�            �o@������������������������       �,�/��?X            �`@                           �?GG߄ �?�           ��@                            @2�F��?`           H�@                          �:@����ug�?�            �y@������������������������       ���c镕�?�            �v@������������������������       �     ��?              H@                           @�4_�g�?j             f@������������������������       �.؂-؂�?L             ^@������������������������       �����S��?             L@                           �?/!�����?!           ��@                            @4����g�?�            pw@������������������������       ���`so��?�            �k@������������������������       �m��!�D�?`             c@                          �;@�Ӷ�1�?0           ~@������������������������       �
�R\��?           `z@������������������������       ������?%            �M@�t�b�values�h4h7K ��h9��R�(KKKK��h��B�       �j@      <@     �A@      :@      Z@     Ȃ@      >@     P�@      *@      @     �W@      P@     H�@     }@      7@     `p@     �a@      *@      <@      6@      S@     �x@      .@     ��@      @      @      P@      B@     �@     pq@       @     `e@     �^@      (@      1@      4@     �M@     pr@      ,@     �{@      @      @      I@      >@     �t@      i@       @     �`@     �O@              "@      @      7@     `c@       @     @g@               @      2@      7@     �f@     �[@      @     �T@      $@               @               @       @              :@                       @      �?     �A@      $@              0@     �J@              @      @      5@     `b@       @      d@               @      0@      6@     `b@     @Y@      @     �P@     �M@      (@       @      0@      B@     �a@      @     �o@      @       @      @@      @     �b@     �V@       @     �I@      8@      (@      @      @      4@      K@      @     �U@       @              6@      @     �M@      >@       @      =@     �A@              @      $@      0@     �U@      @      e@      @       @      $@       @     �V@      N@              6@      3@      �?      &@       @      1@      Y@      �?     Pp@              �?      ,@      @     @f@     �S@              C@      &@      �?      $@      �?      &@     �M@      �?     @Y@                      "@      �?     �R@      F@              ,@      @      �?      @      �?      $@      C@      �?     �I@                       @      �?      @@      2@              &@      @              @              �?      5@              I@                      �?             �E@      :@              @       @              �?      �?      @     �D@              d@              �?      @      @     �Y@      A@              8@      @                      �?      @      :@             @Y@              �?      @      @      K@      =@              7@      �?              �?              @      .@             �M@                                     �H@      @              �?     �Q@      .@      @      @      <@     �i@      .@     `}@      @       @      >@      <@     �p@     @g@      .@     �V@      A@      @      @      �?      0@     �U@      "@     @f@      @      �?      $@      &@     �W@      P@      $@     �K@      5@      @      @      �?      "@     �P@      "@      X@      @      �?      $@      "@     @P@     �J@      @     �H@      5@      @      @      �?      "@      O@      "@     �S@      @      �?       @      "@     �M@      I@      @     �A@                                              @              2@                       @              @      @              ,@      *@       @      �?              @      3@             �T@      �?                       @      =@      &@      @      @      *@       @      �?               @      ,@             �I@      �?                       @      0@      $@      @      @                                      @      @              ?@                                      *@      �?              �?     �B@      $@      �?      @      (@      ^@      @     @r@      �?      �?      4@      1@     �e@     �^@      @      B@      5@      �?      �?      �?      @     �I@      �?     �b@      �?      �?      @      @     �Q@      H@       @      $@      1@      �?      �?      �?      @      ;@      �?     @S@      �?      �?      @       @     �F@      =@       @       @      @                              �?      8@             �R@                              @      :@      3@               @      0@      "@               @       @     @Q@      @     �a@                      ,@      (@     �Y@     �R@      @      :@      0@      "@               @       @      L@      @      ^@                      ,@      (@     �T@     �Q@      @      9@                                              *@              5@                                      4@      @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�^hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�=\q��?�	           ��@       	                   �<@���Q4�?3           l�@                           �?J<��MK�?�           \�@                            �?�E��/K�?�            @j@������������������������       ���:����?)            @Q@������������������������       �-�l�J�?W            �a@                           �?��K��V�?d           �@������������������������       ��`�ה��?�            �s@������������������������       �5}�[�?�           (�@
                           �?�_hD���?O            �`@                            �?�q�q�?             8@������������������������       ���Q��?             $@������������������������       ��)x9/�?             ,@                           @�X;�U��?A             [@������������������������       �<�7�QJ�?+            �R@������������������������       �@�_)P��?            �@@                           �?�����?M           ܠ@                          �5@'�ݞ4K�?�            �v@                          �3@��E���?w            �h@������������������������       �'��O�?R            �`@������������������������       �Ti�?%            �O@                            @�������?k            �d@������������������������       ��8
|y�?Q            �_@������������������������       ��GcT!)�?             C@                            @e֚�1��?k           �@                           @˳���H�?(           �@������������������������       �sdnoo�?�           ��@������������������������       ����&�?W             a@                          �2@���N��?C           �@������������������������       ��m�}k��?L            �]@������������������������       ��g�PM��?�            Px@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        g@      8@     �F@      6@      ]@     ��@      C@     x�@      2@      @     �S@     �O@     ��@     8�@      5@     �p@      Y@      (@     �@@      *@      Q@     �s@      7@     �z@      "@      @      D@      <@     Pr@     �m@      0@     �a@     @V@      &@      >@      *@      P@     �r@      7@     @w@      "@      @     �A@      ;@     `q@      l@      0@     �`@      &@              @      �?      @      4@             �P@      @              @      @     �E@      6@              3@      @                                      @              =@                      @      @      0@      @              @      @              @      �?      @      1@              C@      @              @      @      ;@      0@              .@     �S@      &@      :@      (@      M@     @q@      7@     s@      @      @      <@      4@     `m@     `i@      0@     @\@      *@       @      (@      @      &@     �P@      @     �S@              �?      @      �?      >@      I@       @     �A@     @P@      "@      ,@       @     �G@     @j@      1@     @l@      @       @      9@      3@     �i@      c@      ,@     �S@      &@      �?      @              @      1@              L@                      @      �?      .@      &@               @       @                                       @              @                      @                      @                                                              @              @                      @                                               @                                      @              @                                              @                      "@      �?      @              @      "@             �H@                      �?      �?      .@       @               @      @      �?      @              @      "@              B@                      �?      �?       @      @               @       @                              �?                      *@                                      @      @              @      U@      (@      (@      "@      H@     �u@      .@     ��@      "@      @      C@     �A@     p{@     �q@      @      `@      1@      �?      @              "@     �J@      @     �W@                      @       @     �T@      O@      @      :@      .@              @              �?      8@      �?     �H@                      @              N@      6@      @      1@      (@               @                      1@      �?      E@                      @              C@       @      @      "@      @              �?              �?      @              @                                      6@      ,@               @       @      �?                       @      =@      @     �F@                       @       @      7@      D@              "@       @      �?                      @      9@      @      <@                       @       @      4@      =@              "@                                      @      @              1@                                      @      &@                     �P@      &@      "@      "@     �C@     `r@      $@     ��@      "@      @     �@@     �@@     @v@     �k@       @     �Y@     �L@      &@       @      @     �B@      i@      "@     `x@      @       @      =@      :@     �m@     �f@      �?     @U@     �K@      &@      @      @     �B@     @g@       @     �t@      @       @      6@      7@      k@     �d@      �?     �S@       @               @       @              .@      �?     �M@      �?              @      @      4@      2@              @      $@              �?       @       @     @W@      �?     �i@      @       @      @      @     �]@      C@      �?      1@      @                                      1@              F@                      �?             �D@      $@               @      @              �?       @       @      S@      �?     @d@      @       @      @      @     �S@      <@      �?      .@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJTG�NhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @J'�N2��?�	           ��@       	                     �?Ԙ��]�?�           �@                           �?Sn�*k��?5           f�@                          �0@Q�*pl��?�           ��@������������������������       ��~�F&K�?             K@������������������������       ���Ϫ�y�?�           @�@                           �?�ݾ[#d�?�           T�@������������������������       ���TdD�?�           h�@������������������������       ���:zp��?           @�@
                          �;@C7 -7�?�           (�@                           �?��#\V1�?�           8�@������������������������       �dЅҶ9�?�             r@������������������������       ��� �	��?�            Pv@                           @~it��?#             O@������������������������       �     ��?             @@������������������������       ��0u��A�?             >@                           @)�� ��?�           D�@                           �?�,�B��?"           p�@                           �?7BK]M��?<            @������������������������       ��Ë'o�?�             i@������������������������       ��F����?�            �r@                           @��Ѓ���?�            �w@������������������������       ��D�d@6�?J            �]@������������������������       ��+�\���?�            Pp@                          �:@V�|�&��?�            `l@                           �?�����?u            @f@������������������������       ��K0��?*            �Q@������������������������       �XB1B&�?K            �Z@                           �?ѷī�?!            �H@������������������������       �]�l8b��?            �A@������������������������       �x9/���?	             ,@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      <@     �B@      9@     �]@     @�@      D@     P�@      0@      @     �T@      N@     ��@     �@      ,@     0p@      f@      1@      :@      1@      X@     }@      @@     `�@      .@      @     �R@     �G@     P@      x@      (@     �k@     �`@       @      .@      $@      M@     �w@      4@     X�@      $@              D@      >@     @x@     �p@       @      c@      M@               @      @      ,@     �a@      @     �e@      @              1@      $@     �\@      Q@      @     �H@                      �?      �?      @      .@      @      @                              @      @      *@                      M@              @       @      &@     @_@             @e@      @              1@      @      [@     �K@      @     �H@     �R@       @      @      @      F@     �m@      .@     �y@      @              7@      4@     q@     �h@      @     �Y@     �F@      @      @       @      :@     �Z@      @     @b@      @              "@      (@      Z@     �R@      �?     �D@      >@      @              @      2@      `@       @     �p@       @              ,@       @      e@     @^@      @      O@      F@      "@      &@      @      C@     @V@      (@      `@      @      @     �A@      1@     @\@     �^@      @     @Q@     �C@      "@      &@      @      C@     �T@      &@     �Y@      @      @      A@      1@     @Y@     @\@      @     �P@      ,@      @      @      @      4@     �G@      @     �B@      @      @      @      (@      H@      G@       @      @@      9@      @      @      @      2@      B@      @     �P@      �?      �?      ?@      @     �J@     �P@       @     �A@      @                                      @      �?      :@                      �?              (@      "@               @      �?                                      @      �?      &@                      �?               @      @                      @                                       @              .@                                      @      @               @      >@      &@      &@       @      6@     �f@       @     �x@      �?      �?      @      *@     p@     @^@       @      C@      7@      @      $@       @      3@     �a@      @     0t@      �?              @       @     �j@     �S@      �?      B@      ,@      @      @      @      *@     @S@      @     @g@      �?              @       @     �X@     �K@      �?      3@      @      @      @              "@      B@       @      M@      �?              @      @      A@      ?@      �?       @      @      �?      @      @      @     �D@      @      `@                              @     @P@      8@              &@      "@      �?      @       @      @     @P@      �?      a@                       @             @\@      7@              1@       @              �?               @      8@      �?      =@                                     �H@      @              @      @      �?      @       @      @     �D@              [@                       @              P@      1@              (@      @      @      �?              @     �D@       @     @Q@              �?      �?      @     �F@     �E@      �?       @      @      @      �?              @      @@       @     �F@              �?      �?      @     �A@      D@      �?       @      �?      @      �?              @      (@       @      (@              �?              @      0@      0@              �?      @      @                              4@             �@@                      �?       @      3@      8@      �?      �?      @                                      "@              8@                                      $@      @                      @                                      @              4@                                      @       @                                                              @              @                                      @      �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJS��}hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx         
                   �;@qM�&X�?�	           ��@       	                    !@I��2y�?�           "�@                           �?R�X)w�?�           ��@                            @b�����?�           ��@������������������������       �U��q�G�?�           �@������������������������       ��!���Y�?           `z@                          �8@^4#T��?�           h�@������������������������       �T̤���?1           �@������������������������       �Z�w��4�?�            0q@������������������������       ���Z�Y�?             7@                           @�'lbe��?           �{@                           @�܈�L�?�            �x@                            @��3�?�            �s@������������������������       ���U�o�?�            �k@������������������������       ��9�?�x�?=            �V@                           �?������?2            @T@������������������������       �����!p�?             6@������������������������       �����˵�?$            �M@                          �<@�U_���?             G@                           �?��a�2��?             2@������������������������       ���ˠ�?             &@������������������������       �����X�?             @                            �?h�����?             <@������������������������       ��z�G��?             $@������������������������       �B{	�%��?             2@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      D@     �E@     �@@     �Y@     x�@      B@     x�@      0@      @     �S@      L@     ��@     P�@      (@     @n@      f@     �A@      D@      @@     �W@      �@     �A@     P�@      (@      @      Q@      K@     ��@     ~@       @     �j@     �e@     �A@      D@      @@     �W@     Ѐ@     �A@     8�@      (@      @      Q@      K@     �@     �}@       @     `j@     �S@      3@      :@      3@      K@     �p@      4@      w@      @       @      <@      >@      q@      i@      @      Z@     �L@      (@      3@      1@     �D@     �i@      .@     �n@      @       @      3@      9@     �g@     @b@      @      U@      6@      @      @       @      *@      O@      @     �_@      @              "@      @     �U@     �K@              4@      X@      0@      ,@      *@     �D@     �p@      .@     ��@      @      �?      D@      8@     �x@     0q@      @     �Z@     �U@      (@      ,@      (@     �@@      o@      ,@     @�@      @      �?      A@      5@     �s@     `k@      @     �X@      $@      @              �?       @      5@      �?     @S@                      @      @     �S@      L@              "@       @                                      $@              @                                      �?      @               @      6@      @      @      �?       @     �R@      �?     �f@      @      �?      $@       @      K@     �D@      @      =@      6@      @      @      �?       @      Q@      �?     �b@      @      �?      "@       @     �G@     �D@      @      <@      0@      @      @      �?       @      H@      �?     �_@      @      �?      "@       @     �C@      4@      @      :@      .@      @      �?      �?       @     �B@      �?      U@                      "@      �?      8@      3@      @      4@      �?               @              @      &@              E@      @      �?              �?      .@      �?      �?      @      @                                      4@              8@                                       @      5@               @                                              �?               @                                       @      &@                      @                                      3@              0@                                      @      $@               @                                              @              >@                      �?              @                      �?                                              @              "@                      �?               @                      �?                                              @              @                      �?                                      �?                                                              @                                       @                                                                       @              5@                                      @                                                                                      @                                      @                                                                       @              ,@                                       @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��PDhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B(                             !@X8�(>��?�	           ��@       	                   �;@�!�2�?�	           `�@                            @I����?w           �@                            �?Xs2��?!           ��@������������������������       �T���?�           l�@������������������������       �!����?�           ��@                           @?�p��?V           ��@������������������������       ����%��?O           @�@������������������������       ��h$��W�?             .@
                           �?V^-+�c�?           �z@                           �?�����?$             N@������������������������       �c}h���?             <@������������������������       �     P�?             @@                            @2	����?�             w@������������������������       �+�C3O��?�            @o@������������������������       ������?P            �]@                           @�I+��?             9@������������������������       �     ��?             0@������������������������       ������H�?             "@�t�bh�h4h7K ��h9��R�(KKKK��h��B�	       �k@      7@      C@      @@     �X@     ��@     �A@     ��@      8@      @      S@      N@     H�@     `@      4@     �p@     �k@      7@      C@      @@     @X@     ��@      A@     ��@      8@      @      S@      N@     @�@     @@      4@     pp@      h@      5@     �A@      ?@     �T@     0�@      ?@     @�@      *@      @      N@      M@     8�@     �}@      3@     `n@      d@      1@      <@      <@     �P@     �|@      7@     ��@      (@      @     �K@     �H@     0y@     0v@      3@     `i@      ]@      ,@      2@      5@      F@      v@      0@     �@      $@             �D@     �@@     �s@     `n@      "@     �`@     �F@      @      $@      @      7@      Z@      @      \@       @      @      ,@      0@      V@      \@      $@      Q@      ?@      @      @      @      .@     �c@       @     `u@      �?              @      "@     �j@     �]@              D@      ?@      @      @      @      .@      c@       @     `u@      �?              @      "@     �i@     �\@              D@                                              @                                                       @      @                      <@       @      @      �?      .@     �R@      @      d@      &@              0@       @     @P@      ;@      �?      4@      @      �?                      �?      .@              ,@                      @              @      @              @      @                                      @              @                      @               @       @                      �?      �?                      �?      &@              @                                      @      @              @      5@      �?      @      �?      ,@     �M@      @     @b@      &@              "@       @     �M@      5@      �?      1@      0@      �?      @      �?      "@     �A@      @     �V@      @              "@       @     �E@      2@              ,@      @                              @      8@             �K@      @                              0@      @      �?      @                                      �?      (@      �?      @                                      �?       @              @                                              $@              @                                              �?               @                                      �?       @      �?                                              �?      �?              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�u1KhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �7@cҭG%}�?�	           ��@       	                     @�q�$��?�           ��@                            �?���+�(�?           ��@                           �?Z`B����?�           |�@������������������������       ���uX���?�           �@������������������������       �������?           ��@                          �5@�.r#P��?N           8�@������������������������       ���ŉ��?           Pz@������������������������       �@�[�0��?B            �X@
                          �6@z�=����?�           �@                           @���Q��?�           8�@������������������������       ��R>�V�?=           �}@������������������������       �U���J�?�            �i@                           �?r�q��?,             N@������������������������       ��s�n_�?            �C@������������������������       �"�����?             5@                           �?��Hx��?�            �@                           @^/`���?9           0}@                          �;@C�N ��?$            {@������������������������       �� ˉy��?�            �r@������������������������       ���=��?c            �`@������������������������       �c��[�m�?            �A@                           @��0�;�?�           h�@                           �?��d�v�?�            �w@������������������������       �ZZZZZZ�?�            �m@������������������������       �h�"C�k�?a            �a@                          �=@�M�b���?�            s@������������������������       ����PU��?�            �k@������������������������       ��m�'�*�?2            �T@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@      7@     �D@      7@     �T@     ��@      >@     t�@      2@      (@     �W@     �Q@     Ї@      �@      ,@     pp@     �b@      .@     �C@      .@     �L@     �z@      9@     `�@      &@      @     �Q@     �O@     �@     px@      &@      h@      ^@      (@      ;@      "@     �G@     �s@      5@     �}@      $@      @      O@      K@      x@     �r@      $@     �d@     �V@      $@      2@      @      9@     �m@      1@     �x@      @       @     �F@      C@     Ps@      j@      @      U@     �I@      @      0@      @      4@     �[@      &@     @a@      @       @      ?@      <@     �_@      U@      @     �C@      D@      @       @      @      @      `@      @     0p@      �?              ,@      $@     �f@      _@      @     �F@      =@       @      "@       @      6@      S@      @     @T@      @      @      1@      0@     @S@     �V@      @     �T@      4@      �?      @              0@      Q@      @     �P@       @       @      ,@      ,@     �P@     @P@      @     �R@      "@      �?      @       @      @       @              ,@       @       @      @       @      &@      9@              "@      ?@      @      (@      @      $@     @[@      @     �p@      �?      �?       @      "@     `c@     @W@      �?      :@      ?@      @       @      @      $@     �Y@      @     �o@      �?      �?      @      @     �a@     @S@              9@      9@      @       @      @      @      R@      @      e@      �?      �?      @      @     @W@     �N@              3@      @                      �?      @      >@             �U@                      @      �?      I@      0@              @                      @                      @              .@                       @       @      (@      0@      �?      �?                      @                      @               @                       @              @      *@              �?                                               @              @                               @      @      @      �?              O@       @       @       @      9@     �j@      @     w@      @      @      9@      @     �k@     @^@      @     �Q@      @@      @       @      @      1@     �U@       @     ``@      @       @      @      �?     �T@     �I@              E@      @@      @       @      @      1@     �S@       @      \@      @       @      @      �?     @T@     �H@             �B@      3@       @              @      &@      P@       @     �P@      @       @      @      �?      N@      >@              ;@      *@       @       @              @      .@             �F@      �?              �?              5@      3@              $@                                              @              3@                                       @       @              @      >@      @              @       @      `@      @     �m@      @      @      4@      @     @a@     �Q@      @      <@      9@      @               @       @      N@      @     �a@      �?      �?      $@      @      M@     �C@      @      8@      .@      @                      @     �C@      @      S@              �?      @       @     �@@      <@      @      6@      $@                       @       @      5@              P@      �?              @      �?      9@      &@               @      @      �?              �?              Q@             �X@       @       @      $@      @      T@      ?@              @      @      �?              �?              K@             @S@               @      @      @      G@      8@              @                                              ,@              5@       @              @              A@      @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJW@1hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?6!q2���?�	           ��@       	                   �;@�Y>.F�?W           ؚ@                          �1@�G��<]�?�           �@                           �?�yE��?�            @s@������������������������       �����1�?T            �\@������������������������       ��CD���?|            @h@                           �?;���?           @�@������������������������       �=原�?l            �c@������������������������       �^~Q�+�?�           А@
                            �?�cx��?n            @f@                            �?f�nOwA�?:            �X@������������������������       �2���Q�?             G@������������������������       �;�;��?!             J@                           @�z�Ga�?4             T@������������������������       �(;5��>�?%            �K@������������������������       �����Mb�?             9@                           @�t=Ի4�?X           &�@                            @�˜o7	�?E           ��@                           @�8�$���?�           Є@������������������������       ��:����?B           X�@������������������������       �M:���Q�?a            �a@                           �?}=��l��?�            �o@������������������������       �` � ���?\            �a@������������������������       �d}h���?F             \@                          �:@�3C�;�?           �@                            @(�5���?�           T�@������������������������       �
�I��?�           X�@������������������������       �dH��@�?�            �p@                           @����1�?�            �l@������������������������       ��/M����?t            `h@������������������������       ���a�2��?             B@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        j@     �@@     �E@      5@     �Z@     x�@      A@     ��@      7@       @     �W@      T@     H�@     x�@      2@     0p@     @Z@      5@      ;@      $@      K@     �t@      2@     �x@      ,@      @      F@      F@     �q@     �l@       @      `@      W@      2@      9@      $@      H@     0s@      2@     @t@      *@      @     �A@      E@     �p@     @j@       @     @^@      7@      @       @              $@     �N@      $@      G@       @       @      @      $@     �C@      F@      @     �C@      $@       @      @              @      @@       @      *@       @              �?      @      &@      4@               @      *@       @      @              @      =@       @     �@@               @      @      @      <@      8@      @      ?@     @Q@      ,@      1@      $@      C@     �n@       @     `q@      &@       @      <@      @@     @l@     �d@      @     �T@      &@       @                      @      2@              I@      @              @      �?     �@@      2@              (@      M@      (@      1@      $@     �A@     �l@       @     �l@      @       @      8@      ?@      h@     �b@      @     �Q@      *@      @       @              @      :@              R@      �?              "@       @      0@      4@               @      @      @       @              @      4@              ?@                      "@               @      (@              @                                      �?      &@              4@                      @              @      @               @      @      @       @               @      "@              &@                      @              @       @               @      @                              @      @             �D@      �?                       @       @       @              @      @                              @      @              8@      �?                       @      @      @               @      @                                      �?              1@                                      �?      �?               @      Z@      (@      0@      &@     �J@      v@      0@     ��@      "@      @      I@      B@      {@     �r@      $@     @`@      K@      @      "@      @      6@      a@       @     �p@              �?      (@      .@      k@      [@      @      N@     �G@      @      @      @      0@     @Z@       @      f@                      "@      *@      a@     @W@      @     �H@     �E@      @      @      @      (@      V@      �?     �^@                      @      $@     �[@     @S@      �?     �D@      @              @       @      @      1@      �?      K@                      @      @      :@      0@       @       @      @               @      �?      @      @@              W@              �?      @       @     @T@      .@              &@       @                      �?      �?      $@              H@                      �?      �?      K@      *@              $@      @               @              @      6@              F@              �?       @      �?      ;@       @              �?      I@      "@      @      @      ?@      k@      ,@     �x@      "@      @      C@      5@     �j@     �g@      @     �Q@     �G@      "@      @      @      ;@     �c@      *@     �r@      @       @      >@      3@     `f@     �e@      @      N@     �C@       @      @      @      5@     @_@      (@     �h@      @       @      >@      .@      ^@     `a@      @     �H@       @      �?              �?      @      A@      �?     @Z@      �?                      @     �M@     �A@              &@      @                              @      M@      �?     @V@      @      �?       @       @      B@      .@              $@      @                              @     �D@      �?     �T@      @      �?       @       @      9@      .@              "@                                              1@              @      �?                              &@                      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��ShG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �=@�}����?�	           ��@                           �?�̭bܦ�?+	           ެ@                           !@�aى��?*           �@                           �?ض� `�?#           ��@������������������������       �����!�?[           0�@������������������������       �.z����?�           H�@������������������������       �����2�?             .@                           �?�+q��?           ��@	       
                     @q�G_��?�            �r@������������������������       �z\�ܯ�?�            �k@������������������������       ����(\��?5             T@                           @�����?E           �@������������������������       ��1�.��?%           �@������������������������       ��Ӗ$��?            �{@                           �?w��WZ�?�            @k@                          �>@�Ϣ��3�?0            �Q@                            @��,d!�?             7@������������������������       �*L�9��?             &@������������������������       ��������?             (@                           �?��8��x�?"             H@������������������������       �I�$I�$�?             <@������������������������       ��������?             4@                           @���;���?\            `b@                          @@@)il;��?V            �`@������������������������       ���Ü�o�?=            �V@������������������������       ��R(�?            �E@������������������������       ��]�`��?             *@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@     �D@      C@      2@      Z@     ��@      <@     �@      =@      &@     �T@      M@     �@     x�@      1@     �p@     @g@      D@      C@      2@      X@      �@      <@     ��@      8@      "@     @T@      M@     8�@     �@      1@     �o@     @Y@      4@      ;@      (@     �K@     �t@      0@     �w@      .@      @     �B@      =@     `s@      k@      @     �\@     @Y@      4@      ;@      (@      K@     0t@      (@     �w@      .@      @     �B@      =@     `s@     �j@      @     @\@     �B@       @      3@      @      5@     �T@             @b@      @       @      2@      @     @X@     �P@              C@      P@      (@       @      @     �@@      n@      (@      m@      "@      @      3@      9@     �j@     �b@      @     �R@                                      �?       @      @                                                      �?              �?     @U@      4@      &@      @     �D@     Ps@      (@     ȃ@      "@      @      F@      =@     w@     �r@      (@     �a@      .@               @      �?      *@     �F@      �?     @Q@                      @       @      O@     �K@      @      >@      ,@                      �?      (@     �@@             �C@                      @       @     �H@      E@      @      7@      �?               @              �?      (@      �?      >@                                      *@      *@              @     �Q@      4@      "@      @      <@     �p@      &@     ��@      "@      @      D@      ;@     0s@     �n@       @     �[@      O@      &@      @      @      2@      g@       @      |@      @       @      9@      5@     �l@     �d@      @     @T@       @      "@      @       @      $@      T@      @     �\@      @       @      .@      @      S@      T@      �?      >@      @      �?                       @      >@              U@      @       @      �?              K@      (@              ,@      @                              @       @              ;@                                      &@      @              @      @                              @      @               @                                       @       @                      @                               @      @              @                                                                                                      @                      @                                       @       @                      @                              �?      @              3@                                      "@      @              @       @                                      @               @                                      @      �?              @      �?                              �?                      &@                                       @      @               @      �?      �?                       @      6@             �L@      @       @      �?             �E@      @              @      �?      �?                       @      3@              K@               @      �?             �D@      @              @              �?                              2@              C@                      �?              :@       @              @      �?                               @      �?              0@               @                      .@      @               @                                              @              @      @                               @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ,�M.hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @���e��?�	           ��@       	                    �?6������?�           L�@                            �?�w>�?c�?           ��@                           @1��.�?Y           ��@������������������������       �nE<���?Q           p�@������������������������       ��ѳ�w�?             1@                           @���)���?�             s@������������������������       ��_v����?�            0p@������������������������       �Q2�����?            �F@
                          �;@t��n�?�           ܘ@                            �?^�t���?j           �@������������������������       �V�_V$�?�           �@������������������������       �������?�            �t@                            �?��E\��?s            �f@������������������������       ���XH��?,            @R@������������������������       �5zDن�?G             [@                           �?`*g�N4�?�           ��@                           �?Bx��Z�?3           �}@                           @��L����?3            �U@������������������������       �3�E��?'            @P@������������������������       �v�"���?             5@                           @�3
��L�?            @x@������������������������       ����b���?�            `l@������������������������       ����	�R�?g             d@                          �2@�t����?t           H�@                          �0@�qc&�O�?j            �e@������������������������       �)O���?             2@������������������������       ���	ɕo�?^            `c@                           @��,�5r�?
           �y@������������������������       �d[���?�            �r@������������������������       ����۾%�?L             ]@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@     �B@      B@      A@     @\@     ��@      1@     ��@      5@      0@     �P@      G@     p�@     �@      7@     `p@     �c@      :@      ;@      >@     �U@      �@      *@     ȅ@      1@      (@     �N@      D@     `�@     �x@      4@      j@     @U@      @      0@      1@     �H@     �m@      "@     pp@      &@       @      4@      7@      l@     `e@      @     �\@     �P@       @      (@      $@     �C@     @h@      @     �i@      @      @      .@      1@     �e@      _@      @     �T@     �O@       @      (@      $@     �B@      h@      @     �i@      @      @      .@      1@     �e@     �]@      @      T@      @                               @      �?       @      �?                                              @               @      3@      @      @      @      $@      F@      @      M@      @      @      @      @     �I@     �G@      @     �@@      .@      @      @      @      @     �B@      @      J@      @      @      @      @     �G@     �@@      @      >@      @              �?      @      @      @              @                                      @      ,@              @     �Q@      3@      &@      *@     �B@      q@      @      {@      @      @     �D@      1@     �t@     �k@      *@     �W@      Q@      0@      &@      &@     �B@     �n@      @      w@      @      @     �B@      ,@      r@     �i@       @     @V@     �I@      (@      @      &@      6@     @g@       @     �s@       @              ,@      &@     `m@     �b@      @      M@      1@      @      @              .@     �M@      �?     �J@      �?      @      7@      @     �K@      L@       @      ?@      @      @               @              =@      �?     �P@      @              @      @      E@      .@      @      @       @                                      @              7@      �?               @       @      :@      &@                      �?      @               @              7@      �?     �E@       @               @      �?      0@      @      @      @     �B@      &@      "@      @      ;@     �g@      @     �v@      @      @      @      @     @l@      \@      @     �J@      2@      @      @      �?      4@     �W@      @     @`@      @      �?      @      @     �U@     �P@       @      @@      �?              �?              @      ,@              7@                      �?              (@      4@              $@      �?              �?              @      *@              $@                      �?              "@      0@              $@                                              �?              *@                                      @      @                      1@      @       @      �?      0@     @T@      @     �Z@      @      �?       @      @     �R@     �G@       @      6@      ,@      @       @              $@      I@      @      K@      @      �?              @      D@      =@       @      (@      @      @              �?      @      ?@             �J@                       @              A@      2@              $@      3@      @      @      @      @     @W@      �?     �m@      �?      @       @      @     �a@     �F@      �?      5@      "@               @      @      �?      8@             �L@                      �?             �K@      ,@              @                                               @              "@                                      @      �?               @      "@               @      @      �?      6@              H@                      �?             �I@      *@              @      $@      @      @              @     @Q@      �?     `f@      �?      @      �?      @     @U@      ?@      �?      ,@      "@      @      @              @     �D@      �?     @a@      �?      @      �?              N@      1@              (@      �?      �?                              <@             �D@                              @      9@      ,@      �?       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ>��zhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @��P����?�	           ��@       	                    �?JN#�:�?�           "�@                           @B�lެ��?           �@                          �<@˻�����?@            �@������������������������       ��BeI��?#           �~@������������������������       �du�9d�?            �H@                           @$BӒY�?�           �@������������������������       �By�Oo|�?j            �e@������������������������       ��!�h��?]           ��@
                            �?�^?��?�           @�@                           @�.�.��?�           ��@������������������������       ���y�):�?0            �@������������������������       �ݚ)3�?�             r@                           �?0��/���?�            �v@������������������������       ���Y��Y�?            �C@������������������������       � 8���?�            Pt@                           �?���0Q,�?�           ��@                           @�WG1}�?*           �|@                           @�X���?�             v@������������������������       �����̌�?�             n@������������������������       �s
^N�K�?J             \@                          �8@-��S��?A            �Z@������������������������       ����J�?6            @V@������������������������       �����K�?             2@                           �?��r���?�           h�@                          �;@�����E�?�            @y@������������������������       �� �R��?�            pu@������������������������       �%}}���?"            �N@                          �8@��-�?�             k@������������������������       ��ˠT�?d            @c@������������������������       �lp����?&            �O@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        k@     �@@      C@      3@     �]@     x�@      ?@      �@      &@      @      X@     �O@      �@     P@      2@     s@     `e@      :@      B@      0@     @W@     �}@      :@     ��@      "@      @      R@      M@     �}@     �w@      2@      p@     @U@      *@      <@      @     �J@      m@      (@     @q@      @      @      @@      A@     �i@      f@      (@     �\@     �C@      @      0@       @      5@     �T@      @     �]@       @              .@      "@     �Q@     @W@      @     �O@     �C@      @      ,@       @      1@     �Q@      @      W@       @              .@      "@     @Q@      W@      @      O@                       @              @      *@              :@                                       @      �?              �?      G@      "@      (@      �?      @@     �b@      @     �c@      �?      @      1@      9@     �`@      U@      "@     �I@      $@      �?      @              @      F@      @      F@                      @      @      ?@      ,@      @      @      B@       @       @      �?      <@     @Z@      @     �\@      �?      @      ,@      5@     �Y@     �Q@      @      F@     �U@      *@       @      *@      D@     �n@      ,@     �{@      @      �?      D@      8@     �p@     �h@      @      b@      M@      *@      �?      &@      8@     �h@      (@     `w@      @              2@      0@     �k@     @a@      @     �W@      J@      (@      �?      @      3@     `d@       @     �p@      @              *@      $@     @e@     �\@       @      N@      @      �?              @      @      B@      @     @[@       @              @      @     �I@      7@       @      A@      <@              @       @      0@     �F@       @      R@      �?      �?      6@       @     �G@     �N@       @      I@      @              @      �?       @      �?              @                      @              $@      @              @      8@              @      �?      ,@      F@       @     @Q@      �?      �?      2@       @     �B@      K@       @      G@     �F@      @       @      @      :@     `f@      @     `w@       @              8@      @     �m@     @_@             �G@      >@      @       @       @      1@      U@      @     @^@                      2@      �?     �X@     �I@              =@      <@      @       @              &@     �R@      @      T@                      "@      �?     �S@     �B@              :@      4@      �?       @               @     �I@       @     �H@                      "@             �M@      6@              1@       @       @                      @      7@      �?      ?@                              �?      3@      .@              "@       @                       @      @      $@             �D@                      "@              4@      ,@              @       @                       @      @      @             �C@                      "@              *@      (@               @                                       @      @               @                                      @       @              �?      .@      @              �?      "@     �W@       @     �o@       @              @      @     @a@     �R@              2@      "@       @              �?      @     �O@       @     �f@                      @      @     �Q@      F@              1@      "@       @              �?      @      G@       @      b@                      @      @      Q@      F@              .@                                      �?      1@              C@                                      @                       @      @       @                       @      @@             �Q@       @              @      �?     �P@      >@              �?      @       @                       @      8@             �F@                      @      �?      J@      2@              �?                                               @              :@       @                              .@      (@                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJH[xhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @��̬x�?�	           ��@       	                     �?����?�           ��@                          �0@*������?}           �@                           @     ,�?,             P@������������������������       �^����T�?            �C@������������������������       ��{�Pk�?             9@                          �<@B�$w���?Q           �@������������������������       �p��&^��?           8�@������������������������       ��IQu`��?6            �V@
                            �?���ai�?b           @�@                           @%����?�           Ԑ@������������������������       ��Y8�	�?�           P�@������������������������       �c6=w��?0            �R@                           @ ������?�           ؄@������������������������       �l������?�             i@������������������������       �R���5��?-           0}@                           �?� b�?�           ��@                          �<@�[����?B           �@                          �1@�
:u4��?"           `|@������������������������       � x��6�?)            �P@������������������������       ��b���?�            @x@                          �=@�d��0�?              N@������������������������       ��n����?             2@������������������������       ��!͎�?             E@                           @i�x0�?�           ��@                          �2@��&�{�?�            q@������������������������       �VUUUUU�?=             X@������������������������       �XL!5ڰ�?n             f@                          �>@���r��?�            Pv@������������������������       �JwO��?�            Pu@������������������������       �     @�?	             0@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        j@      2@      B@      =@     �]@      �@     �E@     ��@      0@      @      R@      P@     ��@     �|@      6@     �p@     �c@      ,@      <@      7@     �V@     |@      A@     0�@      (@      @     �P@      M@      �@     �u@      4@     �j@     �F@      @      @      $@      <@     @d@      .@     s@      @              "@      &@     �n@     @]@      @      K@      �?                       @      @       @      @      @                              �?      *@      ,@              $@                                              @      @       @                              �?      @      *@              @      �?                       @      @      �?              @                                      @      �?              @      F@      @      @       @      7@     @c@      (@     �r@      @              "@      $@      m@     �Y@      @      F@     �E@      @      @       @      7@      b@      $@      p@       @              "@      $@     �j@     @X@      @     �B@      �?                                      "@       @      E@      @                              4@      @              @     �\@      @      6@      *@      O@     �q@      3@     Py@      @      @     �L@     �G@     �r@     �l@      .@     �c@     @P@      @      $@      $@      =@     �j@      "@     Pp@       @       @      ?@      7@     `g@     @a@      @     �U@      P@      @      $@      $@      <@     �i@      @     �l@       @       @      ?@      4@     �f@     �_@      @     �S@      �?                              �?      $@      @      ?@                              @      @      &@               @     �H@      @      (@      @     �@@     @R@      $@      b@      @       @      :@      8@     �[@     �V@       @     @R@      $@      @      @      �?      @      2@       @      B@      @              &@      @     �B@      :@      @     �A@     �C@      �?      @       @      <@     �K@       @      [@       @       @      .@      4@     �R@      P@      @      C@      I@      @       @      @      <@     `h@      "@     �y@      @      �?      @      @      n@     @]@       @      L@      <@      @      @      �?      0@     @W@       @      d@       @              @      @     @Z@     �J@              =@      .@      @      @      �?      (@     �U@       @     `a@       @              @       @      Y@     �H@              9@      @      �?      �?              �?      .@      @      9@                      �?       @      @      @              @      &@       @      @      �?      &@      R@      @     �\@       @              @              X@     �F@              4@      *@                              @      @              6@                               @      @      @              @      @                                                      &@                                              @                      "@                              @      @              &@                               @      @      �?              @      6@      �?       @      @      (@     �Y@      �?     @o@       @      �?      �?       @      a@      P@       @      ;@      @              �?       @      @      :@             �_@              �?      �?             @Q@      7@              1@      @                       @              (@             �A@                                     �B@      @              �?                      �?              @      ,@             �V@              �?      �?              @@      2@              0@      2@      �?      �?      @      "@      S@      �?      _@       @                       @     �P@     �D@       @      $@      0@      �?      �?      @      "@     �R@      �?      ^@      �?                       @     �M@     �D@       @      $@       @                                      �?              @      �?                               @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJe�]hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @��Ir���?�	           ��@       	                    �? �3���?�           f�@                            �?w�����?           X�@                           @6|�����?�             z@������������������������       �!�Zz/��?z            @h@������������������������       ���E���?�            �k@                           @�~u���?	           ��@������������������������       �-��6��?�           Ї@������������������������       �<+	���?%             N@
                            �?��H��g�?�           t�@                           @.���|�?x           8�@������������������������       �����?D           P@������������������������       ����i��?4            �T@                           @��O_���?B           ��@������������������������       ���nӹ��?�            `v@������������������������       �tB��3��?S           ��@                           �?����8�?�           X�@                          �1@>caV�?�           X�@                          �0@�:��u��?,            @R@������������������������       �t�@�t�?	             .@������������������������       ���C���?#             M@                          �5@��L���?�           �@������������������������       �m�v�c�?�            �p@������������������������       �(%/���?�            `u@                           @W,{����?6           �~@                          �=@���P�?�            �s@������������������������       ���X��?�            �r@������������������������       ��?             1@                           �?Xo侴 �?o            �e@������������������������       �|���V�?/            �R@������������������������       ��#�U���?@            �X@�t�b�+     h�h4h7K ��h9��R�(KKKK��h��B�       �j@      ?@     �I@      6@      Y@     0�@      A@     D�@      ,@      @     @U@     �P@     �@     `@      0@     �o@      c@      ;@     �D@      2@      U@      @      >@     ��@      &@       @      R@     �J@     �|@     �v@      .@     �i@     @T@      1@      @@       @     �G@      l@      .@     pp@      @      �?      A@      :@     �i@     �c@       @     @[@      8@       @      @      �?      &@     �S@       @     �]@                      (@      "@      O@     �I@       @      B@      .@              �?      �?      @     �G@      �?      N@                      @      @      7@      .@       @      1@      "@       @      @              @      ?@      �?     �M@                       @      @     �C@      B@              3@     �L@      .@      9@      @      B@     `b@      *@      b@      @      �?      6@      1@      b@     �Z@      @     @R@     �L@      .@      9@      @      B@     �a@      $@     @`@      @      �?      6@      1@     �`@     @W@      @     �N@                                              @      @      ,@       @                              &@      ,@              (@      R@      $@      "@      $@     �B@     �p@      .@     �{@      @      �?      C@      ;@     �o@      j@      @     @X@      <@      @       @      @      @     @Z@      @      i@      @              @      "@     �[@     @P@      @      6@      <@      @       @      @      @     �V@      @      e@      @              @      @      X@      J@      @      5@              �?               @      �?      ,@              ?@                               @      .@      *@       @      �?      F@      @      @      @      >@     �d@       @      n@      �?      �?      ?@      2@     �a@      b@       @     �R@      :@      @       @      �?      *@      O@      �?     @W@      �?              @      "@     �Q@      H@              6@      2@       @      @       @      1@      Z@      @     `b@              �?      8@      "@     @R@      X@       @     �J@      N@      @      $@      @      0@     �j@      @      y@      @       @      *@      *@     �n@     �`@      �?     �H@      F@      �?      "@      @      "@     �\@      @     �n@      @       @      @      $@     �]@     @T@      �?      A@       @              �?               @      2@              ,@                      �?      @      ,@      "@               @                                      �?       @                                      �?       @       @      @              @       @              �?              �?      0@              ,@                               @      (@      @              @      E@      �?       @      @      @     @X@      @     �l@      @       @      @      @      Z@      R@      �?      :@      7@      �?      @      @      @     �C@      �?     �X@      �?      �?      @              A@     �C@              0@      3@              @              @      M@       @     �`@       @      �?              @     �Q@     �@@      �?      $@      0@      @      �?      �?      @     �X@      �?     �c@                       @      @     �_@      K@              .@      &@              �?      �?      @     �H@             �\@                      @              U@      A@              $@      &@              �?      �?      @      H@             �Y@                      @             �T@      A@              $@                                       @      �?              (@                                       @                              @      @                      �?      I@      �?      E@                       @      @      E@      4@              @       @       @                      �?      8@      �?      3@                      �?      @      *@      @              @      @      �?                              :@              7@                      �?              =@      ,@               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��OrhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @f�{U��?�	           ��@       	                     �?��4��?�           �@                           �?�m�Ӥ�??           ��@                           �??B��;T�?E           �@������������������������       �gA
����?P            �_@������������������������       �oFl��4�?�           (�@                          �0@�T��|��?�           ��@������������������������       ��u�)�?$            �H@������������������������       �DeGٴ��?�           ��@
                           @��qh��?�           `�@                          �2@�.-3+�?~           ��@������������������������       �дE�7�?{            @j@������������������������       ��k�����?            z@                          �:@x�-�?$             M@������������������������       �t�<�
�?             C@������������������������       ��z�G��?             4@                           �?l[��I�?�           D�@                          @A@rF�CY�?�           ��@                           �?f�\��?�           ��@������������������������       �3̫���?�            `o@������������������������       �[����?�            py@������������������������       �޾�z�<�?             *@                           �?|ϛ̼�?            {@                          �2@h�����?�             l@������������������������       ���B����?&             J@������������������������       �X�j�F�?h            �e@                           @��\��?�            @j@������������������������       �*x9/'�?G             \@������������������������       �`�qT��?<            �X@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @i@      ?@     �F@      <@     �\@     ��@     �E@      �@      0@      &@     �V@     �N@     �@     �@      1@     �n@     `d@      :@      >@      7@     @W@     @~@      B@     ��@      ,@      @     @S@      I@     H�@     �v@      0@      i@     �[@      2@      5@      5@     �K@     �x@      9@     ��@      $@             �I@      <@     �y@     �p@       @     �a@      I@      $@      3@       @     �@@     `f@      *@     @h@      @              8@      ,@     �e@     �\@      �?     �W@      @       @      @      @      $@      "@       @     �C@                      "@      �?      5@      (@              "@     �F@       @      0@      @      7@     @e@      &@     `c@      @              .@      *@      c@     �Y@      �?     @U@      N@       @       @      *@      6@     �j@      (@     0w@      @              ;@      ,@      n@     �b@      @     �G@       @                                      $@              @                       @      �?      1@      "@              @      M@       @       @      *@      6@     �i@      (@     �v@      @              9@      *@     �k@     �a@      @      F@     �J@       @      "@       @      C@     �V@      &@     @a@      @      @      :@      6@      [@      Y@       @      N@      J@       @      @       @      C@     �T@      &@     �\@      @      @      6@      6@     �Y@     �U@       @     �M@      8@      @       @               @     �A@      @      C@              �?      &@       @      8@      1@      @      <@      <@      @      @       @      >@     �G@      @     @S@      @      @      &@      ,@     �S@     @Q@       @      ?@      �?               @                       @              7@                      @              @      ,@              �?                       @                      @               @                      @              @      *@                      �?                                       @              .@                                              �?              �?     �C@      @      .@      @      6@     @g@      @     x@       @      @      ,@      &@      k@     `b@      �?     �F@      ;@      �?      *@      @      2@     �]@      �?     �m@       @      @      "@      @     �Z@     �U@      �?     �A@      :@      �?      *@      @      2@     �]@      �?     @l@       @      @      "@      @     @Z@     �U@      �?     �A@      (@      �?       @              (@      H@             �Q@       @       @      @      @     �B@      B@      �?      (@      ,@              @      @      @     �Q@      �?     `c@               @      @      @      Q@     �I@              7@      �?                                                      $@                                       @                              (@      @       @      �?      @     �P@      @     �b@                      @      @     �[@      N@              $@      @      @      �?      �?      @      ?@      @     �Q@                      @      @     �J@      ?@              "@      �?                      �?              @      �?      "@                       @       @      7@      @              @      @      @      �?              @      :@      @      O@                       @       @      >@      :@              @      @      �?      �?                      B@             �S@                      �?             �L@      =@              �?      @              �?                      2@              C@                                     �C@      *@                      @      �?                              2@              D@                      �?              2@      0@              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJM�}hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�*��n�?�	           ��@       	                   �1@�z>�!1�?N           $�@                            �?N�V���?�            Pr@                           @n(�9W��?p            �e@������������������������       ��A��?X            `a@������������������������       �y�N����?            �@@                           �?�h����?S            @^@������������������������       �	6c����?             1@������������������������       �{�<p��?H             Z@
                          �;@G�R6Z��?�           ��@                           @�I�h��?!           ��@������������������������       ���Fp�?           0�@������������������������       �:P��P��?           �{@                           @�GIl�p�?j            �d@������������������������       ��H�S�?U            ``@������������������������       �4�2%ޑ�?            �A@                          �;@���6��?y            �@                           �?�8���?�           4�@                          �5@��b�= �?�             s@������������������������       ���8���?{            �g@������������������������       �|/}* ��?M            @]@                            @�ު�(��?           l�@������������������������       �H6jF�?�           L�@������������������������       �4��d��?+           �|@                           @�i�b<�?�            `n@                           @/}�\.�?            @h@������������������������       ��F�h��?n            @e@������������������������       ��8��8��?             8@                           @D>�@A�?#            �H@������������������������       �=[y���?             1@������������������������       �     ��?             @@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        j@     �@@      E@      @@     �Z@     (�@     �E@     D�@      2@       @     �R@     �J@     X�@     ��@      6@      o@     �Z@      1@      @@      3@      Q@     �q@      2@     @{@      ,@      @      @@      <@     �r@      n@      &@      `@      9@      �?      @      �?      1@      G@      @     �C@      @      �?      @      "@      G@     �G@      @     �B@      *@              @      �?      $@      6@      @      :@      @      �?       @       @      >@     �A@       @      ,@      (@              @      �?      @      .@      @      .@      @               @       @      <@      @@       @      "@      �?                              @      @              &@              �?                       @      @              @      (@      �?      �?              @      8@       @      *@                       @      @      0@      (@      �?      7@                                      @       @              �?                              �?              @              @      (@      �?      �?              @      6@       @      (@                       @      @      0@      "@      �?      0@     �T@      0@      9@      2@     �I@     �m@      &@     �x@      &@      @      <@      3@     `o@     @h@       @      W@     �P@      *@      5@      2@     �F@     @l@      &@      u@      $@      @      8@      0@      k@      g@       @     �S@     �A@      @      2@      ,@     �@@     �c@      @      n@      @       @      .@      @     �b@     �[@      �?     �D@      @@      $@      @      @      (@     �P@      @      X@      @       @      "@      "@     �P@     �R@      @      C@      .@      @      @              @      &@             �N@      �?              @      @     �A@      $@              *@      (@      @       @              @      $@              K@      �?              @      @      2@       @              (@      @               @               @      �?              @                                      1@       @              �?     @Y@      0@      $@      *@      C@     �t@      9@     �@      @      @      E@      9@      z@      r@      &@     �]@     @X@      *@      $@      &@     �@@     �p@      7@     �@       @      �?     �C@      7@      w@     pq@      $@     @[@      *@              @      �?      @      @@      @     �V@                      @      �?     �P@     �K@       @      <@      (@              @      �?      @      3@       @     �J@                      �?              J@      ;@       @      *@      �?                              @      *@       @     �B@                      @      �?      ,@      <@              .@      U@      *@      @      $@      :@     �m@      3@     @�@       @      �?     �A@      6@      s@      l@       @     @T@     �P@      (@      @      @      6@      f@      2@     �v@      �?      �?      ?@      0@      h@     @g@      @     @Q@      1@      �?      @      @      @     �O@      �?     �g@      �?              @      @     �[@      C@       @      (@      @      @               @      @     �M@       @     �V@       @       @      @       @      H@      "@      �?      $@      @      @                      @     �G@       @      S@               @      @      �?      ?@      "@      �?      $@      @      @                      @     �E@       @      N@               @       @      �?      =@       @      �?      $@                                              @              0@                      �?               @      �?                                               @              (@              .@       @                      �?      1@                                                                       @              @                              �?      "@                                                       @              $@              $@       @                               @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJU/{hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx                              @��ڍy��?�	           ��@       	                   �0@�k����?�           ��@                           @�X<g/�?p            `f@                            �?h ����?O            @_@������������������������       ���X��?!             L@������������������������       �I� ��?.            @Q@                            �?/
k��?!             K@������������������������       ��-����?            �B@������������������������       �/k��\�?             1@
                           �?Yf�}��?p           :�@                          �=@�0J5y�?�           ��@������������������������       �h$�H��?�           �@������������������������       ��:�^���?            �C@                            �?`�u���?�           ��@������������������������       �
wԳ%C�?f           ��@������������������������       ��jp?�?J           X�@                          �@@��jʫ��?�           �@                           @f�����?�           ��@                           �?J��f^��?=           �@������������������������       ��$����?�             p@������������������������       �    ���?�             p@                          �0@���J1��?�           �@������������������������       ��?�0�!�?
             1@������������������������       �S�n0��?v           ��@������������������������       ���k���?             6@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        m@      ;@     �D@      <@     �\@     ��@      @@     ؑ@      1@      @     �T@     �N@      �@     �}@      4@     �p@     �f@      6@      >@      :@     @W@     �}@      :@     ��@      *@      @     �Q@     �K@      }@     `u@      4@     �k@      "@      �?      �?      �?      @     �@@      @      7@      �?       @      @       @      @@     �E@              $@      @      �?      �?      �?      @      :@      @       @                      @       @      ;@      @@              @                              �?      @      &@      @      �?                                      1@      3@              �?      @      �?      �?              �?      .@              @                      @       @      $@      *@              @      @                               @      @      �?      .@      �?       @                      @      &@              @      @                               @      @              .@      �?                              @      @              @      �?                                      @      �?                       @                      �?      @               @     �e@      5@      =@      9@     �U@     �{@      6@     ȅ@      (@       @     �P@     �G@      {@     �r@      4@     �j@      T@      (@      :@      (@     �E@      j@      "@     �p@      @      �?     �A@      =@     �e@      ^@      &@      V@      T@      (@      :@      (@     �D@     �i@      "@     �n@      @      �?     �A@      =@     �e@     @\@      &@     �T@                                       @       @              5@                                       @      @              @      W@      "@      @      *@      F@     `m@      *@      {@      @      �?      ?@      2@     @p@     `f@      "@     @_@     �@@      @              @      @     �Y@      @     �h@       @              &@      @     �Z@     �M@       @      4@     �M@      @      @      @      C@     �`@      "@      m@      @      �?      4@      *@     @c@      ^@      @     @Z@     �I@      @      &@       @      5@     `g@      @     `z@      @       @      (@      @     @n@     @`@              F@     �H@      @      &@       @      5@     `g@      @     Py@      @       @      (@      @     �m@     @`@              F@      2@      �?      $@      �?      "@     �O@      �?     �f@      �?      �?       @       @     �`@     �M@              ;@      "@      �?      @              @     �A@      �?     �T@      �?              @              M@     �@@              3@      "@              @      �?      @      <@             �X@              �?      �?       @     �R@      :@               @      ?@      @      �?      �?      (@      _@      @      l@      @      �?      @      @     �Z@     �Q@              1@      @                               @               @      �?                                      @      �?              @      <@      @      �?      �?      $@      _@      @     �k@      @      �?      @      @      Z@     �Q@              (@       @                                                      1@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJI�dhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @c�+RB��?�	           ��@       	                   �?@C�},��?�           ��@                            �?"��0*�?�            �@                           �?ZP����?           ��@������������������������       ���ߨ�C�?C           H�@������������������������       ������?�           h�@                          �2@�;�ܢ��?�           h�@������������������������       ��'9��?�            @h@������������������������       �a�Y��?8           �~@
                           @��.��T�?*            �P@                           @��%�D��?            �K@������������������������       ����*���?            �@@������������������������       ����J�?             6@������������������������       ����#���?             &@                          �2@xmn5��?�           ܑ@                          �1@����-�?�            �q@                           �?��a!�z�?Z            �`@������������������������       �l-0]V�?            �H@������������������������       �"�]6a��?>            �T@                           �?�k(���?\             c@������������������������       �P"�3[z�?&            �O@������������������������       �x���H�?6            @V@                          �=@�[M A��?           ؊@                           @�������?�           x�@������������������������       �T���?�           ��@������������������������       �ވ��\�?@            �W@                           @b_j���?1             S@������������������������       �v	��H}�?+            @Q@������������������������       �������?             @�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `i@      <@      I@      0@     �Z@     ��@      ?@     4�@      0@      @     �T@     @Q@      �@     h�@      8@     �o@     �b@      7@     �C@      ,@     @U@     �|@      5@     ��@      (@      @     �Q@     �K@     �@      y@      5@     `j@     `b@      7@     �C@      ,@     @U@     �|@      5@     ��@      &@      @     �Q@      J@      @     `x@      4@      j@     @[@      ,@      =@      "@      J@     @v@      1@     ��@      @      �?      I@      A@     Px@      q@      *@     �`@     �M@      @      8@      @      >@      g@      @     �g@      @      �?      9@      6@     �e@     �Z@      "@      O@      I@      "@      @      @      6@     `e@      &@     �u@      @              9@      (@      k@     �d@      @     �Q@      C@      "@      $@      @     �@@     @Y@      @      `@      @      @      5@      2@     @[@     �]@      @      S@      (@       @       @      �?      @      ?@      @     �@@              �?      &@      @      .@      E@      @      6@      :@      @       @      @      ;@     �Q@             �W@      @      @      $@      &@     �W@      S@       @      K@       @                                      @              >@      �?                      @      "@      (@      �?       @                                              @              <@                               @      @      $@      �?       @                                              @              5@                                      @              �?       @                                                              @                               @      @      $@                       @                                      �?               @      �?                      �?       @       @                      K@      @      &@       @      6@      e@      $@     �y@      @              &@      ,@     �p@     �^@      @     �D@      "@              @       @      @      G@       @     �T@                      @      @     @U@      9@              (@      @                              @      7@       @     �D@                      �?      @      @@      .@              @      @                                      @              5@                                      .@      @                      @                              @      2@       @      4@                      �?      @      1@      $@              @      @              @       @      @      7@              E@                      @             �J@      $@               @                       @      �?              (@              3@                                      7@      @              @      @               @      �?      @      &@              7@                      @              >@      @              @     �F@      @      @              .@     �^@       @     `t@      @              @      "@     �f@     �X@      @      =@      D@      @      @              (@     �\@       @     �r@      @              @      "@      c@     �X@              =@      C@       @      @              $@     �X@       @     �p@      @              @       @      a@      V@              4@       @      @       @               @      0@              >@                      @      �?      0@      $@              "@      @                              @      "@              ;@      �?                              <@              @              @                               @       @              7@                                      <@              @                                              �?      �?              @      �?                                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ.�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?��E�qw�?�	           ��@       	                   �:@SBJ��/�?Y           ��@                           @�P_A�?�?�           �@                          �8@�q�$ t�?�           ��@������������������������       �����=t�?�           ��@������������������������       ���^���?<            �W@                            @NN����?�           ��@������������������������       �ly@X<+�?�           ��@������������������������       ���Ά��?U             `@
                            �?�A�����?�             m@                           @�mO1��?$            �I@������������������������       ��|Ӭ��?            �A@������������������������       �     @�?             0@                          �<@�1��!�?{            �f@������������������������       ��W	��?=            @V@������������������������       ��hS<��?>            @W@                          �<@��}?���?r           :�@                           @�crT���?�           �@                            @уm�ϥ�?,           ��@������������������������       ���>�:�?�           ؃@������������������������       ������?�            `k@                           @�a/��?�           ��@������������������������       ���?9R��?�           Є@������������������������       �&��55�?&           `}@                           �?��a �?}            �j@                          �?@���(\��?             D@������������������������       ��0�*�?             9@������������������������       �����2�?             .@                           @�7.��?f            �e@������������������������       �c�O{�?;            �X@������������������������       �lO���?+             S@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      A@      J@      6@      ]@     @�@      6@     `�@      .@      *@      Q@      Q@     ��@     �~@      .@     `m@      \@      7@      A@      ,@     @S@     �t@      (@     �y@       @      "@      <@      A@     �q@     `i@      @     @^@     @W@      0@      =@      *@     �R@      s@      "@     @t@      @      "@      9@      A@     �o@     `f@      @      Y@     �K@      $@      3@      @     �C@     ``@      @     �b@      @       @       @      "@     @Z@     �W@      �?      J@      G@      $@      3@      @     �B@     @Y@      @     �a@       @       @      @      "@     �V@     @R@      �?     �F@      "@                      �?       @      >@               @      �?               @              ,@      5@              @      C@      @      $@       @     �A@     �e@      @     �e@       @      @      1@      9@     �b@     @U@      @      H@     �@@      @      $@      @      @@     �c@       @      `@       @      @      (@      9@     �\@     @S@      @      F@      @       @               @      @      3@      �?     �F@                      @             �A@       @              @      3@      @      @      �?      @      8@      @      V@      @              @              ?@      8@      �?      5@                              �?      �?      @       @      9@                       @              @      @              @                              �?      �?      @       @      1@                       @              @                      @                                               @               @                                              @              �?      3@      @      @               @      3@      �?     �O@      @              �?              :@      3@      �?      0@      @      @      @                      $@      �?      :@       @                              .@       @              &@      *@               @               @      "@             �B@      �?              �?              &@      &@      �?      @     �W@      &@      2@       @     �C@     �w@      $@     ��@      @      @      D@      A@     |@     �q@      $@     �\@      W@      &@      2@       @     �B@     �t@      "@     ��@       @      @      B@      >@     �y@     q@      $@     �[@     �G@       @      @      @      2@     �^@      �?     �p@                      "@      *@     �i@      Y@      @      I@     �D@       @      @      @      1@     �Y@      �?     �e@                      @      &@      c@     @R@      @      E@      @              �?       @      �?      5@              X@                       @       @     �J@      ;@               @     �F@      "@      &@      @      3@      j@       @      u@       @      @      ;@      1@     �i@     �e@      @      N@      :@      @      &@       @      &@      _@       @      h@       @       @       @      &@     @b@     �W@       @      <@      3@      @              �?       @     @U@      @      b@              �?      3@      @     �N@     �S@      @      @@       @                               @      I@      �?     �W@      @      �?      @      @      B@      (@              @      �?                              �?      ,@              ,@      @                      @      �?      �?              �?      �?                                      *@              @                               @      �?      �?              �?                                      �?      �?               @      @                      �?                                      �?                              �?      B@      �?      T@      �?      �?      @      �?     �A@      &@              @      �?                              �?      *@      �?     �J@      �?      �?      @              2@      @              @                                              7@              ;@                              �?      1@       @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��O1hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@Ҁ�s�q�?�	           ��@       	                     @�;�\��?�           �@                            �?�B����?-           ��@                           !@��Z��?�           ��@������������������������       ��TD}�?�           4�@������������������������       ����,�?
             3@                          �7@�����?�           ��@������������������������       ������?D           0@������������������������       �     ��?N             `@
                          �2@q����?^           ��@                           �?|L�]��?�            0r@������������������������       ���T�f�?D            �\@������������������������       ��4_�g��?s             f@                           �?}��K��?�           p�@������������������������       ���C�̷�?t            @f@������������������������       �𵰁���?3           �}@                          �@@j;����?           P|@                           @��2����?           @z@                          @@@%w��&\�?�            �v@������������������������       �r�h��?�            �t@������������������������       ��^v�]�?            �B@                           �?_�#���?!             K@������������������������       �     @�?             0@������������������������       �8�ZY�?             C@                            �?����D��?            �@@������������������������       �*;L]n�?             .@                           @)O���?             2@������������������������       �ףp=
��?             $@������������������������       �      �?              @�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �e@      <@      G@      8@     �Z@     �@     �F@     �@      $@      @     �R@      P@     Ȉ@     h�@      9@      m@     @c@      9@      E@      6@     �W@      �@     �D@     ��@      @      �?     �O@     �N@     0�@     �~@      .@     �j@      ]@      0@      B@      2@     �R@     �{@      B@     ��@      @      �?     �I@      K@     @     Pw@      .@     �g@     �S@      @      =@      *@      J@     `v@      :@     @~@                      ?@      ?@     Px@     Pp@      @     @^@     �S@      @      =@      *@      H@      v@      6@     @~@                      ?@      ?@     0x@     0p@      @     @^@      �?                              @      @      @                                               @       @                     �B@      "@      @      @      7@     �U@      $@      [@      @      �?      4@      7@      [@      \@       @     �P@      >@       @      @      @      .@     �Q@      $@     @S@      @      �?      2@      6@     �S@      X@       @      I@      @      �?              �?       @      .@              ?@                       @      �?      =@      0@              1@      C@      "@      @      @      3@     �d@      @     t@       @              (@      @     �j@     �]@              :@      (@       @       @      @      "@      I@             �R@                      @      @     �S@      C@              .@      @               @      �?              ,@              >@                                      F@      ,@              @      @       @               @      "@      B@              F@                      @      @     �A@      8@              $@      :@      @      @      �?      $@     �\@      @     �n@       @              "@      @     �`@     @T@              &@      "@      @                      @     �B@      @     �L@                      @              <@      9@              @      1@      @      @      �?      @     @S@       @     �g@       @              @      @     �Z@      L@              @      5@      @      @       @      (@     �N@      @     �f@      @      @      &@      @     �T@     �@@      $@      2@      1@      @      @       @      (@     �M@      @     @e@      @      @      &@      @     @S@      6@      $@      2@      1@      @      @       @      (@     �J@      @     �a@      @      @      $@      @     �O@      5@      $@      0@      0@      @      @       @      "@     �H@      �?     �_@      @              $@      @     �O@      3@      @      ,@      �?                              @      @      @      *@       @      @                               @      @       @                                              @              >@                      �?              ,@      �?               @                                                              @                                      @                       @                                              @              7@                      �?              @      �?                      @                                       @              $@                                      @      &@                                                               @               @                                      �?      $@                      @                                                       @                                      @      �?                      @                                                      @                                       @                              �?                                                      @                                      @      �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJRpTuhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @Y��	۪�?�	           ��@       	                    @���|q�?�           �@                           �?j�����?.           ��@                            �?�.�t�h�?|           ��@������������������������       ���^���?!           }@������������������������       ����i;�?[            `a@                           �?��]*#o�?�           8�@������������������������       �� ݫjb�?           �{@������������������������       ��{��Q�?�            �p@
                          �<@��)V`�?�           ��@                           �?�F�B�?�           �@������������������������       ��y1��?�           p�@������������������������       ��h��l��?�           `�@                           @�K�S��?E            @\@������������������������       ����:��?9            �W@������������������������       ��.�s�?             3@                          �2@o�2�@�?�           �@                           @�B�K�T�?�            �o@                           @U��;F��?�             k@������������������������       �     ��?W             `@������������������������       �;n,�R�?5             V@                           @^����T�?            �C@������������������������       ���-�?             =@������������������������       �p=
ףp�?             $@                           �?Z�P�?           ��@                           �?���i�E�?�            `x@������������������������       �;�J��?�            �l@������������������������       �)�c#U:�?d            @d@                          �@@3�f���?           `{@������������������������       �VD��X��?           �z@������������������������       ��g���e�?             &@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `k@      B@     �B@      :@     �^@     ��@     �@@     ��@      4@      @      R@      Q@     x�@     p@      0@     �p@     �e@      <@      <@      8@      X@     `~@      ?@     ��@      1@      @     �O@     �L@     0�@     pv@      ,@     �l@     �U@      (@      .@      2@      O@     �l@      $@     �t@      @              4@      :@     �p@     @^@      @     �[@     �B@      @      $@      (@     �@@     �]@      @     �a@      @              .@      0@     �V@     �O@       @      I@      <@      �?      "@      "@      5@     @X@      @     @^@      @              *@      @      S@     �G@       @      ;@      "@      @      �?      @      (@      6@              5@       @               @      "@      .@      0@              7@     �H@      @      @      @      =@     �[@      @     @g@       @              @      $@     �e@      M@       @     �N@      >@      �?      @      @      1@     @T@             �Z@       @               @      @     �[@     �B@             �D@      3@      @      �?       @      (@      =@      @     �S@                      @      @     @P@      5@       @      4@     @V@      0@      *@      @      A@     p@      5@     @w@      $@      @     �E@      ?@     �o@     �m@      $@     �]@      V@      0@      *@      @     �@@     `m@      5@     `t@      $@      @      D@      <@     �l@     �l@      $@     �\@      E@      "@      "@       @      1@     �]@      $@     @^@      @      @      ,@      *@     �X@     @X@      @      M@      G@      @      @      @      0@     @]@      &@     �i@      @       @      :@      .@     @`@     ``@      @      L@      �?                              �?      6@              G@                      @      @      7@      $@              @      �?                              �?      *@              F@                      @      @      2@      @              @                                              "@               @                                      @      @                      F@       @      "@       @      ;@      g@       @     �v@      @      �?      "@      &@      m@      b@       @      C@      "@      �?      �?      �?      @     �C@              R@                       @      �?     �Q@      C@              0@      "@              �?      �?       @      ?@             �M@                      �?              Q@      >@              ,@       @              �?      �?       @      5@              @@                      �?              >@      :@              (@      @                                      $@              ;@                                      C@      @               @              �?                       @       @              *@                      �?      �?      @       @               @              �?                       @      @              @                              �?      @       @               @                                               @              @                      �?                                             �A@      @       @      �?      7@      b@       @     `r@      @      �?      @      $@     @d@     �Z@       @      6@      <@      @      @              2@      Q@      �?     @\@       @      �?      @      @     �R@     �K@      �?      (@      8@      �?      @              @     �B@             �K@       @      �?       @      @      H@      B@      �?       @      @      @      �?              (@      ?@      �?      M@                       @      �?      :@      3@              @      @      @      @      �?      @     @S@      �?     �f@      �?              @      @      V@     �I@      �?      $@      @      @      @      �?      @     @S@      �?     @f@      �?              @      @     @T@     �I@      �?      $@      �?                                                      @                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJuy�MhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @�&B�k�?�	           ��@       	                   �0@�y�����?�           ��@                           �?@.d�]@�?p             f@                           @��L�n��??            @Y@������������������������       �`ל�<��?            �H@������������������������       ���
ц��?!             J@                           @��UH��?1             S@������������������������       ���%�L�?            �D@������������������������       ����:��?            �A@
                          �1@!��]���?�           H�@                            �?1]$�?�             t@������������������������       ���8u���?D            �Y@������������������������       �ԭ�h�G�?�            �k@                            �?��]��?�           ġ@������������������������       ��*�gA�?^           P�@������������������������       �fP5���?\           p�@                           �?��M4���?�           Б@                           @�l�)M�?/           P~@                          �9@��i>�?�            �m@������������������������       �$�?���?x            �h@������������������������       �
ףp=
�?             D@                           @��tS��?�            �n@������������������������       �]�v���?y            @g@������������������������       �<+	���?"             N@                          �0@�ʽ��?�           x�@������������������������       �r�q��?             8@                          �2@.c����?z           ��@������������������������       �:�uf��?\             b@������������������������       �vG�MGY�?           `~@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@      8@      @@      8@     @Z@     P�@      @@     ��@      4@      @     �R@     @P@     ��@     �@      7@      p@     �b@      .@      7@      6@     @U@     �}@      ;@     p�@      0@      @      P@      L@     `@     Px@      6@     �i@      @      �?       @      �?       @      >@       @      5@      @              @      @     �A@      D@      �?      2@       @      �?       @      �?       @      (@       @      *@      @               @      @      ,@      7@      �?      (@                       @                       @      �?      @                      �?      @      $@      (@      �?      @       @      �?              �?       @      @      �?      @      @              �?              @      &@               @       @                                      2@               @                       @       @      5@      1@              @      �?                                      @              �?                               @      1@      &@              @      �?                                      *@              @                       @              @      @               @     @b@      ,@      5@      5@     @S@     �{@      9@     ȅ@      (@      @      N@      I@     0}@     �u@      5@     �g@      9@      �?      @              ,@     �P@      @      T@                      "@      @      B@      H@      @      5@      &@               @              @      3@       @     �A@                               @      @      &@              @      ,@      �?       @               @      H@      @     �F@                      "@      @      =@     �B@      @      ,@     @^@      *@      1@      5@     �O@     �w@      3@     H�@      (@      @     �I@      F@     �z@     �r@      0@      e@      U@      @      &@      2@      D@     �s@      *@     �@      @             �@@      7@     �t@     �j@      "@     @_@     �B@      @      @      @      7@      N@      @     �Y@      @      @      2@      5@     @X@     �U@      @     �E@     �I@      "@      "@       @      4@      f@      @     �y@      @              &@      "@      p@     @^@      �?     �I@      >@      @      @      �?      ,@     �T@      @      a@       @              $@      @     �Z@      L@      �?      ;@      ,@              @      �?      @      @@      �?      M@      �?              $@      �?     �P@      =@              ,@      ,@              @      �?      @      >@      �?      E@                      $@              J@      :@              ,@                      �?              �?       @              0@      �?                      �?      .@      @                      0@      @                       @      I@       @     �S@      �?                      @     �C@      ;@      �?      *@      0@      @                      @     �B@      �?     �H@      �?                      @      A@      7@      �?      "@                                      @      *@      �?      >@                                      @      @              @      5@      @      @      �?      @     �W@       @     0q@       @              �?      @      c@     @P@              8@                                              @              0@                                      �?       @               @      5@      @      @      �?      @      W@       @     0p@       @              �?      @     �b@     �O@              6@       @              �?               @      2@              G@                              �?     �I@      *@              @      *@      @      @      �?      @     �R@       @     �j@       @              �?      @      Y@      I@              1@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ^�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@H�{����?�	           ��@       	                     @�ݞl`��?�           0�@                            �?���sB/�?6           ��@                            �?�K*��?�           ��@������������������������       ��P���_�?>           p�@������������������������       �g4f�?u           <�@                           �?D����?�           ��@������������������������       �lA����?�            p@������������������������       �	������?�            0u@
                           �?�X/p�C�?R           8�@                          �2@��իF�?M           Ȁ@������������������������       �"�r���?R            �`@������������������������       ��O����?�            @y@                           �?n�3�a�?           �z@������������������������       ��S�r
�?�             l@������������������������       ���:連�?~            �i@                          �@@>���^�?           {@                           �?̋U��,�?�            �x@                           @6
=Ȕ�?i             e@������������������������       �
��d~�?P            @`@������������������������       �ޭg_{�?            �C@                           @xn�M;��?�            @l@������������������������       �� �N0�?z            �g@������������������������       ���Hx��?             B@                           @@�'�@��?             C@                           �?�i��F�?             =@������������������������       ��u]�u]�?             5@������������������������       �      �?              @������������������������       ���"e���?             "@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@      1@     �H@     �A@     �]@     ��@      >@     ��@      .@      &@     �U@     �R@     ؆@     �@      8@      p@     @f@      1@      G@     �@@     �Z@     ��@      ;@     p�@      &@      "@      T@     �Q@     Є@     �}@      4@     �m@     �b@      $@     �A@      <@      V@     px@      4@      �@      $@       @      P@     �K@     �|@     �v@      4@      i@     @]@      @      8@      6@     �O@     t@      0@      �@      @      @     �C@      <@     Pv@      o@      0@      a@     �K@      @      @      0@      ,@     �b@       @     �o@       @              0@      &@     �c@     �`@      @      G@      O@      @      1@      @     �H@     `e@       @      p@      @      @      7@      1@     �h@     @]@      $@     �V@     �@@      @      &@      @      9@     �Q@      @      Y@      @       @      9@      ;@     �Y@     �\@      @      P@      *@       @      @      @      ,@      :@       @     �F@      @      �?      @      ,@      F@      H@      @      ;@      4@       @      @      @      &@      F@       @     �K@      �?      �?      4@      *@      M@     �P@             �B@      <@      @      &@      @      2@     �e@      @     �t@      �?      �?      0@      .@     �i@     �[@             �C@      ,@       @      "@      @      $@     �X@      @     �g@      �?      �?      @      (@      X@      Q@              5@       @              @      @      @      2@             �C@                       @      @      8@      ?@              @      (@       @      @      �?      @      T@      @     �b@      �?      �?      @       @      R@     �B@              2@      ,@      @       @      �?       @     �R@      @     �a@                      "@      @     �[@      E@              2@       @       @              �?      @      F@      @      N@                      "@       @     �J@      6@              ,@      @      @       @               @      >@              T@                              �?      M@      4@              @      7@              @       @      (@      P@      @      g@      @       @      @      @     @P@     �B@      @      3@      5@              @       @      (@     �J@      @     �e@      @       @      @      @      M@      @@      @      2@      2@              @              "@      :@              O@                       @       @      5@      .@              &@      2@              @              "@      6@             �C@                       @       @      2@      &@              @                                              @              7@                                      @      @              @      @                       @      @      ;@      @     �[@      @       @      @      �?     �B@      1@      @      @      @                       @      @      :@      @     �T@      @       @      @      �?      A@      .@      @      @                                              �?              =@                      �?              @       @                       @                                      &@              &@                              �?      @      @              �?       @                                      "@               @                                      @       @              �?       @                                       @              @                                      @                      �?                                              �?              @                                       @       @                                                               @              @                              �?              @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJZ0MmhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?��B����?�	           ��@       	                   �=@�%�'�?H           �@                            @���#�?           ��@                            �?�Z�?�           d�@������������������������       ������2�?0           ȋ@������������������������       ��Hx�U�?�             r@                           @��5$�^�?,            }@������������������������       ��)Hs�?�            �s@������������������������       �`JjԆ��?c            `b@
                           �?��!3�?4            �V@                            �?T`�[k�?!            �J@������������������������       �r�q��?             (@������������������������       �:��d�_�?            �D@                           @)���}�?             C@������������������������       ��nkK�?             7@������������������������       �؂-؂-�?             .@                            @��_�y��?`           �@                           @rG�)$t�?�           ��@                          �4@׃�u	��?�           ̑@������������������������       �*$���?d           h�@������������������������       �,��K�?}           0�@                            �?Ti����?           `{@������������������������       ��0�S�&�?�            �u@������������������������       �'O5��q�?=            �W@                           @<����0�?x           Ђ@                           @ű���?            }@������������������������       ��-
1��?           |@������������������������       ��?�0�!�?             1@                           @����p�?Y             a@������������������������       ���;۝�?P            @]@������������������������       �=�
I��?	             3@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        l@      <@     �C@      6@     @\@     ��@      ?@     �@      7@      @      R@      O@     ��@     ��@      2@     `n@      \@      &@      ;@      *@      P@     �r@      3@      z@      1@      �?     �B@      :@     �q@     �p@      @     �`@     �Y@      &@      ;@      *@     �K@     �r@      3@     0x@      &@      �?     �B@      7@      q@     �o@      @      `@     �R@      $@      .@      &@      D@     �j@      "@     @o@      $@      �?      =@      4@     �g@     �g@      @      [@     �O@      @      ,@       @      <@      d@       @     �i@      @              7@      ,@     �c@      _@      @      R@      (@      @      �?      @      (@     �J@      �?      G@      @      �?      @      @     �@@     �P@       @      B@      ;@      �?      (@       @      .@      U@      $@      a@      �?               @      @     @T@      P@              5@      3@              $@       @      &@     �N@      @     �U@                      @      �?     �N@      E@              0@       @      �?       @              @      7@      @     �I@      �?               @       @      4@      6@              @      $@                              "@      @              ?@      @                      @      $@      *@              @      @                              @      @              2@      @                      @      @                       @                                                              $@                                       @                              @                              @      @               @      @                      @      @                       @      @                               @                      *@                                      @      *@              �?                                       @                      $@                                      @       @                      @                                                      @                                       @      @              �?      \@      1@      (@      "@     �H@     �t@      (@      �@      @      @     �A@      B@     p}@     Pr@      *@     �[@      X@      *@       @       @      A@     �n@      (@     p{@      �?       @      A@      ?@      t@     @m@      (@     �U@     �T@      @      @      @      9@      i@       @     �r@      �?      �?      5@      1@     �l@     `c@      "@     �Q@      G@               @       @      "@     �[@      @     �`@                      $@      $@      X@      W@      @      B@     �B@      @      @      @      0@     �V@      @     �d@      �?      �?      &@      @     �`@     �O@      @      A@      *@      @       @       @      "@     �F@      @     `a@              �?      *@      ,@     �V@     �S@      @      1@       @      @               @      "@     �C@      @     �_@                      &@      $@      Q@     �J@              "@      @               @                      @      �?      *@              �?       @      @      7@      :@      @       @      0@      @      @      �?      .@     �T@              m@      @      �?      �?      @     �b@     �M@      �?      8@      ,@      �?      @      �?      *@     �G@             �g@      @      �?      �?      @      ^@      F@              6@      ,@      �?      @      �?      *@      G@              g@      �?      �?      �?      @     @]@     �E@              3@                                              �?              @      @                      �?      @      �?              @       @      @                       @     �A@              F@                              �?      ?@      .@      �?       @       @      @                       @      =@              D@                              �?      8@      *@      �?       @                                              @              @                                      @       @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�m)hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?m�b�?�	           ��@                            @ouy��?c           |�@                          @@@5���_�?'           l�@                          �=@�jhd�?           �@������������������������       �ޛWe�d�?           ��@������������������������       ���h�C�?             ;@������������������������       ���Q���?
             4@                           @����o�?<            �@	       
                    @�ā��?�            0w@������������������������       ��f��@W�?�            �u@������������������������       ��������?             8@                           @�y�!���?d             b@������������������������       ��^�:|�?9             U@������������������������       �`�4 ը�?+            �N@                           �?�3h
���?Z           Ԡ@                            @
� ��b�?�            �u@                          �0@֍���?�            `n@������������������������       ��zv��?             &@������������������������       ����x۷�?�             m@                           @W�h�+��?B            �Z@������������������������       �2��T��?3            @T@������������������������       �(������?             9@                           !@�n`d��?           4�@                            @�SL˭��?u           �@������������������������       ����XnT�?:           ,�@������������������������       �$�J�9�?;           @������������������������       �$�ɜoB�?
             1@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      6@      C@     �A@     �\@     Ѕ@      @@     đ@      &@      @      R@     @Q@     ��@     �@      &@     �n@     @W@      $@      >@      0@     �R@     �u@      0@     �{@       @      @      B@      >@      r@     @m@      @     �_@      N@      @      6@      0@      L@      n@      .@     �p@       @      @      =@      ;@     �i@      f@      @     �[@      N@      @      6@      0@      L@      n@      .@     Pp@       @      @      =@      ;@      i@     �d@      @     �[@      M@      @      6@      0@     �I@      n@      .@      o@       @      @      =@      ;@     �h@     �d@      @      [@       @                              @                      (@                                      @      �?              @                                              �?              @                                      @      &@                     �@@      @       @              2@      Z@      �?      f@                      @      @     �U@     �L@              0@      @@      @      @              .@     @T@      �?     @^@                              @      M@      F@              @      <@      @      @              .@      S@      �?     @]@                              @      L@     �B@              @      @                                      @              @                                       @      @               @      �?       @       @              @      7@              L@                      @              <@      *@              $@              �?                      �?      &@             �C@                       @              4@      @              @      �?      �?       @               @      (@              1@                      @               @       @              @     @X@      (@       @      3@      D@     v@      0@     ��@      @       @      B@     �C@     P{@     �p@       @     �]@      0@               @       @      "@      F@      @     @Y@                      @      @      P@      O@      @      =@      &@              �?       @      @      <@      @      N@                      @      @     �H@      E@      @      :@      @                                      @                                                       @      �?               @       @              �?       @      @      9@      @      N@                      @      @     �G@     �D@      @      8@      @              �?              @      0@      �?     �D@                                      .@      4@              @      @              �?              @      &@      �?      A@                                      .@      "@              @      �?                              �?      @              @                                              &@                     @T@      (@      @      1@      ?@     Ps@      (@     ��@      @       @      @@      @@     Pw@      j@      @     �V@     @T@      (@      @      1@      ?@     �r@      (@     h�@      @       @      @@      @@     @w@     �i@      @     �V@      Q@      &@      @      *@      =@     �k@      &@     �w@      @      �?      <@      9@     `o@     �d@      @     �S@      *@      �?      �?      @       @     �S@      �?     �j@              �?      @      @     @^@     �D@              &@                                               @              @                                      �?      @                �t�bub�/     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�WhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @{��HT��?�	           ��@       	                     �?#�WYj�?�           ��@                           �?���l��?%           �@                           �?�T�x�9�?H           x�@������������������������       �^䑎���?S            �a@������������������������       �2�j7�?�           �@                           @<z./��?�           �@������������������������       �p^FW4��?�           Є@������������������������       ��y5���?1            ~@
                           �?:�|
H��?�           x�@                           �?m��Š"�?)            @Q@������������������������       ���Jr�?            �@@������������������������       ����[���?             B@                          �;@{��s��?�           P�@������������������������       �"#M���?o           �@������������������������       �؂-؂-�?            �F@                          �;@�ffB0�?�           đ@                           �?twѿ�@�?t           ��@                          �2@���\��?�             s@������������������������       �����W�?D             \@������������������������       ��8��86�?{             h@                           �?ᩴ����?�           �@������������������������       �����<�?�            �q@������������������������       �}�Fػ�?�            �z@                           �?X��$��?Q            �_@                           �?���2���?$            �J@������������������������       �s
^N���?
             ,@������������������������       �ݾ�z�<�?            �C@                          �=@}>���?-            @R@������������������������       ��������?             8@������������������������       �`�a	���?            �H@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      =@     �D@      4@      \@      �@      @@     �@      1@      @     @X@      S@     x�@     (�@      3@     �p@     �c@      6@      ;@      0@      V@     @@      :@      �@      *@       @     @S@      O@     0~@     �x@      2@      k@     �[@      &@      1@      *@     �O@     �x@      4@     ��@      @              E@      ?@     0x@      q@      &@     �a@     �J@      @      ,@      @      G@     �f@      $@     `h@      @              3@      *@      e@     �\@      @     @S@      "@               @       @      "@      0@             �B@                      @      @      A@      1@              @      F@      @      (@      @     �B@     �d@      $@     �c@      @              (@      $@     �`@     @X@      @      R@      M@      @      @      @      1@     �j@      $@     @u@       @              7@      2@     `k@      d@      @     @P@     �@@       @      @      @      "@     �b@      @      h@       @              "@      &@     �^@      S@      @      F@      9@       @              @       @      P@      @     `b@                      ,@      @      X@      U@      @      5@      G@      &@      $@      @      9@     @Z@      @     �a@       @       @     �A@      ?@      X@     �]@      @     �R@      @      @      �?       @       @      @              @      @              @              &@      *@      �?      (@              @      �?              �?      @              @      @                              @      @              @      @                       @      �?      �?              �?                      @               @      "@      �?      @     �E@       @      "@      �?      7@     @Y@      @     �`@       @       @      >@      ?@     @U@     @Z@      @     �O@     �C@       @      "@      �?      7@     @W@      @     @]@       @       @      <@      ?@      S@      Z@      @     �N@      @                                       @              2@                       @              "@      �?      �?       @     �C@      @      ,@      @      8@      f@      @     z@      @       @      4@      ,@     �m@     @_@      �?      H@      ?@      @      *@      @      4@     �d@      @     �u@       @      �?      4@      (@     �j@     �^@              E@      $@      �?      @      �?      @     �E@      @     �U@                      "@      @     �R@      F@              4@      @              @      �?              .@              =@                                      E@      "@              @      @      �?                      @      <@      @     �L@                      "@      @     �@@     �A@              *@      5@      @       @      @      0@     �^@      @     �p@       @      �?      &@      "@     �a@     �S@              6@      $@      @      @              $@     �K@      �?     �U@              �?      @      @      J@      @@              1@      &@       @      @      @      @     �P@       @     `f@       @              @      @      V@      G@              @       @              �?              @      &@             �P@       @      �?               @      5@      @      �?      @      @              �?              @      @              4@       @                       @       @       @      �?      @                                              �?              @                               @      @       @               @      @              �?              @       @              1@       @                              @              �?      @       @                              �?       @              G@              �?                      *@      �?              �?                                              @              .@                                              �?              �?       @                              �?      �?              ?@              �?                      *@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJe/�DhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             @�m�XH��?�	           ��@       	                    �?&a~���?'           ��@                          �1@�~c�iR�?�           ��@                            �?�5��?�             k@������������������������       ����E��?O            @^@������������������������       ��V��?8            �W@                          �:@D�0�	�?x           8�@������������������������       �>�Q,�.�?           ��@������������������������       �u0i����?r            `e@
                           @�W����?(           4�@                            @h+�8B��?�           @�@������������������������       ���x�P��?=            @������������������������       �X�<ݚ�?�             k@                           @6��ݦ�?X           (�@������������������������       �������?N           ؀@������������������������       ���g�_�?
           �z@                            �?�����a�?m           �@                          �;@(a�4(F�?�            @k@                           �?ȿj�MG�?z            `h@������������������������       �x|T
�?/            @R@������������������������       �m�oڑ�?K            �^@������������������������       ��LQ�1	�?             7@                           @e��p��?�           �@                            @ ���?�            �w@������������������������       �e��xp��?�            �t@������������������������       �VUUUU��?             H@                           �?ت���H�?           �z@������������������������       ��Xa����?y            `i@������������������������       ���A�j�?�            �k@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @j@      =@      =@      <@     �`@     �@     �B@     h�@      ,@       @     �Q@     �K@     (�@     P�@      ,@      q@     `c@      :@      4@      :@     @U@     @~@      <@     ��@      &@      �?     �I@      ;@     ��@     �y@      &@     �h@     @S@      6@      *@       @     �D@     �h@      &@     �q@       @      �?      =@      3@     @k@      d@      @     �_@      2@      @      @      �?      @      >@      @      <@      �?              @      @     �B@      ;@      �?     �D@      ,@              @      �?      �?      0@      @      .@      �?               @      @      6@      8@              .@      @      @      �?              @      ,@              *@                      @       @      .@      @      �?      :@     �M@      1@      "@      @      A@     �d@       @     �o@      @      �?      6@      *@     �f@     �`@      @     �U@     �I@      &@      @      @      >@     �a@      @      h@      @      �?      0@      &@     �b@     �]@      @     �R@       @      @       @              @      7@      �?      N@                      @       @     �@@      ,@      �?      &@     �S@      @      @      2@      F@      r@      1@     �@      @              6@       @     �u@     �o@      @     �Q@     �H@      @      @      @      9@     �[@      @     �i@                      @       @      e@      X@       @      ?@     �D@      @      @       @      5@     �T@      @     �]@                      @       @     �[@     @S@       @      7@       @                      @      @      ;@              V@                       @             �L@      3@               @      =@      �?      @      *@      3@     @f@      (@     s@      @              .@      @      f@     �c@      @      D@      6@              �?       @      &@     �X@      $@     �e@       @              @      @     @W@     �R@       @      >@      @      �?      @      @       @     �S@       @     @`@      �?              "@      �?      U@      U@       @      $@     �K@      @      "@       @     �G@      c@      "@     0t@      @      @      4@      <@     @f@     �Z@      @     �R@       @      @              �?      *@      >@              W@                      �?       @      B@      6@      �?      "@       @      @              �?      *@      >@              R@                      �?       @     �@@      6@      �?      "@       @                              @      5@              7@                               @      @      $@              @      @      @              �?      "@      "@             �H@                      �?              :@      (@      �?      @                                                              4@                                      @                             �G@              "@      �?      A@     �^@      "@     �l@      @      @      3@      :@     �a@     @U@       @     @P@      <@              @              ,@      D@      @     �[@      �?      @      (@      4@     �K@      G@       @      ?@      <@              @              ,@      C@      @     @U@      �?      @      &@      4@      E@     �D@       @      >@                                               @              :@                      �?              *@      @              �?      3@              @      �?      4@     �T@       @      ^@       @      �?      @      @     �U@     �C@              A@      *@              @      �?      0@     �A@       @      K@              �?      �?      �?      @@      :@              2@      @               @              @      H@             �P@       @              @      @     �K@      *@              0@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�>7hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?��rI��?�	           ��@       	                    �?Ƿ��@�?9           P�@                           �?��z�YK�?�           ��@                            �?�l�@�s�?9            @W@������������������������       ��ƖJ��?             ?@������������������������       ������?%             O@                          �<@_1d�O�?�           ��@������������������������       �%���-�?o           ��@������������������������       �{9�D�?            �G@
                          �0@؟�4��?v           ��@                            �?�^��T�?              M@������������������������       ��q-�?             *@������������������������       ������?            �F@                           @ ��C7�?V           ��@������������������������       �����O�?�           �@������������������������       ��o<���?�             l@                           @��(�3��?o           j�@                           @G͜���?h           4�@                            @�G����?-           \�@������������������������       �� f`���?(           ؋@������������������������       ��I;Wq�?           �y@                            �?;_�\�?;           `@������������������������       ��+��^��?�            0s@������������������������       �=F��*��?�            `h@                          �?@�ZE�G��?           �z@                            �?k���{��?           �y@������������������������       �]t�E�?9             V@������������������������       ��&����?�            `t@������������������������       ����Q��?             $@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        l@      :@      B@      <@     @\@     �@     �B@     l�@      6@       @     �V@      K@     0�@      @      8@     �o@      [@      ,@      6@      .@     �Q@     �q@      5@     `y@      $@      @      G@      ;@     �r@     �k@      (@      ^@      C@      @      &@      "@     �A@     �`@      @     �b@      @      �?      ;@      (@     `c@     @V@       @     �J@      @              �?              @      @              5@      �?              (@       @      *@      1@              "@      @                              �?      �?              (@                      @              @      @              �?      �?              �?              @      @              "@      �?              @       @      $@      *@               @     �@@      @      $@      "@      >@     �_@      @      `@      @      �?      .@      $@     �a@      R@       @      F@      @@      @      $@      "@      >@      _@      @      Z@      @      �?      (@      $@     �`@     �Q@       @      D@      �?                                       @              9@      �?              @              "@       @              @     �Q@      $@      &@      @      B@     �b@      .@      p@      @      @      3@      .@     �b@     ``@      $@     �P@       @                              �?      @              @                               @      $@      1@               @                                              �?              @                                              @              �?       @                              �?      @              �?                               @      $@      (@              @      O@      $@      &@      @     �A@      b@      .@      o@      @      @      3@      *@     @a@     �\@      $@     �M@      H@      $@      @      @      8@      ]@      .@     �d@      @      @      2@      (@      Z@     @W@      @     �D@      ,@              @       @      &@      =@              U@              �?      �?      �?      A@      5@      @      2@     @]@      (@      ,@      *@      E@     �v@      0@     (�@      (@       @     �F@      ;@     p{@     @q@      (@     �`@     �X@      $@      "@      $@      <@      r@      ,@     ��@       @       @      ;@      9@      v@     @m@      @     @X@     �S@       @      @      @      7@      k@      @     �y@      @       @      @      2@      q@     `c@      @     �S@      P@      @      @      @      1@      d@      @      m@      @              @      ,@     �f@     @]@      @     @P@      .@      �?       @              @      L@       @     `f@       @       @              @     �V@      C@              ,@      3@       @      @      @      @     @R@      @     �f@      @              4@      @     �T@     �S@              2@      (@      �?              @      @      A@      @      _@       @              ,@      @      G@     �F@              *@      @      �?      @              �?     �C@      �?     �L@      �?              @      @      B@      A@              @      3@       @      @      @      ,@     �Q@       @      ]@      @              2@       @     @U@      E@      @      B@      3@       @      @      @      ,@      P@       @      ]@                      2@       @     @U@      E@      @      B@       @      �?                      �?      @      �?      >@                       @              6@      ,@      @      @      1@      �?      @      @      *@      M@      �?     �U@                      0@       @     �O@      <@      @      >@                                              @                      @                                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�hPhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@�����?�	           ��@                            @���Q���?~           *�@                           !@{a�Ţ&�?           ��@                           @��Q��?           ��@������������������������       �^�T��$�?�           $�@������������������������       ����l��?O           �@������������������������       �ݾ�z�<�?             *@                           �?B�{y�?_            �@	       
                    @
�jL�>�?           @z@������������������������       �"�2�Ot�?�            pt@������������������������       �o�׼t�?D            @W@                           @v:�����?N            �@������������������������       �t����?�            py@������������������������       �7|]�4�?O             a@                           @�PO�.��?           @{@                            �?�21N�?�            �v@                          �=@iQJ��>�?>            �W@������������������������       �@�(ݾ��?              J@������������������������       �^b�m�?            �E@                            @����P�?�            �p@������������������������       ����[פ�?`            �b@������������������������       �������?L            @^@                           �?��{���?2            �Q@                           @W3g	�?            �@@������������������������       ��]�`��?
             *@������������������������       �
ףp=
�?             4@                          �=@�<J�L�?            �B@������������������������       �g\�5�?
             *@������������������������       ��q�q�?             8@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        k@      3@      C@      5@     @[@     ��@     �C@     h�@      3@      &@      V@     @P@     ��@     �~@      2@     0p@     @h@      1@     �A@      4@      Y@     ؂@      B@     X�@      0@      "@     �S@      M@     ��@     �|@      0@     @m@     �c@      $@      ;@      .@      V@     P{@      @@     �@      .@      @     @Q@     �H@     `{@     �u@      0@     @h@     �c@      $@      ;@      .@     �T@     0{@      >@     �@      .@      @     @Q@     �H@     `{@     �u@      0@     @h@     �U@       @      3@      $@      I@     @k@      &@     �p@      @       @      3@      =@      k@     �`@      @      U@     �Q@       @       @      @     �@@      k@      3@     @u@      &@      @      I@      4@     �k@     `j@      &@     �[@       @                              @       @       @                                                       @                     �A@      @       @      @      (@     �d@      @     �t@      �?      @      $@      "@     �k@     �\@              D@      8@      @      @      �?       @     @W@      @      Z@              @      @      �?     �V@     �I@              9@      6@      @      @              @     �R@      @     @Q@              @      �?      �?      R@      G@              4@       @                      �?      �?      3@             �A@                      @              3@      @              @      &@       @      @      @      @     @R@      �?      l@      �?              @       @     ``@     �O@              .@      @      �?      @      @      @      J@      �?     �c@      �?              �?       @     �Y@      J@              ,@      @      �?                      �?      5@             �P@                       @              <@      &@              �?      6@       @      @      �?      "@      Q@      @     �e@      @       @      "@      @     �R@      >@       @      9@      2@       @      @              @     �J@      @     �c@      �?       @      "@      @      J@      9@       @      8@      @                              @      @      �?      K@                              �?      1@      @              @      @                              �?      @              8@                                      (@       @              @                                       @      �?      �?      >@                              �?      @      @                      .@       @      @              @      G@       @      Z@      �?       @      "@      @     �A@      4@       @      4@      "@       @      @               @      <@       @      G@                      "@      @      3@      $@      �?      ,@      @                               @      2@              M@      �?       @              �?      0@      $@      �?      @      @                      �?       @      .@              1@       @                              7@      @              �?      @                               @                      "@                                      (@      @              �?      @                                                      @                                      @       @                      �?                               @                      @                                      "@      @              �?                              �?              .@               @       @                              &@                                                      �?               @              @                                      @                                                                      *@               @       @                              @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJJוMhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx         
                     @�0sf ��?�	           ��@       	                    !@�&)�!��?�           ��@                            �?�*[���?�           ��@                            �?ܰx+o��?2           j�@������������������������       ���	k�?�           ,�@������������������������       �}�j�/��?�           ��@                           @�`'<���?�           X�@������������������������       ���9e�c�?�            �q@������������������������       ��S���?�             w@������������������������       ���Q���?
             4@                           �?�i.��?�           ԑ@                           �?��θR�?�           ��@                          �8@IUY�?�            �o@������������������������       �D���@s�?v            `h@������������������������       �JC�ɯ�?*            �L@                          �;@��U���?�            �y@������������������������       �V�J����?�            pv@������������������������       �)ݾ�z��?%             J@                           �?�,O>��?,           �}@                          �4@�Z$���?�            �m@������������������������       ���$��?K            �]@������������������������       ��%�X��?H             ^@                           @6�h$`�?�             n@������������������������       ���`�#�?Y            `b@������������������������       ��V�z^�?@            @W@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @l@      >@      :@      8@     @W@     Ȅ@      @@     x�@      <@      "@     @T@      J@     �@     `@      :@     pp@     `e@      6@      7@      5@     �R@     �}@      :@     P�@      5@       @     �P@      E@     �~@     Px@      9@     �i@     `e@      6@      7@      5@      R@     �|@      8@     @�@      5@       @     �P@      E@     �~@     0x@      9@     �i@     �`@      ,@      "@      2@     �G@     pw@      0@     8�@      1@      �?      G@      8@     �x@     �p@      0@     �a@     �I@       @       @      $@      0@     `g@      $@     �s@       @              3@      &@     �g@     �b@      $@     �H@     �T@      @      @       @      ?@     �g@      @     �p@      "@      �?      ;@      *@     `i@     �]@      @      W@      C@       @      ,@      @      9@      V@       @      `@      @      @      5@      2@     �W@      ^@      "@     @P@      "@      @      @      �?      "@      =@             �P@       @      @      "@      @      H@     �H@      @     �@@      =@      @       @       @      0@     �M@       @     �O@       @      @      (@      *@      G@     �Q@      @      @@                                      @      "@       @       @                                       @       @                     �K@       @      @      @      2@      h@      @     @y@      @      �?      ,@      $@      o@     @\@      �?     �L@      E@      @       @       @       @      ]@      @     �l@      @      �?      @      @     �_@     �S@      �?      ?@      :@      �?                      @      J@       @     @R@      @              �?              B@     �C@              (@      $@                              @     �E@       @     �O@      �?              �?              ;@      ?@              (@      0@      �?                              "@              $@      @                              "@       @                      0@       @       @       @      @      P@      @     �c@       @      �?       @      @     �V@     �C@      �?      3@      0@       @       @       @       @      H@      @     �`@       @               @      @     @U@     �B@      �?      2@                                      �?      0@              :@              �?                      @       @              �?      *@      @      �?      �?      $@     @S@      �?     �e@                      &@      @     �^@     �A@              :@      @       @      �?      �?      "@     �D@      �?     �P@                      $@       @     �L@      2@              8@      @      �?              �?      @      ;@      �?      B@                      @       @      3@      @              (@       @      �?      �?              @      ,@              >@                      @              C@      *@              (@      @      @                      �?      B@             �Z@                      �?      �?     @P@      1@               @      @                              �?      (@              S@                              �?     �F@      @               @      @      @                              8@              ?@                      �?              4@      $@                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�0IhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@�˾�OR�?�	           ��@       	                     @߆��Uo�?�           �@                           @1�R�y��?&           8�@                          �9@��nb��?�           8�@������������������������       ���\��?�           T�@������������������������       �F�E��?N            @^@                          �0@j��*�(�?N           p�@������������������������       ��6�i��?(             N@������������������������       ��[7��?&           ��@
                           �?������?v           ��@                          �9@�ˍL��?�            @s@������������������������       ��*;�?�?�             r@������������������������       ���ӭ�a�?	             2@                           �?�>?2e��?�           ��@������������������������       ��(����?�            �p@������������������������       �$�
��?           �z@                           �?���v��?           �{@                           �?�]����?-            �S@                          �<@�tk~X��?             B@������������������������       �$��Z=;�?             6@������������������������       �
^N��)�?             ,@                           �?e�J���?             E@������������������������       ��q�q�?             (@������������������������       �ϊF��?             >@                           @�^-����?�            �v@                            @��|mV�?�            @t@������������������������       ����/t�?�            �j@������������������������       ���t�h�?G            �[@                           @
oΕ�c�?            �E@������������������������       �fP*L��?             6@������������������������       ���+��?             5@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �f@      >@      ?@      5@     �Y@     x�@      :@     ��@      8@      �?     @Q@     �P@     �@     (�@      0@     �n@     �c@      :@      :@      4@     @W@     �@      9@     �@      1@      �?      L@      P@      �@     �~@      ,@     �l@     �]@      .@      5@      0@      T@     0|@      3@     `�@      ,@      �?     �H@      K@     �{@     Pv@      ,@     `g@     �R@       @      .@       @      N@      r@       @     0z@      @      �?      7@      B@     @r@     `h@      @     @\@      P@      @      .@      @      M@     0q@      @      x@      @      �?      6@      B@      p@      g@      @     @[@      &@       @              @       @      *@      @     �@@       @              �?              B@      &@              @      F@      @      @       @      4@     `d@      &@      i@      "@              :@      2@     �b@     @d@      $@     �R@      @              �?       @      �?      @              $@                              �?      2@      @       @      "@      D@      @      @      @      3@     �c@      &@     �g@      "@              :@      1@     �`@     `c@       @     @P@      D@      &@      @      @      *@     �c@      @     `u@      @              @      $@      m@     �`@             �D@      (@      @              �?      @     �C@       @     �V@                      @              X@      A@              2@      (@      @              �?      @      C@       @     �U@                      @             @U@      A@              1@                                              �?              @                                      &@                      �?      <@      @      @      @      $@      ^@      @     `o@      @               @      $@      a@      Y@              7@      &@      @       @              "@      K@      @     �R@      �?              �?      @     �D@     �K@              (@      1@      �?      @      @      �?     �P@      �?      f@       @              �?      @      X@     �F@              &@      6@      @      @      �?      $@     @S@      �?     �d@      @              *@       @     @W@      :@       @      1@      @      �?                       @      0@              3@                      @              7@      @              @      @                                      @              $@                      @              (@       @                       @                                       @              @                      �?              (@                              �?                                      @              @                      @                       @                      �?      �?                       @      &@              "@                                      &@      @              @      �?                                      @               @                                       @                                      �?                       @      @              @                                      "@      @              @      2@      @      @      �?       @     �N@      �?     @b@      @              "@       @     �Q@      4@       @      ,@      2@      @      @      �?       @     �M@      �?      ]@      @               @       @      O@      3@       @      *@      (@      @      @      �?      @      >@      �?     @T@      @               @      �?      A@      .@      �?      (@      @              �?              �?      =@             �A@      @                      �?      <@      @      �?      �?                                               @              >@                      �?               @      �?              �?                                              �?              1@                      �?              �?      �?              �?                                              �?              *@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�܌.hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?t�i�?�	           ��@       	                     @����"�?H           Л@                           @0�xu~�?           ��@                          �1@��GD~�?�           ؑ@������������������������       �HTvϳ��?�            �m@������������������������       �K��G�:�?A           P�@                          �7@��aG��??            @]@������������������������       ���N����?'            �P@������������������������       ��A�f��?             I@
                           @�O&��?3           H�@                           �?@��@q��?�            pp@������������������������       �=�#>��?l            �h@������������������������       �[�6z���?)            @P@                          �6@����s�?�             p@������������������������       ��A�a�?b             d@������������������������       ��o5T)Q�?<            @X@                            @�;Q4�	�?:           ��@                            �?�XHQ��?�           �@                           @�����?�           ��@������������������������       ��U��<�?J           p�@������������������������       �j���� �?�             q@                           @te�Ӂ�?�            �s@������������������������       ��U�x�?�            @p@������������������������       ��Õty��?"             M@                           @ࠔ6J�?{           Ȃ@                          �3@`�ޚ@�?�            �u@������������������������       �{n`��?]            �a@������������������������       ������V�?�             j@                          @@@���?�            `o@������������������������       ��Q�O�
�?�            �m@������������������������       ���8��8�?             (@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `k@      A@     �E@     �@@     �]@     (�@      A@     Đ@      0@      @     �N@      M@     ��@     `�@      3@     �m@     @Z@      1@      =@      *@      S@     @t@      5@     �{@       @      @      A@      A@     �r@     �l@      "@      a@     �S@      $@      7@      &@      N@     `k@      2@     �q@      @      @      ;@      ;@     @i@      f@      @     �[@     �S@      $@      5@      &@     �K@     @i@      0@     @p@      @      @      ;@      ;@     @f@     �c@      @      U@      0@      �?      "@      �?      *@      7@      @     �D@      �?       @       @      $@      J@     �@@       @      4@      O@      "@      (@      $@      E@     `f@      (@     `k@      @      �?      3@      1@     �_@     @_@      @      P@      �?               @              @      1@       @      5@      �?                              8@      2@              :@      �?               @              @      &@       @      "@      �?                              .@      ,@              @                                              @              (@                                      "@      @              3@      :@      @      @       @      0@     @Z@      @      d@      �?      �?      @      @     �X@      J@      @      :@      0@              @       @      @      D@      @     �R@                      @       @      Q@      8@              .@      (@              �?               @      A@      @     �J@                      @       @     �J@      3@              ,@      @              @       @      @      @              6@                       @              .@      @              �?      $@      @                      &@     @P@             @U@      �?      �?              @      ?@      <@      @      &@      @      @                      "@      >@             �P@              �?              @      4@      *@              "@      @      @                       @     �A@              2@      �?                              &@      .@      @       @     �\@      1@      ,@      4@     �E@     v@      *@     ��@       @      @      ;@      8@     �|@     �r@      $@     �Y@      X@      *@       @      .@     �A@     p@      (@     �y@      @      �?      9@      5@     �r@     �m@      "@     �U@     �Q@      $@      @      ,@      :@     �j@      $@     pv@      @              0@      &@      m@     `f@      @     �L@     @P@       @       @      &@      3@     �f@      @     `o@      @              &@       @     �g@     �b@      @     �B@      @       @      �?      @      @     �A@      @      [@      @              @      @      E@      ?@       @      4@      9@      @      @      �?      "@      E@       @      I@      �?      �?      "@      $@     �Q@     �L@      @      =@      3@      @      @      �?      @      B@       @     �B@      �?      �?      @      $@      J@      L@      @      6@      @                              @      @              *@                      @              2@      �?              @      2@      @      @      @       @      X@      �?     �k@      �?       @       @      @     @c@      N@      �?      1@      @      �?      @      @      @     �C@             �a@               @       @      �?     �Z@      :@              &@      @                       @       @      &@             �C@                                      O@      1@              @      @      �?      @      @      @      <@             @Y@               @       @      �?     �F@      "@              @      &@      @      @               @     �L@      �?     �T@      �?                       @     �G@      A@      �?      @      &@      @      @               @      K@      �?     @T@      �?                       @      D@      A@      �?      @                                              @               @                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ$n8yhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @j}��lo�?�	           ��@       	                    �?��y:��?�           إ@                           @��_lw�?�           D�@                           @o�9�s��?M           `�@������������������������       ��7.�'�?;           �@������������������������       ��B����?           {@                            �?+>aj�?�            Pr@������������������������       ��A�e�?7            @W@������������������������       �0L�
F%�?{             i@
                            �?�Q��`�?�           l�@                          �0@�1x�y��?�           ��@������������������������       ��]�l�?%             Q@������������������������       ��!��&��?�           ��@                           @�=�����?�            @w@������������������������       �     �?T             `@������������������������       ��e���n�?�            �n@                           �?��R����?�           t�@                          �2@�ď�'@�?�            �s@                           @؁sF���?=             Y@������������������������       �<Cb�ΐ�?(            �P@������������������������       �JєX�?             A@                           �?6��컉�?�             k@������������������������       �     ��?Q             `@������������������������       ��
Z�b��?8            @V@                           @�I+��?            �@                           @��ϜR�?|           0�@������������������������       �#(����?Z            �a@������������������������       ���p֓�?"           �{@                           �?z5���?�            @k@������������������������       �p=
ףp�?             $@������������������������       �T!�����?�             j@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        l@      @@      A@      ;@     @W@     0�@     �@@     �@      3@      (@     �V@     �R@      �@     ~@      0@     �m@      f@      7@      4@      9@     @R@      }@      <@     x�@      ,@       @      T@     �P@     �~@     �v@      (@     �h@     �U@      "@      ,@      1@     �F@     �j@      (@     �q@      "@      @     �A@     �A@     `i@     �c@       @      X@     �P@      @      &@      1@     �D@     �d@       @     �j@      @      @      ?@      >@     �c@      Z@      @     �S@      :@      @      @      &@      7@     @U@      �?     �`@      �?              6@      @     �V@      J@      @     �E@      D@       @      @      @      2@     �S@      �?     �T@      @      @      "@      8@      Q@      J@       @      B@      4@      @      @              @      I@      $@     �Q@      @      @      @      @      F@     �J@       @      1@      @      �?                      @      &@      @      =@                       @       @      &@      2@      �?       @      1@      @      @                     �C@      @      E@      @      @       @      @     �@@     �A@      �?      "@     �V@      ,@      @       @      <@     �o@      0@     }@      @      �?     �F@      ?@     @r@     `i@      @     �Y@     �P@      *@       @      @      .@     @i@      0@     x@      @              9@      2@      m@     �a@      @     �P@      @                                      $@              ,@                      �?       @      1@      $@              $@      O@      *@       @      @      .@      h@      0@     0w@      @              8@      0@     �j@     @`@      @      L@      9@      �?      @      @      *@      I@              T@      �?      �?      4@      *@      N@     �O@      �?      B@      @              �?      �?      �?      (@              8@      �?      �?      "@      @      @@      1@              3@      3@      �?      @      @      (@      C@              L@                      &@      "@      <@      G@      �?      1@      H@      "@      ,@       @      4@     �f@      @     `y@      @      @      &@      "@      n@     @^@      @      C@      "@              @              @      J@      @     �X@                      @      �?     �T@     �B@              6@      �?              @                      $@              ;@                                     �E@      $@              @      �?              @                       @              5@                                      4@      "@              @                                               @              @                                      7@      �?               @       @                              @      E@      @     �Q@                      @      �?      D@      ;@              0@      @                              �?      =@      @      >@                      @      �?      4@      3@              ,@      �?                               @      *@             �D@                       @              4@       @               @     �C@      "@      &@       @      1@      `@       @     @s@      @      @      @       @     �c@      U@      @      0@      C@      @      "@      �?      &@     �X@      �?      j@      @      @      @       @     �Z@     �P@      @      ,@       @              @      �?      @      &@             �N@       @              @       @     �@@      $@               @      >@      @      @               @     �U@      �?     `b@      �?      @              @     �R@      L@      @      (@      �?       @       @      �?      @      >@      �?      Y@       @               @             �I@      2@               @                                               @              @                                      �?                              �?       @       @      �?      @      <@      �?     @W@       @               @              I@      2@               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�"bHhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �<@�BU]�?�	           ��@       	                    �?��"\u�?�           �@                            @�Z~"�?�           �@                           �?�ӟѰs�?�           ��@������������������������       �@�0�!��?Z             a@������������������������       �x/�ް~�?s           ��@                           �?e3�����?           �|@������������������������       �د!\�a�?3            �U@������������������������       �$����?�             w@
                          �0@��:�p��?�           ̞@                            @���D�?A            �Y@������������������������       �g(��Ү�?2            �S@������������������������       ��q�q�?             8@                           @I�'��?�           0�@������������������������       �Z�a�M�?           �@������������������������       ������}�?u           X�@                           �?�ҽe��?�             u@                           �?M��Cʨ�?U            �`@                            �?z͆����?"            �M@������������������������       ����:��?            �A@������������������������       �9��8���?             8@                            @k{L��N�?3            �R@������������������������       �2���h��?             C@������������������������       �������?             B@                           �?2(
�j�?|            `i@                            �?�ZI��?            �A@������������������������       �     ��?	             0@������������������������       ����Դ�?             3@                           @Sy'��?f             e@������������������������       �>v�禺�?M            �`@������������������������       �9��8���?             B@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @g@     �@@     �C@      :@     @Y@     ��@      =@     �@      9@      "@      N@      L@     ��@     @~@      .@     �q@     �d@     �@@      C@      :@     �V@     ��@      ;@     ؏@      6@      @     �J@      L@     ؅@     }@      ,@     �p@      U@      1@      9@      $@      J@     @q@      6@     �x@      1@      @      9@      8@     �q@     �l@      @      a@     �P@      &@      3@      $@      F@     �g@      1@     `o@      0@       @      1@      6@     �h@     �e@      @     @Z@      @      @      �?              @      .@             �C@      @              @              <@      ,@              1@      O@       @      2@      $@     �C@     �e@      1@     �j@      $@       @      ,@      6@     @e@     �c@      @      V@      1@      @      @               @     �U@      @     �a@      �?       @       @       @      U@      M@              @@       @               @              @      8@              2@                       @       @      ,@       @              (@      .@      @      @              @      O@      @      _@      �?       @      @             �Q@      I@              4@     �T@      0@      *@      0@      C@      t@      @     ��@      @       @      <@      @@     z@     @m@      @      `@      @                      @              9@              :@                              @      &@      *@              0@      @                      @              5@              &@                              @      "@      (@              ,@                                              @              .@                                       @      �?               @     @S@      0@      *@      *@      C@     pr@      @     ��@      @       @      <@      =@     `y@     �k@      @     @\@     �D@      "@      &@      $@      =@     `i@      @     pz@      @       @      (@      *@      s@     �b@       @     �O@      B@      @       @      @      "@      W@       @      f@      �?              0@      0@      Y@     �Q@      @      I@      3@              �?              &@      Q@       @     �_@      @      @      @              M@      3@      �?      2@      1@              �?              @      3@             �G@      �?               @              5@      $@      �?      @      @                              �?      (@              8@      �?              �?              (@       @              @      @                              �?      &@              &@                      �?              @      �?              @                                              �?              *@      �?                               @      �?                      ,@              �?              @      @              7@                      �?              "@       @      �?      @      �?              �?              @      @              &@                      �?              @      @              @      *@                              �?      @              (@                                      @       @      �?      �?       @                              @     �H@       @     �S@       @      @      @             �B@      "@              &@                                       @       @               @                                      @       @              @                                              @              @                                      �?      @              @                                       @      @              @                                      @      @              �?       @                               @     �D@       @     �Q@       @      @      @             �@@      �?              @       @                               @      :@       @      O@       @      @      @              5@      �?              @                                              .@              "@                                      (@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJq��(hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             @�Hr|�x�?�	           ��@       	                    �?�^��x�?W           "�@                          �<@����a8�?^           t�@                            �?)�Tc>�?'           �@������������������������       �F`��C)�?�            �s@������������������������       �ͻ�mz�?g           0�@                            �?��˜�G�?7            �V@������������������������       �`!�2���?            �G@������������������������       �D��2(�?             F@
                           �?�|}F��?�           И@                            @6?,R��?f            �@������������������������       �C�W�0t�?           �{@������������������������       �j@����?U            ``@                           �?6����j�?�           ��@������������������������       �NQf���?W            �a@������������������������       ���9����?<           8�@                          �;@wyqW�?c           ��@                          �0@�ܺ���?           8�@                           @���H�~�?              G@������������������������       ��P�a�r�?             >@������������������������       �     @�?
             0@                            @��4t4��?�           Ȉ@������������������������       �������?�           ��@������������������������       ������?z            `g@                          �@@��Wk�?G            @\@                           �?������?@            �Y@������������������������       �}��7�?             6@������������������������       �:�ci�~�?4            @T@������������������������       �H�z�G�?             $@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      7@     �C@      ;@     @^@     Ѓ@      ?@     ��@      ,@      "@     �T@     �P@     p�@     p@      2@     �o@     `d@      3@      @@      8@     �Z@     �{@      3@     H�@      @      @      Q@      J@     X�@     0v@      .@     �g@     @T@      ,@      5@      .@     �Q@     @j@       @     �t@      @       @      A@      @@      q@      e@      @     �Y@     �R@      &@      3@      .@      O@     @i@       @     pr@      @       @      =@      ?@      p@     �d@      @     �Y@      7@      �?      �?       @      "@     �H@       @     �W@      �?              @      $@      Q@     �C@       @       @     �I@      $@      2@      *@     �J@      c@      @      i@      @       @      6@      5@     �g@     �_@      �?     �W@      @      @       @              "@       @              B@                      @      �?      ,@      @       @      �?      @      @       @              @      @              *@                      @              "@      �?                      @                              @       @              7@                              �?      @       @       @      �?     �T@      @      &@      "@      B@     `m@      &@     ��@       @      @      A@      4@     �s@     @g@      $@     �U@      E@      �?      @      @      .@     @V@      �?     �e@                      @      "@      `@     @R@      �?      <@      E@      �?      @       @      ,@     �R@      �?     @]@                      @       @     @X@     �K@      �?      6@                               @      �?      ,@             �L@                              �?      @@      2@              @      D@      @       @      @      5@     @b@      $@      w@       @      @      ;@      &@     @g@     @\@      "@      M@      @              @      @      @      6@             �Q@              @      @              3@      @              @      B@      @      @       @      1@      _@      $@     �r@       @      �?      7@      &@     �d@      [@      "@     �K@     �D@      @      @      @      ,@     �g@      (@     pp@      @      @      .@      ,@     `d@     �b@      @     �P@      C@      @      @      @      ,@     �d@      (@     `j@      @      @      .@      ,@     �a@     �`@      @     @P@      @              �?               @      "@              @                               @      @      ,@       @       @      @              �?                      @              @                               @      @      @       @       @      �?                               @       @                                                       @      "@                     �@@      @      @      @      (@     �c@      (@      j@      @      @      .@      (@      a@     �]@      �?     �O@      ;@      @      @      @      (@     �^@      (@      b@      @      @      ,@       @      X@     �V@              M@      @      �?       @                     �A@             �O@                      �?      @     �D@      <@      �?      @      @                                      6@              J@                                      4@      .@              �?       @                                      6@             �H@                                      4@      "@              �?                                              @              @                                      �?      @                       @                                      .@              E@                                      3@       @              �?      �?                                                      @                                              @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJMBhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @ң���?�	           ��@       	                    �?�*���?�           �@                            �?SQ�4md�?           ̓@                          �=@��/z�1�?P           ��@������������������������       ���U��G�?6           x�@������������������������       ��������?             D@                           �?���?�            �s@������������������������       �J�_cV�?             ;@������������������������       �x������?�            r@
                           @���4V�?�           D�@                           �?X6��@b�?N           0�@������������������������       ��.�6���?�             w@������������������������       ���a�i��?d           ��@                           @"����!�?�           X�@������������������������       ��*'b�?�            Px@������������������������       �}-�ì��?�            �l@                           @X���?�?�           �@                          @@@b�Њ6*�?�           ��@                           �?��Y=�?�           �@������������������������       ���3�[d�?�            �s@������������������������       ��JV=�?�            �v@������������������������       �4և����?	             ,@                           �?=Ea<*�?           @y@                          �;@B�X5�p�?�            �m@������������������������       ��2�^�?�            �g@������������������������       ��i�q���?              I@                          �5@p�r��?n            �d@������������������������       ���Z=;�?<             V@������������������������       �3�m���?2            �S@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        j@      ;@      I@      5@     �_@     P�@      8@     x�@      *@      @     @T@     �L@     Ї@     ~@      8@     �p@     �d@      2@      B@      4@      X@     �~@      .@      �@      (@      @     @R@     �E@     �@     �v@      5@     @j@     �U@      $@      5@      &@      Q@     @n@      @     �q@      "@       @     �B@      8@     �j@      b@      "@      Y@     �Q@      @      *@      "@      L@     �h@      @     �k@      @      �?      =@      0@      d@     @X@      @      P@     @Q@      @      *@      "@     �I@      h@      @     �h@      @      �?      =@      0@     `c@     @W@      @      P@      �?                              @      @              6@                                      @      @                      0@      @       @       @      (@      G@      �?     @P@      @      �?       @       @      J@      H@      @      B@                      @               @      �?               @      @                              @      �?              @      0@      @      @       @      $@     �F@      �?     �L@      �?      �?       @       @     �H@     �G@      @     �@@     �S@       @      .@      "@      <@     `o@      $@     `|@      @       @      B@      3@     pr@     �k@      (@     �[@      K@      @      &@      @      2@     �c@      @     �p@      @       @      *@      *@      g@      [@       @     �R@      1@      @              �?      $@     �L@       @     �T@                      @      @      U@      J@      @     �D@     �B@       @      &@      @       @     @Y@      @     `g@      @       @      @      @     @Y@      L@      @     �@@      9@      @      @      @      $@     @W@      @      g@                      7@      @     �[@     �\@      @      B@      2@      �?      @       @      @      N@      �?     @[@                      *@      @     @P@     �U@      @      0@      @       @               @      @     �@@       @     �R@                      $@       @     �F@      ;@      �?      4@     �E@      "@      ,@      �?      ?@     �c@      "@     �w@      �?      �?       @      ,@     �o@     �\@      @     �K@      8@      @      $@      �?      6@      V@      @     �l@      �?              @      $@     �f@     @P@              D@      5@      @      $@      �?      2@     �U@      @     �l@      �?              @      $@     �f@     @P@             �B@      (@      @      @              0@      L@      @      T@                      @      �?     �R@      B@              3@      "@              @      �?       @      ?@             �b@      �?              @      "@      [@      =@              2@      @                              @      �?              @                                                              @      3@      @      @              "@     @Q@      @     `b@              �?      �?      @     @R@     �H@      @      .@      ,@       @      @              @     �A@      @     �X@              �?               @      A@      >@      @      @      &@       @      @              @      6@      @     @R@              �?               @      <@      >@      �?      @      @                                      *@              :@                                      @               @              @      @                      @      A@      �?      H@                      �?       @     �C@      3@              "@      @      �?                       @       @      �?      @@                      �?       @      5@      $@              @              @                       @      :@              0@                                      2@      "@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�cB0hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @��Ȣn�?�	           ��@                            �?k�n���?�           �@                           !@_�\�Vc�?$           D�@                           �?�<�F^�?           ,�@������������������������       ��#���)�?9           ��@������������������������       ��r�r���?�           \�@������������������������       ��8��8��?             (@                           @VIϩE��?�           ��@	       
                   �2@*
��V��?J           �@������������������������       ��W�o���?j            �e@������������������������       �Q�`�S��?�             w@                          �:@�+^ �?q            �f@������������������������       ��"e����?^             b@������������������������       ����e�?            �C@                           �?5����?�           L�@                           @S�0qX�?0           �}@                          �0@�c���?�            @x@������������������������       �      �?             0@������������������������       �80V���?�            @w@                          �4@�Eq�Ȟ�?=            �V@������������������������       ��x?r���?            �@@������������������������       ��d�����?'            �L@                           @�Yd��?�           ��@                           @�Z&rA��?/            }@������������������������       �t<iE���?�            �x@������������������������       ��Kh/���?2             R@                           @Y��I�?f            �d@������������������������       �a'q���?[            �b@������������������������       �     ��?             0@�t�b��     h�h4h7K ��h9��R�(KKKK��h��B�       @i@      9@      D@      =@     �[@     `�@      9@     ��@      2@      *@     @T@      N@     ��@     (�@      "@     �n@     �c@      1@      <@      7@      U@     �}@      7@     ؆@      *@      &@     �Q@     �I@     �@      y@      "@     `i@      [@      (@      *@      4@     �L@     �v@      2@     ��@      $@       @     �F@      ;@     �x@     0q@      @      `@      [@      (@      *@      4@     �L@     �v@      ,@     ��@      $@       @     �F@      ;@     �x@     0q@      @      `@      K@      @      *@      *@     �H@      e@      @     �j@      @       @      :@      $@     �c@      [@      �?     @P@      K@      @              @       @      h@      $@     �w@      @              3@      1@      n@     �d@      @      P@                                              @      @                                               @                             �H@      @      .@      @      ;@     �[@      @     �`@      @      "@      9@      8@     �[@     @_@      @     �R@     �D@       @      $@      @      5@     �V@      @     @U@       @      @      3@      5@     @U@     @V@      �?      N@      .@              @      �?      @     �A@       @      ;@                      $@      &@      "@      ;@              :@      :@       @      @       @      .@      L@       @      M@       @      @      "@      $@      S@      O@      �?      A@       @      @      @              @      3@      �?      I@      �?       @      @      @      9@      B@      @      ,@      @      @      @              @      1@      �?      ;@      �?              @      @      4@      >@      @      ,@      �?                                       @              7@               @                      @      @                     �F@       @      (@      @      ;@     �e@       @     �x@      @       @      &@      "@      o@     @]@              F@      3@      @      $@      �?      3@     @U@      �?     @a@      @      �?      $@      @     �W@      N@              :@      1@      @      "@      �?      1@      Q@             �Y@      @              "@       @     @T@     �I@              6@                                                              @                      �?       @      @      @              �?      1@      @      "@      �?      1@      Q@             �X@      @               @              S@     �G@              5@       @      �?      �?               @      1@      �?      B@              �?      �?       @      *@      "@              @              �?                       @       @      �?      2@                      �?       @       @       @               @       @              �?                      .@              2@              �?                      &@      @               @      :@       @       @      @       @     �V@      �?      p@      �?      �?      �?      @     @c@     �L@              2@      0@               @      @      @     �K@      �?     �i@      �?      �?              @     �]@     �C@              &@      (@               @      @      @     �F@      �?     �f@      �?      �?              �?     @W@      ?@              &@      @                                      $@              7@                               @      9@       @                      $@       @                       @     �A@              J@                      �?       @      B@      2@              @      $@       @                       @      ;@             �I@                      �?       @      A@      .@              @                                               @              �?                                       @      @               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�VXhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @>��Q���?�	           ��@       	                   �4@�!�u��?N           ��@                           @�LW$���?           ��@                           @&���W�?�           8�@������������������������       �xP�#NM�?D           �@������������������������       �l~X�<�?<             [@                            �?P��z	�?�            `m@������������������������       ��Z:$l�?J            �]@������������������������       ��Rpo�?J             ]@
                           �?�/����?:           ��@                          �;@����?�            @y@������������������������       ��E�_��?�             u@������������������������       �ʜoB��?,             Q@                          �>@c��-���?E           �@������������������������       ��/&���?*           �|@������������������������       �},܋;��?            �I@                           �?/�4�~�?e           Π@                          �<@0��F���?U           ��@                           @<��4��?-           �@������������������������       ���\\��?�           �@������������������������       �     ��?R             `@                           @�Z�LY��?(            �N@������������������������       �R?��yq�?            �A@������������������������       ��q-�?             :@                          �;@�t|�9�?           ��@                          �9@�� 
���?�           �@������������������������       ��T�n�?o           ��@������������������������       ���߭Q�?6            �T@                           @X^g�}��?k            �d@������������������������       ��iQT�?3            �U@������������������������       �1�N!T�?8            �S@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      9@      <@      8@     �Z@      �@     �A@     ܐ@      2@      @     �V@     �O@     x�@     h�@      4@     0r@     @[@      *@      2@      *@      J@      r@      (@      }@      "@       @     �B@      ?@     �v@     �i@      @     �`@     �O@      @      @       @      >@     ``@      @     �h@      �?              1@      1@     �h@      \@      �?     �O@     �D@      @      @      @      2@     @X@      @      `@                      @      @     �e@      T@             �E@      ;@      �?      @      @      ,@      V@      @     �\@                      @      @     �`@     �Q@              B@      ,@       @              @      @      "@              *@                      �?       @     �E@      "@              @      6@              �?      �?      (@      A@              Q@      �?              $@      $@      7@      @@      �?      4@      0@                              @      0@             �D@      �?              �?      @      ,@      *@      �?      @      @              �?      �?      @      2@              ;@                      "@      @      "@      3@              0@      G@      $@      ,@      @      6@     �c@      @     �p@       @       @      4@      ,@      e@     �W@      @      R@      6@      @      (@       @      &@     @Q@       @      Z@      @      �?      (@      @     @Q@      H@      @     �B@      0@               @       @      "@      O@       @     �T@       @      �?      @      @      O@      E@      @      A@      @      @      @               @      @              6@      �?              @              @      @              @      8@      @       @      @      &@      V@      @     �d@      @      �?       @      $@      Y@     �G@             �A@      7@      @       @      @      "@      S@       @     �c@                       @      @      V@      G@              ?@      �?                               @      (@       @       @      @      �?              @      (@      �?              @     �X@      (@      $@      &@      K@     @x@      7@     8�@      "@      @      K@      @@      v@     �s@      .@     �c@     �H@      @       @      �?      ;@     �e@      *@     @l@      @      �?      2@      (@     �c@      _@      @     �P@      E@      @       @      �?      8@     @e@      *@     �h@      @      �?      1@      (@      c@      ]@      @     �P@     �A@      @       @      �?      1@     �`@      "@     `d@      @              0@      (@     `a@     @Y@      @     �L@      @                              @     �A@      @      B@              �?      �?              *@      .@              "@      @                              @      @              ;@                      �?              @       @       @      �?      @                              @      @              *@                      �?              �?      @       @      �?       @                                                      ,@                                      @      @                     �H@      @       @      $@      ;@     �j@      $@     Px@      @      @      B@      4@      h@     @h@       @     @V@     �H@      @       @      $@      ;@     `f@      $@     ps@       @      @      @@      3@     @e@     �f@      @     @T@     �G@      @       @      @      6@      e@      $@     �r@       @       @      =@      2@     @b@     `d@      @     @S@       @                      @      @      &@              $@              �?      @      �?      8@      3@              @                                              A@             �S@      @              @      �?      7@      (@      �?       @                                              4@              B@      @                              .@      @      �?       @                                              ,@              E@      �?              @      �?       @      "@                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�5hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?��D E��?�	           ��@       	                   �:@�6n�5�?e           �@                           �?�6u�Q�?�           ��@                           @��6�R�?�            @l@������������������������       �T��Ǐ�?~            `j@������������������������       �ƒ_,���?             .@                            �?x�FXB�?S           4�@������������������������       ������?�           8�@������������������������       �f恰B�?�           0�@
                            @x=i��?�            �j@                          �=@UUUUUU�?`             b@������������������������       �I�����?D            �Z@������������������������       �,���y4�?             C@                          �=@s��\;0�?,            @Q@������������������������       ��˔�&E�?            �F@������������������������       ��q�q�?             8@                            @�V%��?H           ��@                            �? #51��?�           ܗ@                            �?���$�?�           �@������������������������       �&���^��?l            �@������������������������       ��lb��?g           ��@                           @��}ڥ��?�            �w@������������������������       ���	,��?�            q@������������������������       �p�U��?E            �Z@                           @�ad�	�?�           p�@                           @f�:G�)�?f           �@������������������������       �I���2�??           �~@������������������������       ��lV}��?'             I@                           5@��s���?            �H@������������������������       ���uJ���?             3@������������������������       �4�ͫ��?             >@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        j@      E@      B@      <@     @_@     �@      B@     ̐@      7@      @     @W@     �G@     ��@      �@      5@     @p@     �\@      6@      :@      $@     �Q@     �t@      2@     {@      0@      @      G@      9@      r@     �m@      @      b@     �X@      1@      9@      $@     �P@     Ps@      1@      v@      .@      @     �C@      8@     �o@      k@      @      `@      $@      @       @      �?      *@      ?@       @      O@      &@              &@       @      A@      :@              1@      $@      @       @      �?      &@      ?@       @      K@      &@              &@       @      =@      :@              1@                                       @                       @                                      @                             @V@      *@      7@      "@     �J@     `q@      .@     @r@      @      @      <@      6@     �k@     �g@      @     �[@     �G@      @      &@      @     �@@      f@       @      c@      @              (@      ,@      \@     �V@      @     �Q@      E@      $@      (@      @      4@     @Y@      @     `a@      �?      @      0@       @      [@     @Y@       @     �D@      0@      @      �?              @      8@      �?     �S@      �?              @      �?      B@      5@              0@      $@      @      �?              @      0@      �?      H@      �?              @              5@      1@              ,@      @      @      �?               @      *@      �?      =@      �?              @              4@      (@              *@      @                              @      @              3@                                      �?      @              �?      @       @                               @              ?@                              �?      .@      @               @       @       @                              @              8@                                      @      @              �?      @                                       @              @                              �?       @      �?              �?     �W@      4@      $@      2@      K@      u@      2@     �@      @       @     �G@      6@     `{@     `q@      .@      ]@     �R@      .@      "@      ,@     �D@     @p@      1@      y@      @       @      F@      4@      s@      j@      &@      X@     �G@      (@      @      &@      9@     �j@      ,@     pt@      @              5@      *@     �n@     �a@       @      P@      2@      @      @      "@       @     @Y@      &@     �f@      @              @      @     �_@     @T@      �?      5@      =@      @      �?       @      1@     �\@      @     `b@       @              2@      $@     �]@      O@      �?     �E@      ;@      @      @      @      0@     �F@      @     �R@      �?       @      7@      @      O@     �P@      "@      @@      5@      @       @      @      (@      >@       @     @P@                      .@      @      H@      C@      @      9@      @              @              @      .@      �?      $@      �?       @       @      �?      ,@      <@      @      @      4@      @      �?      @      *@      S@      �?      n@                      @       @     �`@     @Q@      @      4@      4@       @      �?      @      *@     �Q@      �?     �j@                      @       @     @_@      O@      @      2@      3@      �?      �?      @      *@      M@      �?      h@                      @       @     �]@      L@      @      1@      �?      �?                              *@              6@                                      @      @              �?              @                              @              9@                                      @      @               @              @                                              *@                                      @                                                                      @              (@                                      @      @               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJeIhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@�vb5`�?�	           ��@       	                    �?��p.���?z           �@                           @O�W���?Y           ��@                          �3@	�����?�            �u@������������������������       �Gsd���?^            @_@������������������������       � ߦ�5�?�            `k@                            �?v��~{�?w            �h@������������������������       ����?J            �^@������������������������       �x������?-            �R@
                            @��v��?!           ܦ@                           @���p}��?,           �@������������������������       ���vy8��?�           ��@������������������������       �A�Q�,�?c           ��@                          �2@�D�̐��?�           �@������������������������       ��~��B�?�             m@������������������������       �JSMI��?`           ��@                           �?�۴d�?           �{@                           �?�@G���?�            `o@                           @'����??            @X@������������������������       �2B�f�?0            �R@������������������������       ��\@˜��?             7@                           �?p1/CD�?]            @c@������������������������       �*wj��?             G@������������������������       ��3�\���?B             [@                          �@@Yy�o���?y            @h@                           �?�A����?s            `g@������������������������       ��W4�	�?3            �S@������������������������       �j�pW�$�?@             [@������������������������       ��$I�$I�?             @�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@      ;@      8@      9@      \@     ؅@      1@     4�@      *@      @     �T@     �I@     ��@     �}@      .@     �q@      e@      :@      6@      9@     �Y@     �@      1@     p�@      $@      @     �R@      G@      �@     p{@      (@     Pp@      4@      �?      @      @      5@      O@      �?     �e@      @              ,@      @      [@      P@      �?      K@      *@              @      @      0@      E@             �W@       @              $@      @     �Q@      A@              H@      @                              @       @              G@                      �?       @      >@      0@              (@      @              @      @      (@      A@             �H@       @              "@      @     �D@      2@              B@      @      �?       @       @      @      4@      �?      T@       @              @             �B@      >@      �?      @      @      �?               @      @      (@      �?      J@                      @              ?@      $@               @       @               @               @       @              <@       @                              @      4@      �?      @     �b@      9@      .@      4@     �T@     (�@      0@     ��@      @      @      N@     �D@     ��@     pw@      &@     �i@     �_@      4@      ,@      0@      S@     �y@      &@      �@      @      @      I@      >@      y@     Pr@      &@     �e@     �Q@      "@      "@      0@      9@     �m@      @     @p@      �?       @      0@      @     `n@      e@      @     �T@      L@      &@      @             �I@     `f@      @      p@       @      @      A@      9@     �c@     @_@       @      W@      7@      @      �?      @      @     �`@      @     `o@      @      �?      $@      &@     �h@     �T@             �@@      (@                      @       @      >@      �?     @Q@                      �?       @     @U@      3@              "@      &@      @      �?      �?      @      Z@      @     �f@      @      �?      "@      "@     �[@     �O@              8@      7@      �?       @              "@      V@             �c@      @               @      @     @U@     �B@      @      6@      .@      �?       @              @     �M@              U@                      @      @      A@      0@      @      4@      "@               @              @      (@              ?@                      @      �?      &@      @      �?      *@      @               @              @      (@              5@                      @      �?      "@      @      �?       @       @                                                      $@                                       @      @              @      @      �?                      �?     �G@             �J@                       @      @      7@      "@       @      @      @                                      0@              &@                              �?      @      @              @      @      �?                      �?      ?@              E@                       @       @      0@      @       @      @       @                               @      =@             �R@      @               @      �?     �I@      5@               @      @                               @      =@             @R@      @               @      �?     �I@      1@               @      @                              �?      &@              =@                                      5@      $@                                                      �?      2@              F@      @               @      �?      >@      @               @      �?                                                       @                                              @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJN�ckhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @��\��?�	           ��@       	                   �;@�Ú,,�?�           �@                            �?G3V��=�?           ��@                          �:@�I=��?�           P�@������������������������       �M�%e��?u           l�@������������������������       ���-���?"            �L@                           @:|E�L�?�           ��@������������������������       �<7_#/T�?&           �}@������������������������       �òrr}�?]            �d@
                           �?g{Iͤ�?�             r@                           @K�%���?L            �^@������������������������       ��Q#1�?             �G@������������������������       �.窷�?,             S@                           @�6~�7�?m            �d@������������������������       �c��7w�?[            �`@������������������������       �ʤ��IF�?            �@@                           @eh��k��?�           T�@                          �0@&���^��?�           ��@������������������������       ������?             7@                           �?��\m���?�           ȅ@������������������������       �	��fUH�?�             u@������������������������       �tv��M �?�            pv@                           �?��&Q��?�            Px@                           �?     ��?)             P@������������������������       �36�v[�?             7@������������������������       ��E��{�?            �D@                           @������?�            Pt@������������������������       �nt{����?�            �o@������������������������       �%ޑ���?*            �Q@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      B@     �C@      ;@      [@     �@      ?@     ��@      0@      @     �S@     �Q@     x�@      �@     �A@     �o@     `d@      9@      ;@      7@      U@     �|@      :@     ��@      *@      @     �P@      N@     �@     px@      @@     �k@      c@      5@      8@      7@     @T@     Py@      9@     ��@      (@      @      N@     �K@     �|@     �v@      @@     @i@     @\@      (@      .@      0@     �E@     pt@      3@     P~@       @      �?      A@     �@@     �v@     @p@      3@     �`@     @\@      (@      .@      0@      E@     0t@      1@     @}@       @      �?      A@     �@@     pu@     �o@      3@      `@                                      �?      @       @      1@                                      5@      @              @      D@      "@      "@      @      C@     �S@      @      [@      $@      @      :@      6@      X@     �Y@      *@     @Q@      C@      @      @      @     �A@      Q@      @      S@      @      @      0@      4@      R@     �P@       @     �G@       @       @      @              @      $@      �?      @@      @              $@       @      8@     �B@      &@      6@      $@      @      @              @     �J@      �?     �[@      �?              @      @      G@      <@              3@      @       @      @              �?      0@              F@                      @              1@      1@              *@      @              @                      "@              4@                       @              @       @              @      @       @                      �?      @              8@                      �?              *@      .@              $@      @       @                       @     �B@      �?     �P@      �?              @      @      =@      &@              @      @       @                       @      9@      �?     �K@      �?              @      @      3@      &@              @                                              (@              &@                                      $@                             �E@      &@      (@      @      8@      g@      @     �z@      @      �?      &@      $@     �j@     @_@      @      ?@      @@      @       @      @      2@     @\@       @     pp@       @              "@      @     �d@     �S@              3@                                              �?              1@                              �?      @      �?                      @@      @       @      @      2@      \@       @     �n@       @              "@       @     @d@     �S@              3@      5@       @      @      @      0@     �Q@       @     �W@      �?              @             �N@     �D@              (@      &@      �?      �?      �?       @     �D@             �b@      �?              @       @     @Y@     �B@              @      &@       @      @              @      R@      @     �d@      �?      �?       @      @      H@      G@      @      (@      @               @              @      @              :@                                      @      (@               @      @                               @      �?              $@                                       @      @               @       @               @              @      @              0@                                      @      "@                      @       @       @              �?     �P@      @     `a@      �?      �?       @      @      E@      A@      @      $@      @       @       @              �?      I@      @     �\@      �?      �?      �?      @      :@      6@      @      "@                                              0@              8@                      �?              0@      (@              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��2hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @$N�R�?�	           ��@       	                    �?cc>�y��?�           ԥ@                          �=@�&�I�l�?	            �@                           @\�N04��?�           D�@������������������������       ���G[Iy�?�           �@������������������������       �F]t�E�?             &@                           �?�-%*��?            �K@������������������������       ���_[��?             ?@������������������������       �      �?             8@
                           @�Ub�'�?�           ��@                            �?�y��y��?�            �@������������������������       ��>'ʇ�?5            @������������������������       �*	a�.��?k            �e@                           @ѳڻ N�?-           �@������������������������       �n{�7��?�           (�@������������������������       ��9+���?b            �c@                          �;@$��=R��?�           |�@                           @���2�?o           0�@                          �0@�Q�ޒ��?�           p�@������������������������       �     ��?             @@������������������������       �*�փ��?�           p�@                           @R�n��?�             k@������������������������       �L�Zͺ(�?�            �h@������������������������       �>
ףp=�?             4@                           �?b�H�/��?Z             c@                           �?�>4և��?$             L@������������������������       �^����T�?            �C@������������������������       �$�ɜoB�?             1@                           @81�P��?6            @X@������������������������       ���E���?)             R@������������������������       ����H�?             9@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      ?@      G@      :@     @Z@     ��@      <@     H�@      2@      @     �T@     �L@     ȇ@     �~@      6@     @l@     @d@      6@      @@      8@     �T@     �{@      6@     ��@      *@      @     �R@     �H@     ��@     0w@      0@      g@     �U@      .@      6@      &@      H@      j@      (@     �q@      "@       @      A@      <@     �j@     �d@       @     @T@      U@      .@      6@      &@      G@     �i@      (@     �o@      "@       @      A@      <@     @j@      c@       @     @S@     �T@      .@      6@      &@      G@     @i@       @     �o@      "@       @      A@      <@     @j@     �b@       @     @S@       @                                       @      @                                                      @                      @                               @      @              :@                                      @      (@              @      @                              �?      @              1@                                              @              @                                      �?                      "@                                      @      "@              �?     �R@      @      $@      *@     �A@     �m@      $@     �}@      @      �?     �D@      5@     �s@     �i@       @     �Y@      E@      @      �?      @      (@     �X@      @     �i@      �?              .@      @      e@     @P@       @      E@      A@       @              @      "@      U@      @     @d@      �?              "@      @      \@      H@      �?      9@       @       @      �?      �?      @      .@             �E@                      @      @      L@      1@      �?      1@     �@@      @      "@      "@      7@     �a@      @      q@      @      �?      :@      ,@     �b@     �a@      @     �N@      >@       @      @      @      7@     �\@      @     �j@      @      �?      4@      (@     @]@     �_@      @     �L@      @      �?      @      @              :@      �?     �M@                      @       @     �@@      ,@              @      F@      "@      ,@       @      6@      h@      @     �y@      @      @      @       @     �l@     �]@      @      E@     �A@      "@      *@       @      1@     @d@      @     u@      @      �?      @       @     �j@      \@      @      C@      =@      @      $@       @      .@     @]@      @     @q@      �?              @      @     �e@     �S@              @@                                              �?              4@                                      @      @              �?      =@      @      $@       @      .@      ]@      @      p@      �?              @      @     �d@     �R@              ?@      @      @      @               @     �F@       @     �N@       @      �?      �?      @      D@      A@      @      @      @      @      @               @      B@       @      M@       @      �?      �?      @      B@      >@      @      @                                              "@              @                                      @      @                      "@              �?              @      >@             �R@       @       @                      1@      @       @      @       @              �?              @      @              7@      �?                               @      @       @       @       @                              @      @              ,@      �?                              @      @       @                              �?                      �?              "@                                      @      �?               @      �?                               @      :@             �I@      �?       @                      "@      @               @      �?                               @      &@              E@      �?       @                      "@       @               @                                              .@              "@                                              �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�I�YhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @���Y���?�	           ��@                            �?G�ɺd"�?�           ܥ@                           !@��2��?8            @                           @b�М��?0           ��@������������������������       ��s仠��?[           ��@������������������������       �X�@�C��?�           �@������������������������       ���X��?             ,@                          �;@ؐ���?�           h�@	       
                   �2@mSV_��?�           ��@������������������������       ���
цO�?�             j@������������������������       �w�*Qޤ�?            x@                           @'#rp���?(            �M@������������������������       �2�A���?             �H@������������������������       ����(\��?             $@                           �?�E�(�&�?�           l�@                           @z��7#�?�           ��@                           �?w.U��?�            �r@������������������������       �?�����?|            @h@������������������������       ����/��?A            �Y@                           �?�K�`�?�            0w@������������������������       ����(�#�?C            @X@������������������������       ��u�N��?�             q@                           @ϵ1�#��?           �{@                           �?�$V.�H�?�            �h@������������������������       �H���0��?H            �Z@������������������������       �\��m�?<            �V@                           �?
�Q���?�             o@������������������������       �5���_�?F             ]@������������������������       ��W�����?T            �`@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �l@      :@     �@@      ;@     �Z@     @�@     �C@     �@      :@      @     @W@      N@     ��@     p�@      2@     �p@      f@      5@      <@      7@      W@      ~@      >@     X�@      2@      @      S@      J@      @     Px@      1@     �j@     �_@      1@      7@      3@      P@     0x@      7@      �@      *@      �?      G@      >@     0x@     Pq@      $@      b@     �_@      1@      7@      3@     �O@     �w@      5@     ��@      *@      �?      G@      >@     x@     Pq@      $@      b@     @R@      @      4@      $@      ;@     �g@      "@     �p@      @              6@      (@     �e@      \@       @      K@      K@      &@      @      "@      B@     �g@      (@     0s@       @      �?      8@      2@     �j@     �d@       @     �V@                                      �?       @       @      �?                                       @                             �H@      @      @      @      <@     @W@      @     �Z@      @      @      >@      6@     @[@      \@      @     �P@     �F@      @      @      @      <@      U@      @      U@      @      @      <@      5@     �X@     �Z@      @     @P@      9@      �?      @      �?      $@      <@       @      5@               @      (@      (@      4@     �D@      @      9@      4@      @       @      @      2@      L@      @     �O@      @       @      0@      "@     �S@     �P@              D@      @                                      "@              7@                       @      �?      &@      @       @       @      @                                      "@              3@                       @      �?      @      @       @       @                                                              @                                      @      �?                     �J@      @      @      @      ,@      e@      "@     �x@       @       @      1@       @     �l@      a@      �?      K@      B@       @      @      @      @      W@      @      o@      @       @      $@      @     �\@      X@      �?     �A@      "@              @       @      @      <@             @\@      @      �?       @       @     �M@      C@              8@      @               @              @      7@             �Q@                      �?       @      E@      <@              4@      @               @       @       @      @             �E@      @      �?      @              1@      $@              @      ;@       @      �?      �?       @      P@      @      a@      @      �?       @      @      L@      M@      �?      &@       @                               @      ,@       @      B@                       @              $@      2@              @      3@       @      �?      �?              I@      �?      Y@      @      �?              @      G@      D@      �?      @      1@      @              �?      @      S@      @     �b@      �?              @      @      ]@     �D@              3@      *@                      �?      �?      6@       @     �P@                      @      �?     �O@      0@               @      @                      �?              0@       @      ?@                      @              9@      ,@               @      @                              �?      @              B@                              �?      C@       @                      @      @                      @      K@      @     �T@      �?              @       @     �J@      9@              &@                                      @      ;@      @      =@                               @      @@      @              $@      @      @                              ;@              K@      �?              @              5@      3@              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @B�)��?�	           ��@       	                     @��u8,��?�           ��@                           @@���-�?\           ��@                          �0@����?7           �@������������������������       �s��i;��?6            @S@������������������������       �9����?           ܒ@                            �?�Z"��?%           D�@������������������������       ����	���?           |@������������������������       �X�YEx�?           ��@
                           @G�6��?�           $�@                           �?1NW�u��?!           8�@������������������������       �rO�?�            x@������������������������       �r���.�?&           `|@                           @F�d�+��?z            @h@������������������������       ���N8�?             5@������������������������       ��ҵ�f��?l            �e@                          �<@�@'��?�            �v@                           @!� ��?�            �s@                            �?�� F(�?�            �q@������������������������       �B{	�%��?)             R@������������������������       ��E�nnE�?�             j@                            �?�"��r�?             ?@������������������������       �t�E]t�?	             &@������������������������       ��p=
ף�?             4@                           �?�������?            �I@                            �?H��	,�?             7@������������������������       �      �?              @������������������������       ��h$��W�?             .@                           @
^N��)�?             <@������������������������       �@4և���?             ,@������������������������       �d}h���?             ,@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `f@     �@@      C@     �B@     �Z@     ��@      >@     ��@      ,@      "@     �R@     �R@     ��@     X�@      6@     @p@     �d@     �@@     �B@      B@     @Y@     h�@      8@     �@      ,@      "@     �P@     @R@     ��@     P}@      6@     �l@     �^@      :@      =@      <@     @U@      |@      2@     p�@      &@       @      L@     �O@     p{@      v@      4@     �g@     �Q@      1@      4@      3@     �I@      n@      "@     �s@       @       @      5@     �@@     �l@     @b@      "@     �V@       @                              @      <@      �?       @                      �?      @      *@      "@              @      Q@      1@      4@      3@     �F@     �j@       @     `s@       @       @      4@      <@      k@      a@      "@     �U@      J@      "@      "@      "@      A@     �i@      "@      s@      @      @     �A@      >@     @j@     �i@      &@     �X@      *@      @       @      �?       @      T@       @     �`@      �?               @      @     �U@     �R@      @      8@     �C@      @      @       @      :@     �_@      @     `e@       @      @      ;@      7@     �^@     ``@      @     �R@      F@      @       @       @      0@     �e@      @     �v@      @      �?      &@      $@     `k@     @]@       @     �D@     �@@      @      @       @      (@      _@      @      s@      �?               @      @     `h@     @X@      �?     �@@      6@      @      @       @       @      R@      @     �[@                      @       @     �S@     �K@      �?      1@      &@      �?      @      @      @      J@       @     �h@      �?              �?      @      ]@      E@              0@      &@      @      �?              @     �H@      �?     �N@       @      �?      @      @      8@      4@      �?       @                                              @              "@       @                       @      �?      @              �?      &@      @      �?              @      G@      �?      J@              �?      @      @      7@      1@      �?      @      *@              �?      �?      @      E@      @     �`@                      @       @     �Q@      K@              =@      *@              �?      �?      @      A@      @      Y@                      @       @      N@      K@              =@      *@              �?      �?      @      ?@      @     �T@                      @       @     �L@      H@              ;@       @                      �?      �?      &@       @       @                      �?              4@      &@              "@      @              �?              @      4@      @     �R@                      @       @     �B@     �B@              2@                                              @              1@                                      @      @               @                                              �?              @                                       @                      �?                                               @              $@                                      �?      @              �?                                               @             �@@                                      $@                                                                      @              "@                                      @                                                                      �?               @                                      @                                                                      @              @                                       @                                                                      �?              8@                                      @                                                                      �?              *@                                                                                                                              &@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJu�	DhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�I[۷{�?�	           ��@       	                     �?�C�_��?�           �@                           @    ��?�            �@                           @
�+t"�?8           ؋@������������������������       �M��]��?           �z@������������������������       �.Z٢�-�?+           }@                           �?��NO�?T            �`@������������������������       �     ��?&             P@������������������������       �z%�ZV��?.            @Q@
                           @ILֹQ�?q           ؛@                           �?F-<Z�?           @�@������������������������       ���o��?�           x�@������������������������       �d�4���?           �@                            �?\��[�?d            �d@������������������������       �4�Ű��?=            @Y@������������������������       �l������?'            @P@                           �?�]���?�           L�@                           �?�Ű���?�           ��@                           �?�PQ����?�            �p@������������������������       ��2����?:            @V@������������������������       �����2�?t            �f@                          �;@
RԱQq�?�            �v@������������������������       �BGW�i��?�            0t@������������������������       �!�g�1a�?            �E@                           @H^�J�?            p}@                           �?#Y��R�?�            �u@������������������������       �Ê(N:!�??            @Z@������������������������       �������?�             n@                           @�`7l[��?M            @_@������������������������       �A��?�?             K@������������������������       �ͫ���/�?.            �Q@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      ;@     �@@      6@     �V@     H�@      F@     |�@      2@      *@     �V@     �M@     ��@     �@      5@     �o@     �c@      2@      6@      5@     @R@     @~@     �A@     x�@      "@      $@     @S@      I@     �@     �x@      2@     @j@     �G@      @      @      @      3@     @f@      .@      s@       @              7@      (@     `k@      _@      @     �L@      G@      @      @      @      1@     �b@      *@     �o@       @              6@      &@     �i@     @Y@       @      J@      9@      �?       @      @      "@     �T@      @     �]@      �?              @      @      Z@      B@       @      9@      5@      @      @      @       @     �P@      @      a@      �?              .@      @     �Y@     @P@              ;@      �?                               @      >@       @     �I@                      �?      �?      *@      7@      @      @      �?                              �?      8@              .@                                      @      .@              @                                      �?      @       @      B@                      �?      �?      $@       @      @              \@      ,@      1@      ,@      K@      s@      4@     �y@      @      $@      K@      C@      r@     �p@      (@      c@      [@      ,@      ,@      ,@      K@      r@      .@     Pv@      @      $@     �D@     �B@      q@     �m@      (@     �`@      P@      &@      $@      "@      ?@     �a@      &@     �c@      @       @      8@      *@     �_@     �U@      "@      S@      F@      @      @      @      7@     `b@      @      i@      �?       @      1@      8@      b@      c@      @      M@      @              @                      0@      @      L@       @              *@      �?      2@      =@              3@      �?                                      @      @      C@                      @      �?      (@      1@              .@      @              @                      "@              2@       @               @              @      (@              @     �F@      "@      &@      �?      1@     �h@      "@      y@      "@      @      *@      "@      l@      \@      @      F@      B@      @      @      �?      @      ]@      @     �j@      @      @      @       @     @^@     �R@      @      <@      4@       @      @              @     �L@       @      P@      @      �?      @      �?      M@      A@      �?      (@      @               @              @      4@              3@                      @      �?      .@      *@              @      *@       @      @              @     �B@       @     �F@      @      �?                     �E@      5@      �?      @      0@      �?      �?      �?             �M@       @     �b@      @       @      @      @     �O@     �D@       @      0@      .@      �?      �?      �?              I@       @     �^@      @              @      @      M@     �D@       @      0@      �?                                      "@              :@               @                      @                              "@      @      @              $@     @T@      @     �g@       @              @      �?      Z@     �B@              0@       @      @      @               @     �J@      @     �b@                      @      �?      U@      5@               @      @       @                       @      6@       @      :@                      �?             �@@       @              @      @      @      @              @      ?@       @     �^@                       @      �?     �I@      *@              @      �?      �?       @               @      <@      �?      D@       @              @              4@      0@               @                       @              �?      "@              *@                      @              $@      (@              @      �?      �?                      �?      3@      �?      ;@       @              �?              $@      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJKhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �:@|��'֦�?�	           ��@       	                     @�Qq��?H           ��@                          �0@�n0E.�?�           ��@                            �?��
#;S�?k            @e@������������������������       ���p;���?)            @P@������������������������       ��D�=��?B            @Z@                            �?0�P3�?�           ,�@������������������������       ���I�O��?           ��@������������������������       ���!���?o           ��@
                           �?:�����?V           �@                           �?"�87e��?[           ��@������������������������       ��ٴ��?�             k@������������������������       ��oM��z�?�            @v@                           �?���	 ��?�            x@������������������������       �$Vn\1��?|             g@������������������������       ���Ρ@��?             i@                           @�6 �J#�?g           `�@                            @�"�,���?�            �y@                           �?{��hX�?�            �p@������������������������       ����9���?U            �`@������������������������       �s�	U���?P             a@                           @��*ڸH�?Z            �a@������������������������       ��Aռ(��?C            �Z@������������������������       �����[�?             B@                           @���!pc�?h             f@                          �?@��T~F��?=            @Y@������������������������       �:O̖6K�?2            �T@������������������������       �h/�����?             2@                           �?z\�|��?+            �R@������������������������       ���!pc�?	             &@������������������������       �     ��?"             P@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      9@     �H@      7@      ]@     x�@      @@     ̐@      *@      &@      R@     @R@     ��@     �@      5@     �r@     �e@      5@     �D@      6@     �Z@     P�@      ;@     �@      (@      &@     �O@     �P@     ��@     �|@      1@     �o@     �`@      .@     �@@      3@     �U@     0{@      3@     ��@      @       @     �I@      J@     �x@     �s@      .@     @k@      @      �?      �?      @      @      A@      @      2@              �?      @      @      ?@      B@      �?      2@                               @      @      (@      @      @                              �?      2@      0@              @      @      �?      �?      �?      �?      6@              *@              �?      @      @      *@      4@      �?      *@     @_@      ,@      @@      0@     �T@     y@      0@     �@      @      @      G@     �F@     �v@     �q@      ,@      i@     �U@      @      2@      ,@     �J@      t@      (@     P|@      @       @      =@      ;@     �q@     �g@       @      `@      C@      @      ,@       @      >@     @T@      @      W@      @      @      1@      2@     @T@      W@      @     �Q@      E@      @       @      @      3@     �b@       @     �r@      @      @      (@      .@     @j@     `a@       @      B@      ;@              @       @      "@      V@      @      g@      @      @      @      (@     �[@      V@       @      7@      (@              @              @      E@             �P@      �?      @      @      @     �@@      >@              *@      .@              @       @      @      G@      @     �]@      @              @      "@     @S@      M@       @      $@      .@      @      �?      �?      $@     �O@      @     @\@                      @      @      Y@     �I@              *@       @      @              �?      $@      A@      @      E@                      @       @     �B@      :@              &@      @      �?      �?                      =@             �Q@                      �?      �?     �O@      9@               @      0@      @       @      �?      $@     @Y@      @     �j@      �?              "@      @     �\@      J@      @     �E@      *@      @       @      �?       @     �R@      @     �_@      �?              @      @     �W@      >@      @     �@@      "@      @      @      �?      @     �H@      @     �Q@                      @      @     �O@      6@       @      <@      @      @      @              @      1@      @      D@                      @      �?      4@       @       @      6@      @                      �?      �?      @@              ?@                       @       @     �E@      ,@              @      @      �?      @              @      9@              L@      �?                       @      ?@       @       @      @       @              @              @      0@              H@      �?                       @      1@       @              @       @      �?                              "@               @                                      ,@               @              @                               @      ;@       @     �U@                       @      �?      4@      6@              $@      @                                      2@       @      E@                      �?               @      3@               @       @                                      1@       @     �@@                      �?               @      (@               @      �?                                      �?              "@                                              @                                                       @      "@             �F@                      �?      �?      (@      @               @                                       @      @              �?                                       @                                                                      @              F@                      �?      �?      $@      @               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJf,ShG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?T�v�4��?�	           ��@       	                     @i���/�?8           �@                           @Dz��.s�?           ܓ@                           @0�_P�?M           ��@������������������������       �f1s �,�?
           ��@������������������������       �sᮾI��?C             [@                           @�.��|�?�            �u@������������������������       �S����p�?�            �o@������������������������       ����@Y��?6            �V@
                           @����6�?$           �|@                          �2@T,TG?<�?�            �r@������������������������       �����K��?5            �U@������������������������       ���9��Q�?�            �j@                           @N�d�:��?d            �c@������������������������       �>�>��?)             N@������������������������       ��$�zE��?;            �X@                          �;@�=���?o           
�@                            @ �ϓ�?�           ��@                            �?x?r����?�            �@������������������������       ��ٮ�h��?�           p�@������������������������       ����q��?�            @v@                           �?h~�bx�??           p~@������������������������       �֋�ܓ��?3            �T@������������������������       �d�����?           @y@                            @�ߤN6��?�            �q@                           @)�1D]�?s            @g@������������������������       ���fL�?`             c@������������������������       ��"��?            �@@                           @-����?:             Y@������������������������       ����J��?0            �U@������������������������       ��)x9/�?
             ,@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      @@      >@      :@      X@     ��@     �C@     Ȑ@      4@      $@     �Q@     @R@     X�@     x�@      0@     �p@     @X@      3@      :@      &@     �F@     r@      6@     @y@      $@      @      E@     �C@     0t@     �o@       @     �a@     �P@      ,@      7@      &@     �B@     @k@      1@      q@      @      @     �A@     �@@      l@      g@      @      ^@      G@      &@      .@       @     �A@     �c@      @     �j@      @      �?      A@      4@     @e@     �\@      @      W@     �D@      @      .@       @      @@      b@       @     @h@       @      �?      =@      .@      c@     @Y@      @     @R@      @      @                      @      ,@       @      2@      �?              @      @      2@      ,@              3@      5@      @       @      @       @      N@      *@      N@       @       @      �?      *@      K@     �Q@      @      <@      0@      @      @      @      �?      H@      (@      A@      �?       @      �?      "@     �B@     �M@      @      2@      @               @              �?      (@      �?      :@      �?                      @      1@      &@              $@      >@      @      @               @     �Q@      @     �`@      @      �?      @      @     �X@      Q@      �?      4@      1@      @      @              @     �M@      �?     @S@      @              @       @      Q@     �E@              &@      @               @              �?      4@              1@                      �?       @      >@      @              @      ,@      @      �?              @     �C@      �?      N@      @              @              C@      B@              @      *@      �?                      �?      (@      @     �K@       @      �?              @      ?@      9@      �?      "@       @      �?                      �?      @       @      1@                                      $@      $@      �?      @      @                                      @       @      C@       @      �?              @      5@      .@              @     @Y@      *@      @      .@     �I@     �t@      1@     ��@      $@      @      =@      A@     �z@      u@       @     �_@     @W@      &@      @      ,@      H@     @q@      &@     ��@      @      @      7@      @@     �w@     �s@      @     @]@     �S@       @      �?      "@     �D@     �j@      $@     �w@      @      @      6@      :@     pp@     `o@      @     �X@     �I@       @              "@      2@      e@      @      t@       @               @      *@     @j@      e@      @     �O@      <@              �?              7@     �F@      @     �K@      �?      @      ,@      *@     �J@     �T@             �A@      ,@      @      @      @      @     �O@      �?     �f@                      �?      @     @]@     �O@       @      3@      @              @              @      @      �?      ;@                                      *@      2@              "@      $@      @              @      @     �M@             �c@                      �?      @      Z@     �F@       @      $@       @       @              �?      @     �M@      @     �[@      @      @      @       @      F@      8@       @      "@      @       @              �?              ;@      @      Q@      @              @       @      B@      2@       @       @      @       @                              2@      @      N@                      @       @      9@      2@       @       @                              �?              "@               @      @                              &@                               @                              @      @@              E@      @      @                       @      @              �?       @                              @      ?@              B@              @                      @      @              �?                                              �?              @      @                               @       @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ,�tphG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?c�@y\��?�	           ��@       	                     @��� �:�?H           8�@                            �?G���x�?           �@                           @�t%���?           �z@������������������������       ���]��o�?�             t@������������������������       �����2�?;            �Y@                          �:@^P��)��?           ��@������������������������       ���+�:��?�           �@������������������������       ���A��?7            @T@
                           @�� �<�?1           0}@                          �1@4Qev�?�            @w@������������������������       ��8��8��?              H@������������������������       ��Z�~�F�?�            @t@                           @槡}�x�?@            �W@������������������������       � n�r��?1            �R@������������������������       �ffffff�?             4@                            @���ٗ��?^           ��@                            �?��/m���?�           ԗ@                            �?�����?�           �@������������������������       ��2mq"0�?u           ��@������������������������       ��6b�v�?m           ��@                          �>@�!��c�?�            w@������������������������       ��#.(�?�            0v@������������������������       �:/����?
             ,@                           @JR Uw��?�           0�@                           @�������?&           �}@������������������������       �V_`C�?           �|@������������������������       ��������?	             1@                          �;@�:V.���?c            �d@������������������������       ��m�P�?N            ``@������������������������       �B{	�%��?             B@�t�b��      h�h4h7K ��h9��R�(KKKK��h��B�       �l@      @@      =@      9@      ^@     �@      ?@     ��@      7@       @     �S@     �T@     ��@     @~@      2@      p@     @`@      5@      2@      *@     @R@     �r@      4@     0{@      (@      @      =@     �A@     �p@     �m@      @     `a@     �X@      ,@      ,@      (@     �J@     @k@      .@     `r@      $@      @      6@      ?@     �e@     @h@      @     �\@      :@       @      @      @      4@      R@       @     @`@       @              &@      $@     �I@     �H@       @      ?@      7@       @      �?      @      1@      J@       @     �Z@       @              "@      "@      D@      @@      �?      5@      @              @              @      4@      @      8@                       @      �?      &@      1@      �?      $@     @R@      (@      "@      @     �@@     @b@      @     �d@       @      @      &@      5@      _@      b@       @     �T@     �N@       @       @      @     �@@      a@      @     `b@      @      @      $@      5@     �Z@     ``@       @     �S@      (@      @      �?                      "@              1@      �?              �?              2@      ,@              @      ?@      @      @      �?      4@     @T@      @     �a@       @      �?      @      @     �W@     �E@      �?      9@      8@      @      @      �?      2@     �Q@      @     @Y@       @              @      @     �S@     �@@      �?      7@      �?                              @      &@              &@                              �?      @      @              @      7@      @      @      �?      *@     �M@      @     �V@       @              @       @     �R@      :@      �?      0@      @      @                       @      &@      �?      D@              �?      �?      �?      .@      $@               @      @      @                       @       @      �?      ?@              �?      �?      �?      $@      "@               @       @                                      @              "@                                      @      �?                      Y@      &@      &@      (@     �G@     pw@      &@     ��@      &@      �?     �H@      H@     @z@     �n@      *@     �]@     �T@      $@       @      $@     �D@     �p@      $@     �z@      @      �?      E@     �D@     �q@     @g@      $@     �X@     �M@      @      �?       @      6@     �j@      "@      w@      @              9@      4@     `k@     �`@      @      O@      :@      @              @      "@     �]@      @      j@      @               @       @     �Z@     �P@      @      8@     �@@      �?      �?       @      *@     �W@      @     �c@      @              7@      (@     @\@     �P@      �?      C@      7@      @      @       @      3@      M@      �?     �M@      �?      �?      1@      5@      O@     �J@      @      B@      7@      @      @       @      3@      M@      �?      J@      �?      �?      1@      4@      M@     �J@      @     �A@                                                              @                              �?      @              �?      �?      2@      �?      @       @      @      Z@      �?     �p@      @              @      @     `a@     �N@      @      5@      .@              @       @      @     �N@      �?     �i@      @              @      @     �[@      G@              0@      .@              @       @      @      N@      �?     @i@      �?              @      @     �Z@      F@              ,@                                              �?               @      @                      @      @       @               @      @      �?                      �?     �E@             @P@                       @      �?      <@      .@      @      @      @      �?                      �?      :@             �I@                       @      �?      9@      *@      @      @                                              1@              ,@                                      @       @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�6hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @eI����?�	           ��@       	                     @#4B"h��?Y           ,�@                            �?e}��W;�?           �@                           �?pJ�Y��?>           `�@������������������������       �8�gg��?�           �@������������������������       �H����?�            �p@                           �?�>����?�            `u@������������������������       �c���{f�?f            �e@������������������������       ��� �~�?g            �d@
                           �?zyʹ�K�?N           H�@                          �5@�����{�?�            p@������������������������       ��E���-�?[             b@������������������������       �,��i�?L            @\@                          �6@��HJ�}�?�            �p@������������������������       �c`�K�?p            �e@������������������������       �̟�Hr��?7            �V@                            @+�}�?o           ��@                           @	�E����?�           ��@                            �?��/���?G           ،@������������������������       �V�ѩ�A�?�           �@������������������������       ��Q�U���?a             c@                           @�y�J>�?�           x�@������������������������       ��X�jcV�?R           ��@������������������������       �N��4�?M             _@                           �?�5�P��?�           ��@                          �;@�L+\�?D            �Z@������������������������       �7�A��?9             V@������������������������       ��lO���?             3@                           @DM�v+��?E           �~@������������������������       �!߾��?           pz@������������������������       ��|n�k��?,            �P@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      <@     �E@      <@     �Z@     ��@      @@     �@      <@      @      Z@     �P@     І@      �@      <@     �m@     @[@      1@      @@      4@     �J@     0r@      $@     �|@      (@      @     �E@      <@     @w@      g@       @     @X@     �S@      0@      2@      2@     �G@     @j@       @     �q@      $@       @     �C@      9@     �n@      `@       @      S@     �K@      (@      $@      *@      6@     �d@       @     �m@      @              :@      .@     �e@     �U@      @     �E@      H@       @       @       @      3@     @Z@       @     `e@      @              3@      *@     �Z@     @P@      @      ;@      @      $@       @      @      @     �M@             �P@                      @       @     �P@      6@      �?      0@      8@      @       @      @      9@      G@              H@      @       @      *@      $@     �R@      E@      �?     �@@      &@      @      @      @      .@      7@              5@      @       @      @      @      @@      :@      �?      1@      *@      �?      @      �?      $@      7@              ;@                      "@      @      E@      0@              0@      >@      �?      ,@       @      @     @T@       @     �e@       @      �?      @      @     @_@      L@              5@      8@      �?      (@              @     �I@       @     �Q@       @              @             �G@      <@              &@      .@      �?      @              @     �A@      �?     �B@                      @              <@      "@              @      "@              @              �?      0@      �?     �@@       @              �?              3@      3@              @      @               @       @      �?      >@             �Y@              �?              @     �S@      <@              $@      @               @       @      �?      8@              L@                                     @P@      0@              @      @                                      @             �G@              �?              @      *@      (@              @      X@      &@      &@       @     �J@     0w@      6@     ��@      0@      @     �N@     �C@     `v@     �t@      4@     �a@      T@      @       @      @      E@     pp@      3@      z@      (@      @      N@      A@     @m@     p@      .@     @_@      C@      �?      @      @      4@     �c@       @      n@      @       @      C@      "@     �c@     �d@      @      N@      =@      �?      @      @      2@     �^@      @     �k@      @              6@      @     �`@     �a@      @     �F@      "@              �?               @     �@@      �?      3@       @       @      0@       @      7@      :@       @      .@      E@       @      @              6@     �Z@      &@     �e@      @      �?      6@      9@      S@     �V@      "@     @P@     �A@       @      @              3@     @W@      &@      a@      �?      �?      5@      5@      P@     �R@      "@     �D@      @                              @      ,@             �C@      @              �?      @      (@      0@              8@      0@       @      @      �?      &@      [@      @      k@      @              �?      @      _@     �R@      @      1@       @              �?              �?      "@              F@                              �?      3@      3@              @      @              �?              �?      @              @@                              �?      3@      1@              @      @                                       @              (@                                               @                       @       @       @      �?      $@     �X@      @     �e@      @              �?      @     @Z@     �K@      @      (@      @      @       @      �?      $@     �V@      @      c@      @                      @     �U@     �D@      @      &@       @       @                               @              3@                      �?              3@      ,@              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJa��*hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @����(z�?�	           ��@       	                     �?��蟑��?�           ��@                           �?���j��?�           ��@                          �:@2G�����?            z@������������������������       �ӌ���?�             w@������������������������       �9��8���?             H@                          �<@i�0P1�?           ��@������������������������       ��`؈x�?^            �@������������������������       �"~2��?!            �H@
                           @v�P��M�?J           l�@                          �2@_�
��g�?�           @�@������������������������       �;ٝ��?8           0@������������������������       �}JY#�?�           t�@                           @�4��i�?V            `a@������������������������       ���e(A�?E            @\@������������������������       ��q-�T�?             :@                          �7@F5UA*#�?�           �@                          �2@e��K�d�?�           X�@                           �?5���;�?�            �q@������������������������       �� ����?F            @\@������������������������       ��H����?o            �e@                           @ '�	g�?&           �|@������������������������       ����JKI�?�            �v@������������������������       ���|J>l�?8            �W@                           �?��(F0�?�            �x@                           @^6k@I��?a            �d@������������������������       �a㟌�V�?I            �^@������������������������       ��3_<�?             E@                           �?�
e͡��?�            @m@������������������������       ��Œ_,��?             >@������������������������       � �ʹ��?}            �i@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      <@      D@     �A@     �[@      �@      <@     ��@      0@       @     �R@     �K@     �@     �@      2@      p@     �d@      4@      9@      =@     �T@     0}@      5@     p�@      (@      @      P@      I@     �@     �v@      0@     �j@      J@      "@       @      .@      9@     `d@      "@     @s@      @              .@      &@     �k@     @^@      @      J@      5@      @      �?      @      3@     @R@      @     �[@      �?              (@      $@     �R@     �I@       @      =@      5@      @      �?      @      1@     �P@      @     �U@      �?              $@      $@     �Q@     �H@       @      9@                               @       @      @      �?      8@                       @              @       @              @      ?@      @      �?      $@      @     �V@      @     �h@      @              @      �?     �b@     �Q@       @      7@      ?@      @      �?      $@      @      V@      @     �e@                      @      �?     �`@     �P@       @      7@                                               @              9@      @                              0@      @                     @\@      &@      7@      ,@     �L@      s@      (@     �y@       @      @     �H@     �C@     0r@     �n@      (@      d@     @\@      &@      6@      ,@      L@      q@      &@     �v@      @      @      G@     �A@     q@     �l@      (@      b@      I@      �?      "@      @      ,@     �T@      �?      T@      �?      @      7@      5@      T@     �S@       @     �E@     �O@      $@      *@      "@      E@      h@      $@     �q@      @      @      7@      ,@      h@     �b@      @     @Y@                      �?              �?      >@      �?     �G@       @              @      @      2@      0@              0@                      �?              �?      9@      �?     �D@       @              @      @      (@       @              .@                                              @              @                                      @       @              �?      L@       @      .@      @      =@     �e@      @      z@      @      �?      $@      @     �k@     �a@       @      G@      9@      @      *@      @      5@     �_@      @      o@       @      �?      "@       @      e@     @U@              ?@      "@       @      @      �?      $@      E@       @     @V@                      @      �?      U@      ;@              *@      @              @                      *@             �@@                                     �H@       @              @      @       @      �?      �?      $@      =@       @      L@                      @      �?     �A@      3@              "@      0@       @      "@      @      &@      U@      @     �c@       @      �?      @      �?      U@      M@              2@      0@       @      "@      @      @      N@      @     �^@       @      �?              �?      T@      H@              &@                                       @      8@              B@                      @              @      $@              @      ?@      @       @               @     �G@      �?     @e@       @              �?      @     �K@     �L@       @      .@      4@      �?       @              @      1@      �?      M@      �?              �?              7@      9@       @       @      4@               @               @      .@      �?     �E@      �?              �?              &@      6@       @       @              �?                      @       @              .@                                      (@      @              @      &@      @                      @      >@              \@      �?                      @      @@      @@              @                                      �?      @              (@                                      �?      $@                      &@      @                       @      8@              Y@      �?                      @      ?@      6@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJk�'hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�рn�?�	           ��@       	                    �?8ӣ�o��?           ��@                            @f�͞�?�            �@                          �3@��?�x��?           0{@������������������������       ��S����?�             i@������������������������       �2�����?�            @m@                           �?�F1'
U�?m            �e@������������������������       ���[��?;            �Y@������������������������       ����IP��?2            �Q@
                            @rx��?x           (�@                            �?�햸���?           `z@������������������������       ��;�*B�?�            �s@������������������������       ���N��N�?I             Z@                          �2@�q��?`            �c@������������������������       �M����?&            @P@������������������������       �D�A�@1�?:            �W@                            @���W�%�?�           H�@                            �?L)T֋�?�           �@                           �?r)S�?�           x�@������������������������       ��ȸ���?p           p�@������������������������       �X�x�N6�?-           ��@                           @⡅����?           �y@������������������������       ���P
�?�            �u@������������������������       �߼�xV�?*             N@                           @O�o7���?�           X�@                           �?�=x��?l           ��@������������������������       �ܶm۶=�?�             l@������������������������       ���y&4�?�            �w@                          �0@�߽�?�            `j@������������������������       ��G�z��?             $@������������������������       �%|�y��?�             i@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @h@      A@      C@      7@     @[@     �@     �A@     ԑ@      4@      "@     @R@     �Q@     X�@     H�@      2@     �m@     �R@      @      0@      &@      A@     @g@      @     �r@      $@       @      =@      ;@      m@     �d@      @     �U@      A@      @      ,@      @      9@     �Y@      @      a@      @       @      3@      2@     �W@     @T@      @     �J@      :@      @      &@      @      5@     @R@      @     @U@      @       @      ,@      1@     �O@      P@      @     �B@      @       @      "@       @      2@      8@       @     �E@      �?       @      @      @      9@     �C@      �?      .@      4@      �?       @      @      @     �H@      �?      E@      @               @      &@      C@      9@       @      6@       @      @      @              @      >@       @      J@                      @      �?      @@      1@              0@      @              @               @      ,@       @     �D@                              �?      ,@      (@              $@      @      @                       @      0@              &@                      @              2@      @              @     �D@      �?       @      @      "@     �T@             @d@      @              $@      "@     @a@     �T@       @     �@@     �B@      �?       @      @       @      R@             �X@      @              $@      @     @V@     �N@       @      ;@      =@                      @       @     �M@             @U@      @               @       @      N@      J@              ,@       @      �?       @      �?      @      *@              ,@                       @      @      =@      "@       @      *@      @                              �?      &@             �O@                              @     �H@      6@              @      @                                      @              6@                                      <@      @              �?      �?                              �?      @             �D@                              @      5@      .@              @     �]@      ;@      6@      (@     �R@     p|@      >@     P�@      $@      @      F@      F@     �@     Pv@      *@      c@     �U@      3@      (@      (@      M@     pr@      5@     X�@      $@      @      D@      @@      u@     �q@      "@     ``@     @P@      ,@      @      $@     �C@     @m@      ,@      }@      @       @      8@      4@     �q@     �k@      @     �V@      A@      @      @      @      :@     �X@      @      a@      @       @      (@      (@     �]@     �T@      @     �D@      ?@      $@      �?      @      *@     �`@      "@     pt@      @              (@       @     �d@     `a@      �?      I@      6@      @      @       @      3@     �N@      @     �V@      @      @      0@      (@      J@     �P@      @      D@      5@      @      @       @      0@      K@      @     @P@      @      @      $@      (@      H@     �M@      @     �A@      �?              �?              @      @              :@                      @              @      @              @      @@       @      $@              1@      d@      "@     �q@                      @      (@      f@     �Q@      @      6@      ?@      @      "@              .@     @]@      @     `g@                      @      (@      a@      J@      @      4@      5@      @      @              &@     �F@       @     �H@                       @      @      D@      9@       @      *@      $@      @      @              @      R@      @     @a@                       @       @      X@      ;@       @      @      �?      �?      �?               @     �E@      @      Y@                                      D@      2@               @                                              @      @       @                                       @                              �?      �?      �?               @      D@             �X@                                      C@      2@               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�� MhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?��}(|�?�	           ��@       	                     @ߎ��(�?\           p�@                           @� �(S{�?$           ��@                            �?6& ���?A           ��@������������������������       �����"`�?�            �@������������������������       ���s�?�            �i@                           @��[�_��?�            �u@������������������������       ��[{��?`             c@������������������������       ���bS��?�            �h@
                           �?o��3��?8           �~@                           �?lן=5W�?�            `p@������������������������       �r�q'�?C             X@������������������������       ��:���?c            �d@                           �?BvD��?�            �l@������������������������       ���� �?2            �Q@������������������������       �����?`             d@                          �;@Z �b��?R           ڠ@                           !@d��uG��?�           ��@                            @"PQF��?�           \�@������������������������       ��}Ƞ��?L            �@������������������������       ��c�A#V�?[           x�@������������������������       ��q�q�?             (@                            �?D��T��?�            �p@                           @     ��?2             X@������������������������       �]�i��n�?'            �R@������������������������       �Y�����?             6@                            �?7g����?q            @e@������������������������       ���?��?-            �P@������������������������       ��TȲ��?D            �Y@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@      6@     �F@      <@     @[@     8�@      <@     �@      4@      @     �Q@     �R@     �@     @�@      1@     pq@      [@      (@      ?@      &@     �N@     �s@      1@     �y@      $@      @      :@     �D@     �r@     `p@      @      b@     �T@      @      6@      &@      H@      l@      .@      q@      "@      @      8@      A@     `h@     �g@      @      ^@     �M@      @      1@      &@      @@     @d@      &@      g@       @       @      5@      ;@     �c@     @_@      @     �U@      I@      @      1@      &@      2@     ``@      @     @c@      @              *@      1@     �_@     �V@       @      N@      "@      �?                      ,@      ?@      @      >@      @       @       @      $@      ?@      A@      �?      ;@      7@              @              0@     �O@      @     �V@      �?       @      @      @      C@     �O@       @     �@@      "@              @              @      ?@      �?     �D@      �?      �?      �?      @      .@      8@       @      1@      ,@               @              (@      @@      @     �H@              �?       @      @      7@     �C@              0@      :@      @      "@              *@     @V@       @     �a@      �?               @      @     @Y@     �R@              8@      7@              "@              @      F@             @Q@      �?              �?      @      I@     �G@              "@      @              @              @      ,@             �A@                              �?      2@      *@              @      3@              @               @      >@              A@      �?              �?      @      @@      A@              @      @      @                       @     �F@       @     �Q@                      �?      @     �I@      ;@              .@      @      @                      �?      3@              (@                                      .@      &@              @              �?                      @      :@       @     �M@                      �?      @      B@      0@              $@     @W@      $@      ,@      1@      H@     �t@      &@     ��@      $@       @      F@     �@@     Py@      p@      (@     �`@     �V@       @      ,@      .@     �E@     �q@      "@     `�@      @       @      E@      >@     �v@      n@      &@     �^@     �V@       @      ,@      .@     �E@      q@      "@     X�@      @       @      E@      >@     �v@     �m@      &@     @^@      R@      @      $@      &@      D@     �h@       @      x@      @       @      C@      8@      o@      h@      @      [@      2@       @      @      @      @     �R@      �?      m@      �?              @      @      \@      G@      @      *@                                               @              �?                                               @              �?      @       @               @      @     �J@       @      \@      @               @      @     �F@      2@      �?      *@      �?                                      "@             �F@       @              �?       @      3@      (@              @      �?                                      "@             �@@                      �?       @      &@      (@              @                                                              (@       @                               @                               @       @               @      @      F@       @     �P@      @              �?      �?      :@      @      �?       @      �?       @               @              7@              2@      �?              �?              &@      @              @      �?                              @      5@       @     �H@       @                      �?      .@       @      �?      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ2��XhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?I��M���?�	           ��@       	                    �?�~ηXF�?S           Ԛ@                            �?˵����?�            @n@                            �?��#Y���?S            @^@������������������������       �����(�?0            @R@������������������������       ��qǱ�?#             H@                          �2@�!'�F�?Q            @^@������������������������       ���?��?             :@������������������������       �0�F����??            �W@
                          �=@ J��I�?�           �@                          �1@N��B�?�           �@������������������������       �-2����?�            �p@������������������������       ��T��
�?�           ��@                           @�-��9P�?-            @R@������������������������       �,x4T��?"            �K@������������������������       �n�����?             2@                           @C���?Z           (�@                           �?=VFr��?I           ��@                           �?�Fw����?�           ��@������������������������       ����	���?g           `�@������������������������       �l�ˮ���?R            �`@                            @[n�n��?�            �l@������������������������       �|}p�i�?e            @d@������������������������       ��_�}2�?+             Q@                           !@�DH�%�?           ��@                           �?�+7g.�?	           ��@������������������������       �`����]�?u            �f@������������������������       �nXt(�7�?�           �@������������������������       �*D>��?             *@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      E@     �F@      4@      \@     P�@      E@     ��@      2@      @     �P@     �P@     p�@     p�@      6@     �n@      Z@      9@      @@      @      R@     �s@      9@     �x@      &@      @     �A@      ;@      s@     �l@      "@      ^@      .@      @      @      �?      @      9@      �?     @R@       @              *@      @     �F@      >@              3@      $@      �?      �?      �?      @       @      �?     �C@      �?              (@      �?      1@      ,@              $@      @      �?                              @      �?      ;@                      "@      �?      &@      "@              @      @              �?      �?      @      @              (@      �?              @              @      @              @      @       @      @               @      1@              A@      �?              �?      @      <@      0@              "@                                      �?       @               @                      �?      @      @      �?              �?      @       @      @              �?      "@              :@      �?                              9@      .@               @     @V@      6@      <@      @     @P@     Pr@      8@     �s@      "@      @      6@      7@     Pp@     �h@      "@     @Y@     @T@      6@      <@      @     �K@      r@      8@     �r@      @      @      6@      6@     �n@      g@      "@     �X@      .@      @      @       @      (@     �G@       @      C@               @      @      @      H@     �G@      @      >@     �P@      2@      8@      @     �E@     `n@      0@     Pp@      @      @      2@      1@     �h@     @a@      @     @Q@       @                              $@      @              4@       @                      �?      ,@      *@               @      @                              $@      @              ,@       @                      �?      &@       @               @      @                                                      @                                      @      @                     �Y@      1@      *@      *@      D@     �v@      1@     ��@      @      �?      @@      D@     �{@     �r@      *@     �_@      J@      @      "@      @      1@     �b@      @     �q@       @              ,@      *@      j@     �Y@      @     �I@     �D@      �?      @      @      (@     �]@      @     `k@       @              &@      &@     �a@     �T@      @      @@      @@              @      �?      $@     @W@       @      e@       @               @      $@     �]@     �R@      @      ;@      "@      �?               @       @      :@      �?     �I@                      @      �?      8@       @              @      &@      @      @       @      @      ?@             �O@                      @       @     �P@      4@              3@      &@      @               @      @      6@              C@                       @      �?      F@      .@              2@                      @                      "@              9@                      �?      �?      7@      @              �?     �I@      (@      @       @      7@     �j@      ,@      x@      @      �?      2@      ;@     `m@     `h@      "@     �R@     �I@      (@      @       @      7@      j@      ,@     �w@      @      �?      2@      ;@     `m@     @h@      "@     �R@      @               @       @      @      0@      @     �N@                      @              ?@      E@       @      @      H@      (@       @      @      0@      h@       @     �s@      @      �?      .@      ;@     �i@      c@      @      Q@                                              @              @                                              �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���`hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�B�ܖ�?�	           ��@       	                    @�{�a�?6           (�@                           �?4��_��?�           �@                           �?h �T�7�?}           ��@������������������������       ��r���?�             m@������������������������       ��*��?;�?�            �v@                            �?*}r���?           �z@������������������������       ��z�<p�?�            @p@������������������������       �_�7���?l            �d@
                           �?Hdc�S�?�           8�@                            �?3+4�!v�?�            �q@������������������������       �#""�?W            �c@������������������������       �J�L�� �?H            �^@                            @+����?           �z@������������������������       �V6d�F�?�            0v@������������������������       �V�\j�?/            �R@                            @��c�?T           ��@                           @�����?�           ��@                            �?~g>]��?�           @�@������������������������       �}	`x(�?5           `�@������������������������       �g>]{x��?�            @r@                           @�9`�E�?�            �u@������������������������       ���c> ��?�            @o@������������������������       ������?<            �W@                           @��<��&�?�           ��@                           �?g�L���?'            ~@������������������������       ��N$���?�            �t@������������������������       �60���?a            �b@                           �?�[��?h            �f@������������������������       �=�
I��?             3@������������������������       ��.�/�U�?Y            @d@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@     �C@     �D@      8@     �V@     ��@     �@@     �@      4@       @     �R@     �L@     @�@     ��@      5@     �o@     �Y@      ;@      <@      @      I@     �u@      0@     �w@      (@      @      ;@      ?@     �t@      l@      $@     �`@     @P@      6@      6@      @      8@      l@      &@     @l@      "@              .@      "@     �f@      `@      @      T@      F@      &@      3@      @      (@      `@      @     �`@       @              &@      @      X@     �R@      @      I@      (@              @      �?      @      E@      �?     �N@      @              @      @     �D@      ;@       @      3@      @@      &@      .@       @      @     �U@       @     �Q@      �?              @       @     �K@     �G@       @      ?@      5@      &@      @      �?      (@     @X@       @     �W@      �?              @      @     @U@     �K@      �?      >@      0@       @       @      �?      @      N@      @      K@      �?              @      @      O@      <@      �?      0@      @      "@      �?               @     �B@      �?      D@                      �?      �?      7@      ;@              ,@      C@      @      @      @      :@     �_@      @     �c@      @      @      (@      6@      c@      X@      @     �J@      7@      �?      @       @       @      I@       @     �H@       @       @      @      @      M@      D@      @      9@      0@              @      �?      @      >@              C@       @              �?       @      9@      1@              0@      @      �?      �?      �?      �?      4@       @      &@               @      @      @     �@@      7@      @      "@      .@      @      �?      �?      2@      S@      @     �Z@      �?      �?       @      .@     �W@      L@       @      <@      .@      @      �?              0@      L@      @      T@      �?      �?       @      .@     �R@     �J@       @      :@              �?              �?       @      4@              ;@                                      3@      @               @     �W@      (@      *@      1@      D@     0u@      1@     (�@       @      @      H@      :@     �}@     �r@      &@     @^@      S@      "@      &@      &@      A@     `m@      0@     0x@      @      @     �G@      6@     0t@     �k@      $@      Y@      Q@      "@      @       @      3@      g@      $@     �q@      @      @     �C@      0@     @o@     �g@       @     �Q@      G@      @      @      @      $@     �a@      @     �m@       @              6@      &@      i@      a@      @     �G@      6@      @      @      @      "@     �E@      @      G@       @      @      1@      @     �H@      K@      @      7@       @              @      @      .@     �I@      @      Z@      �?               @      @     @R@     �@@       @      >@      @              @      @      &@     �C@      @     @T@      �?              @      @     �L@      ,@       @      1@       @                              @      (@              7@                       @      @      0@      3@              *@      3@      @       @      @      @      Z@      �?      p@      @       @      �?      @      c@      T@      �?      5@      "@      @       @      @      @     �P@      �?      i@      @       @      �?      @      \@      H@              3@      @      @      �?      @      @      H@      �?     �a@      @       @      �?      @     �O@      >@              2@      @              �?                      3@              N@                                     �H@      2@              �?      $@                              �?     �B@             �L@                              �?      D@      @@      �?       @      @                              �?      @               @                                      �?      "@                      @                                      A@             �K@                              �?     �C@      7@      �?       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ&�0hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @��5΀�?�	           ��@       	                    �?��u��?�           �@                           @���c_�?           ��@                          �=@�D�K�?�           h�@������������������������       ��kiP|\�?�           ԑ@������������������������       ����~ӝ�?            �B@                          �8@��`d���?8            �U@������������������������       �D��H��?+            �P@������������������������       ��������?             4@
                          �;@��h�V��?�            �@                           @�rh4��?_           ��@������������������������       ��m�Ш�?�           ��@������������������������       �a$�o��?�           ��@                           �?@���5��?n            �d@������������������������       �x�5?,R�?             B@������������������������       �"Y^��?Y             `@                          @@@E����?�           D�@                           @H��*��?�           ��@                           �?������?c           p�@������������������������       ��d�,�?           �x@������������������������       �j*,LL��?a           ��@                           �?<!t����?V            �^@������������������������       �z���2�?            �E@������������������������       �\���(�?7             T@                          �@@��Q��?             D@������������������������       �����Gc�?
             3@                          @A@�ՙ/�?             5@������������������������       �H�z�G�?             $@������������������������       ����!pc�?             &@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `i@      B@     �C@      >@     �[@     ��@     �A@     @�@      ,@      "@     @P@     �G@     ��@     ؀@      7@      o@     �c@      ;@      ?@      9@     @W@     P@      ;@     Ѕ@      &@      @     �L@     �A@      @     Py@      5@      k@     @R@      .@      3@      *@      L@      l@      .@     �q@       @      @      9@      4@     �i@     �g@      $@      Y@      Q@      .@      .@      *@     �G@     �j@      (@     �p@       @      @      9@      4@     �g@     �f@      $@     @U@     �P@      .@      .@      *@      F@     `j@      (@      o@       @      @      9@      4@     �g@      f@      $@     �T@       @                              @      @              5@                                       @      @               @      @              @              "@      &@      @      .@                                      .@      "@              .@      @              @              "@      @      @      @                                      ,@      "@               @                                              @               @                                      �?                      @      U@      (@      (@      (@     �B@     @q@      (@     �y@      @       @      @@      .@     @r@     �j@      &@      ]@     @T@      $@      (@      &@     �A@     �n@      $@     Pv@      �?       @      =@      (@     `p@      i@      $@      Y@      J@       @       @       @      2@      [@      @     �d@                      $@      @     �_@      Q@      @      F@      =@       @      @      "@      1@     @a@      @     �g@      �?       @      3@      @      a@     �`@      @      L@      @       @              �?       @      >@       @      L@       @              @      @      >@      ,@      �?      0@       @      �?                              $@              @                               @       @      @              @      �?      �?              �?       @      4@       @      J@       @              @      �?      6@      $@      �?      &@      G@      "@       @      @      2@     �g@       @     `y@      @      @       @      (@     �k@     �`@       @     �@@     �F@      "@       @      @      1@     �f@       @     �w@      @       @       @      (@      k@     �`@       @      ?@     �D@      @       @      @      ,@     �c@      @     �u@       @       @      @      &@     �h@     @]@       @      :@      ;@      @      @              "@      Q@      @      ^@      �?       @      �?      @     �T@     �I@      �?      ,@      ,@      �?       @      @      @      V@       @      l@      �?              @      @      ]@     �P@      �?      (@      @      @               @      @      ;@      �?      C@      �?              @      �?      2@      1@              @      @                              �?      @              $@                              �?      @      &@               @              @               @       @      4@      �?      <@      �?              @              &@      @              @      �?                              �?      @              8@              �?                      @                       @                                      �?      @              $@              �?                                               @      �?                                                      ,@                                      @                              �?                                                      @                                      @                                                                                       @                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���4hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @A�ھ�g�?�	           ��@       	                    �?��$
.��?�           :�@                          �?@�ƆgV�?�           p�@                           �?&L�"�h�?�           �@������������������������       �ͬ����?�            �t@������������������������       �����&�?%           ��@                           �?x�5?,�?             ;@������������������������       �f�t���?             1@������������������������       ���(\���?             $@
                          �2@s���p�?�           �@                            �?��O,���?�            0x@������������������������       �P���y �?�            �q@������������������������       ��� i�?=            @Y@                            �?�[���(�?�           ��@������������������������       ������?H           ��@������������������������       �O]Ķ��?�            �p@                           �?-�޷��?�           ��@                           @��ꏊ��?+           `}@                          �9@�Zw���?�            �u@������������������������       ��H�9�?�             q@������������������������       ���t�n�?/            �S@                           @"�jݨ��?L            �]@������������������������       �`!8�e|�?;            �V@������������������������       �bΊx��?             =@                          �;@�&�˝�?{           ��@                           @#P�M��?K           X�@������������������������       ����ӵ�?�            �x@������������������������       �     v�?R             `@                           �?L�����?0            �R@������������������������       ���ͦ-��?              K@������������������������       ��U̠ç�?             5@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@     �@@      ?@      5@     �U@     h�@      5@     ��@      0@      @     �W@     �N@     ��@     ��@      1@      o@      e@      6@      8@      4@     �O@     P~@      3@     `�@      *@      @      U@      I@     ��@     �z@      ,@     �i@      T@      $@      1@      (@     �D@     �k@      (@     Pq@      "@       @      @@      <@     `i@     `h@      @      Y@     �S@      $@      1@      (@     �D@     �j@      (@     Pp@      "@       @      @@      <@     `i@      h@      @      Y@      0@      @      $@      @      (@     �H@       @     �Q@      @              1@       @      A@      J@      @      G@     �O@      @      @      "@      =@     �d@      $@     �g@      @       @      .@      4@      e@     �a@       @      K@      �?                                      @              0@                                              @                                                              @               @                                               @                      �?                                                       @                                              �?                     @V@      (@      @       @      6@     �p@      @     p{@      @       @      J@      6@     Pt@      m@      "@     �Z@      ?@      �?       @       @      @      V@              U@                      1@       @      N@     �N@      @      6@      :@      �?               @      @      Q@             �R@                      @      @     �K@     �B@              $@      @               @               @      4@              $@                      (@      @      @      8@      @      (@      M@      &@      @      @      0@      f@      @     0v@      @       @     �A@      ,@     �p@     `e@      @     @U@     �D@       @      @      @      (@     �b@      @     �r@      @              7@      *@     �i@      `@      @      H@      1@      @      �?              @      <@      @      K@      �?       @      (@      �?      N@      E@             �B@      C@      &@      @      �?      8@      i@       @     �y@      @              &@      &@     �h@     @[@      @     �D@      7@      "@      @              $@     �Y@       @     �b@      @               @      @      T@      L@              1@      5@       @      @              @     �S@      �?     �Z@      @              @      @      M@      F@              *@      0@      @      @              @     �Q@      �?     �Q@       @              @      @      G@      @@              (@      @      @      �?              �?      @              B@      �?                              (@      (@              �?       @      �?                      @      8@      �?     �F@                      @              6@      (@              @       @      �?                       @      4@              ?@                      �?              5@      "@              @                                      �?      @      �?      ,@                      @              �?      @              �?      .@       @      @      �?      ,@     �X@             p@                      @      @     �]@     �J@      @      8@      ,@       @      @      �?      $@      U@             �j@                      @      @     @[@     �I@      @      7@      &@              @      �?      $@      K@             �d@                       @      @     �V@     �C@              .@      @       @                              >@             �H@                      �?       @      2@      (@      @       @      �?                              @      ,@             �E@                                      $@       @              �?      �?                              @       @              B@                                      @                      �?                                      �?      @              @                                      @       @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�;&hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�)��#s�?�	           ��@       	                    @��8��?           ��@                           @��;����?R           ��@                            �?&hOBh��?7           2�@������������������������       ��f��P�?�           ��@������������������������       ���:���?]           `�@                           �?�{���w�?            �F@������������������������       �ƵHPS!�?             *@������������������������       �      �?             @@
                           �?���ȫ��?�           ��@                          �1@*�����?�            @l@������������������������       ��V���?             6@������������������������       �3����?�            �i@                           @*گT��?           �z@������������������������       �З`1��?�            �p@������������������������       ���밆:�?i             d@                          �;@���a���?�           ̑@                           �?�^�RA�?w           P�@                           @I��n�5�?           �z@������������������������       ����F�'�?�            �r@������������������������       ��U/�?P            ``@                          �2@�Ͻ��X�?i           ��@������������������������       ����@^�?a            �c@������������������������       �g\�5��?            z@                           @�y�~���?S             a@                           �?�o,���?'            @R@������������������������       �"?ӧ
��?             ?@������������������������       �Bu��?             E@                          �>@     8�?,             P@������������������������       ��=F?�!�?             E@������������������������       �F]t�E�?             6@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@     �C@     �B@      9@      Z@     ��@     �B@     p�@      3@       @     @S@     �L@     �@     �@      $@     @n@     @a@      >@      <@      8@     �T@     �}@      =@      �@      0@      @     �P@     �H@     `@     �y@      @     `i@     �]@      8@      3@      7@      Q@     w@      1@     h�@      &@      @      G@      C@     �x@     q@      @     @c@     @]@      8@      3@      4@      Q@     �v@      1@     ��@      &@      @      G@      B@      x@      q@      @     �b@     �S@      0@      (@      (@      E@     0r@      "@      {@      "@              ;@      4@     `r@      g@      @     �U@     �C@       @      @       @      :@      S@       @     �X@       @      @      3@      0@      W@      V@              P@      �?                      @               @              ;@                               @      @      �?              @                              @               @               @                               @      @                      �?      �?                                                      9@                                      @      �?               @      4@      @      "@      �?      .@     @[@      (@     `b@      @      �?      4@      &@     �[@     �a@             �H@       @      �?      "@               @     �D@      @     �L@      @      �?      "@      @      >@      B@              5@       @              @                      @      �?       @       @                               @      @                      @      �?      @               @     �B@       @     �K@       @      �?      "@      @      <@      ?@              5@      (@      @              �?      *@      Q@      "@     �V@      �?              &@      @      T@     @Z@              <@      @      @                      @     �D@      @     �D@                      "@      @      L@      T@              (@      @                      �?      @      ;@       @     �H@      �?               @       @      8@      9@              0@     �I@      "@      "@      �?      5@      h@       @     �y@      @       @      &@       @     �m@     ``@      @     �C@     �D@      "@      "@      �?      4@     `d@       @     u@      @      �?      &@       @     �l@     @_@      �?     �B@      7@      @      @      �?      (@     �T@      @     �^@       @      �?      @      @     �U@      L@              2@      .@      @      @      �?      &@      N@      @     @T@                      @      �?     �O@     �D@              $@       @      �?       @              �?      6@       @     �D@       @      �?      �?      @      8@      .@               @      2@      @       @               @     @T@      @     �j@      �?              @      @     �a@     @Q@      �?      3@      @               @               @      8@             �C@                      @             �L@      4@              @      *@      @                      @     �L@      @      f@      �?               @      @      U@     �H@      �?      .@      $@                              �?      =@             �R@              �?                       @      @      @       @      @                              �?      $@             �H@              �?                       @       @              �?      @                                      @              .@                                      �?       @              �?                                      �?      @              A@              �?                      �?                              @                                      3@              :@                                      @      @      @      �?       @                                      .@              1@                                      @      @              �?      �?                                      @              "@                                      @              @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�|�ThG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             @*���v��?�	           ��@       	                     @�����?C           ��@                            �?f[�È�?3           >�@                           �?Jk��9��?�           X�@������������������������       �i�J`��?�            px@������������������������       ��<[���?�            @v@                          �<@>��j��?J           Д@������������������������       ���Uvx��?           ��@������������������������       ��qec8��?1            �R@
                           �?��q�m�?           ��@                           @h��.<�?�            Px@������������������������       ���v��S�?�            �p@������������������������       ��P�r�^�?O             _@                           @	�䂐��?           0{@������������������������       ���#�;�?�            �u@������������������������       ��F��s��?:            �V@                          �;@pL��?�           ��@                           �?�щ����?<           �@                            @tܟ�Q�?�            `x@������������������������       �����C�?�            �s@������������������������       �u#�����?2             S@                           @O��?A           p@������������������������       �R]Kܺ�?�            �w@������������������������       ������?P             _@                          �@@& Q����?N            @]@                            �?���	�?F            �Y@������������������������       ��?���0�?(            �M@������������������������       �ˠT�x�?             F@������������������������       �>4և���?             ,@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      D@      =@      8@      Y@     ��@      B@     P�@      *@      "@     @R@     @Q@     p�@     (�@      7@     `r@      e@      ?@      5@      1@     �T@      �@      5@     `�@       @      @     �J@      I@     �@     �t@      0@     �l@     �`@      :@      .@      .@     �Q@     �v@      ,@     P@      @      @     �G@      D@      x@     �o@      .@     �g@      D@      @      �?      @      4@     �a@      "@      m@                      &@      $@      b@     �R@      @      E@      >@              �?      @      @     �T@      @     �`@                      @      $@     �N@      @@      @      2@      $@      @              @      ,@      N@       @      Y@                       @              U@     �E@      @      8@     @W@      5@      ,@      "@      I@     �k@      @     �p@      @      @      B@      >@     �m@     `f@       @     �b@     �U@      1@      *@      "@     �H@     �h@      @     �o@      @      @     �@@      <@     @m@     �e@      @     �a@      @      @      �?              �?      8@      �?      *@      �?              @       @      @      @      �?       @      B@      @      @       @      (@     `b@      @     pq@       @              @      $@      h@     @S@      �?     �D@      8@      @      @       @       @     @S@      @      Y@                      @       @      V@      H@      �?      8@      5@      �?      @              @      L@      @      Q@                       @       @     �H@      D@      �?      ,@      @       @      �?       @      @      5@              @@                      @             �C@       @              $@      (@       @       @              @     �Q@      @     `f@       @              �?       @     @Z@      =@              1@      "@       @                      @     �J@             �b@       @              �?      @     �S@      5@              1@      @               @                      1@      @      =@                               @      :@       @                      ;@      "@       @      @      2@      g@      .@     �p@      @      @      4@      3@     �e@     @g@      @     �O@      :@      "@       @      @      1@     �d@      .@     `j@      @      @      2@      2@      c@      e@      @      N@      3@      @      @      �?       @     �V@      $@     @Q@      @      @       @      0@     �O@     �O@      @      7@      2@      �?      @      �?      @      T@      $@      E@      @       @      @      ,@     �H@     �J@      @      6@      �?       @      �?              �?      $@              ;@      �?       @      @       @      ,@      $@              �?      @      @       @      @      "@      S@      @     �a@      �?      �?      $@       @     @V@     �Z@      @     �B@      @      @       @      @       @      P@      @     �Z@      �?      �?      @      �?      R@     �T@      @      4@      @       @                      @      (@      �?     �A@                      @      �?      1@      7@              1@      �?                              �?      2@             �J@                       @      �?      5@      1@              @      �?                              �?      2@              I@                       @              4@       @              @                                      �?      @              :@                       @              2@      @              �?      �?                                      *@              8@                                       @       @               @                                                              @                              �?      �?      "@                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ4��4hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?��H4��?�	           ��@       	                    �?���?H           ��@                            �?*���-�?�           �@                          �3@�:m�Z��?q            �f@������������������������       �_j�����?.             S@������������������������       �I'��)�?C            �Z@                           �?�� m��?N           P�@������������������������       ��rO���?;            @������������������������       ��8��8��?             8@
                          �=@@�[���?�           ��@                           @n�;���?h           p�@������������������������       �M�+���?g           Ȃ@������������������������       �E!�'�?           Py@                           @��?��?!             J@������������������������       �/�5���?            �D@������������������������       �}��7�?             &@                           �?�����?W           ̠@                            @�aWg&�?t           p�@                          �4@�����?           �|@������������������������       ���|�(<�?�            �k@������������������������       ��+�l��?�            �m@                           @��J�3+�?Y            @`@������������������������       ��E��_��?S            �]@������������������������       ��zv��?             &@                           !@�BLy��?�           `�@                          �;@�w��$��?�           8�@������������������������       �R®�*�?N           ��@������������������������       ��:
�f��?�            @m@������������������������       �p=
ףp�?             $@�t�b�+     h�h4h7K ��h9��R�(KKKK��h��B�       �l@      5@      =@      1@     �]@     `�@      ;@     ��@      .@      *@      Q@     �O@     ��@     �@      0@     �p@      \@       @      7@      @     �P@     �v@      *@     �y@      $@      @      D@     �A@     pr@     �l@      "@      a@     �C@       @      ,@      @      9@     �b@      @     @c@      @       @      6@      0@     �^@      S@       @     �P@      ,@              �?               @     �F@              L@                      @       @     �@@       @      �?      0@      @              �?              �?      $@              <@                              �?      2@      @              @      "@                              �?     �A@              <@                      @      �?      .@       @      �?      $@      9@       @      *@      @      7@     �Z@      @     �X@      @       @      1@      ,@     �V@      Q@      �?      I@      9@      �?      (@      @      4@      Z@      @     @V@      @       @      0@      ,@      U@     �P@      �?      I@              �?      �?              @       @              "@                      �?              @      �?                     @R@      @      "@       @     �D@     @j@      "@     0p@      @      @      2@      3@     �e@      c@      @     �Q@      P@      @      "@       @     �A@     �i@      "@      n@      @      @      2@      3@      e@     �a@      @      Q@     �D@       @      @       @      .@     �a@      @      `@      @      �?      @       @      ]@     �V@      @     �A@      7@      @      @              4@     �P@      @      \@       @      @      .@      &@     �J@      J@      @     �@@      "@                              @      @              3@                                      @      $@               @      @                              @      @              2@                                       @      @              �?      @                                                      �?                                      �?      @              �?     �]@      *@      @      &@     �J@     0v@      ,@     ��@      @      @      <@      <@     �{@     0q@      @     �`@     �F@               @              0@     @U@             @c@      �?              @      ,@     `c@     �R@              D@      F@               @              .@     �R@              [@      �?              @      (@     @[@      M@             �@@      9@                              @     �G@              L@                              @     �G@      3@              3@      3@               @              (@      ;@              J@      �?              @      @      O@     �C@              ,@      �?                              �?      &@              G@                               @      G@      0@              @                                      �?       @              F@                                     �E@      0@              @      �?                                      @               @                               @      @                             �R@      *@      @      &@     �B@     �p@      ,@     `@      @      @      8@      ,@     �q@      i@      @     �W@     �R@      *@      @      &@     �B@     pp@      ,@     P@      @      @      8@      ,@     �q@     �h@      @     �W@      R@      (@      @      $@      A@     �j@      (@     Py@      �?      @      2@      ,@     �m@      g@      @     @U@       @      �?              �?      @      H@       @      X@      @       @      @             �G@      ,@              "@                                              @              �?                                               @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJP�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?2�
�y�?�	           ��@       	                   �=@�>-�?K            �@                            @L����2�?           ��@                          �4@"<�<3{�?           8�@������������������������       ��C�$��?�           H�@������������������������       �SL���?v           (�@                           @�];j���?           {@������������������������       �Ư�,�?�            �i@������������������������       ��
d� ^�?�            @l@
                            �?�Gw��?-            @R@                            �?�z�G��?             D@������������������������       �d�����?             3@������������������������       �������?             5@                           @��3cڟ�?            �@@������������������������       �n�����?	             .@������������������������       �2�tk~X�?	             2@                           @Cv�l߹�?T           �@                           �?oRe3�v�?            x�@                          �<@0��b�/�?�             n@������������������������       ������I�?�            �k@������������������������       ��&5D�?
             1@                           @�cOM�C�?f           ��@������������������������       ���ww�C�?I           ��@������������������������       ����`5�?             K@                           !@���<�?T           �@                            �?�d��)7�?L           ��@������������������������       �)�mO?��?�            Ps@������������������������       ��vSo�p�?�            �k@������������������������       �      �?             0@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@      =@     �B@      6@     �Z@     ��@     �C@     ��@      4@      @      R@      P@     ��@     �~@      5@     `q@      X@      &@      9@       @     �R@     `t@      4@     �y@      "@      @      A@      C@     �r@     `l@      "@     �b@     @U@      &@      9@       @     @Q@     �s@      4@     �w@       @      @      A@      B@      r@     �k@      "@     `b@     �L@      "@      5@      @      L@     �n@      1@     �o@       @      @      <@      A@     �g@     �d@      "@     @_@     �B@      @      ,@      @     �A@     �[@      "@      _@       @      @      *@      7@      R@      Z@      "@      K@      4@      @      @      @      5@      a@       @      `@      @              .@      &@     �]@      O@             �Q@      <@       @      @      �?      *@      R@      @     @_@                      @       @      Y@     �K@              6@      .@      �?      @      �?       @      A@       @     �F@                      @              M@      @@              $@      *@      �?                      &@      C@      �?      T@                      @       @      E@      7@              (@      &@                              @      @              >@      �?                       @       @      @              @      �?                              @      @              3@                                      @      @              �?                                      @      @              $@                                       @      �?                      �?                              �?       @              "@                                       @      @              �?      $@                              �?       @              &@      �?                       @      @                       @                                      �?                       @      �?                       @      @                              $@                                       @              @                                      �?                       @     @X@      2@      (@      ,@      @@     �t@      3@     H�@      &@      @      C@      :@     �|@     pp@      (@      `@     �S@      ,@       @      &@      8@     �n@      &@     X�@      @       @      9@      3@     �v@     `d@      &@     �W@      .@       @       @      �?      @     �C@      �?     �N@                      @              O@      6@      @      9@      .@       @       @      �?      @      C@      �?     �I@                      @              N@      6@      @      6@                                      �?      �?              $@                                       @                      @      P@      (@      @      $@      4@      j@      $@     �~@      @       @      6@      3@     �r@     �a@       @     �Q@      P@      (@      @      $@      2@     `i@      $@     p}@      @       @      5@      .@     r@     �a@       @     �O@                                       @      @              7@       @              �?      @      "@      �?              @      2@      @      @      @       @     �T@       @     �c@      @      �?      *@      @     @Y@      Y@      �?     �@@      2@      @      @      @       @     @S@       @     �c@      @      �?      *@      @     �X@     �W@      �?      @@      $@       @              @      @     �D@      @     �[@       @               @      @     �I@      F@              6@       @       @      @              @      B@      �?     �G@      @      �?      @      �?     �G@     �I@      �?      $@                                              @              �?                                      @      @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ$FOhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @���c��?�	           ��@       	                   @@@7wPq��?H           �@                           �?x"�˞�?5           ��@                           �?�{�C#d�?�           `�@������������������������       ���U��?�            pq@������������������������       �,[P���?�            Py@                            �?��}����?�           ��@������������������������       ����2�"�?u           �@������������������������       �#Q_���?           �{@
                            @�5��?             ;@������������������������       ���
ц��?	             *@������������������������       �/����?
             ,@                          �;@�����~�?_           �@                           �?9�B���?�           �@                            @܆��C�?�           H�@������������������������       ���eӗ�?|           ��@������������������������       �h���_�?�            `j@                           @U_�N�?�           `�@������������������������       �t.���?�           ��@������������������������       ���ƄIU�?            �E@                            �?�Iwo��?�            0p@                           �?J��J7�?7            @T@������������������������       ����<,�?             9@������������������������       �$I�$I��?)             L@                           @z/sT{�?q            @f@������������������������       �9��8�c�?`             b@������������������������       ���U�(�?             A@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @j@      ?@     �D@      4@     �W@     �@      A@     \�@      ,@      @     �V@      N@     ��@     �@      ;@     �p@     �Z@      3@      9@      *@     �H@     �q@       @     @@      @      @      C@      :@     �t@     @g@      @     �`@     �Z@      3@      9@      *@      G@     �q@       @     ~@       @      @      C@      :@     �t@     @g@      @     �`@      F@      (@      (@      @      ,@     �X@      @     `k@                      2@      (@     �[@     @S@             �L@      *@      @      (@      @      @      E@       @     @U@                      .@      $@      @@     �@@              2@      ?@      @               @      @      L@       @     �`@                      @       @     �S@      F@             �C@      O@      @      *@      @      @@     @g@      @     `p@       @      @      4@      ,@     @k@     @[@      @      S@     �B@      @      @      @      3@     �_@      @     �c@                      $@      @     @^@      H@      @      @@      9@      @      @      @      *@     �M@      �?      Z@       @      @      $@      "@     @X@     �N@       @      F@      �?                              @      �?              3@      �?                               @                              �?                                      �?              "@      �?                              �?                                                              @                      $@                                      �?                             �Y@      (@      0@      @      G@     Pv@      :@     �@      &@      �?     �J@      A@     �x@     0v@      5@     �`@     �V@      (@      0@      @     �E@     Ps@      8@     �@      @      �?     �I@     �@@     �u@     pt@      1@     �^@     �I@      @       @      @      9@      a@      .@     `e@      @      �?      3@      *@     �a@     `b@      *@      L@      E@       @      @      @      4@     @Y@      *@     �\@      @      �?      2@      (@     @X@      [@      *@      F@      "@      @      �?              @      B@       @     �L@                      �?      �?      F@     �C@              (@      D@      @       @      @      2@     �e@      "@     0u@      @              @@      4@     @j@     �f@      @     �P@      C@      @       @      @      1@     �c@      "@     �t@      @              @@      4@     �h@     �e@      @      P@       @                              �?      .@              @                                      (@      @               @      (@                              @      H@       @     @Y@      @               @      �?      E@      <@      @      (@                                      @       @              B@       @              �?      �?      .@      .@              @                                                              *@                                      �?      @              @                                      @       @              7@       @              �?      �?      ,@      "@              �?      (@                                      G@       @     @P@       @              �?              ;@      *@      @      @      (@                                      C@       @     �F@       @              �?              5@      *@      @      @                                               @              4@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ½�ahG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @Px�u�?�	           ��@       	                     �?e�1���?�           ��@                           @x]r����?           ��@                          �?@O�]���?�           x�@������������������������       �|�(�7�?�           ��@������������������������       ����3�E�?             :@                          �0@���]��?�             j@������������������������       ���<,��?             9@������������������������       �zפ����?{            �f@
                           @և��P\�?e            �@                          �1@����v�?�           |�@������������������������       �^�����?�            �t@������������������������       ����b(=�?5           X�@                           �?�H8}9��?h             d@������������������������       �      �?             0@������������������������       ��O�j�?]             b@                           @������?�           (�@                           �?�K4����?=           �@                          �2@��9	C�?�            �t@������������������������       ��lu���?K            @]@������������������������       ��m�ؘ��?�             k@                          �6@���'��?j            �e@������������������������       �� V�?A            �Y@������������������������       �VUUUUU�?)            @Q@                          �?@���ۺ�?|           ��@                           �?k	���?l           ��@������������������������       �o��O>�?�            �k@������������������������       ���q>�?�            �u@������������������������       ��~j�t��?             9@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      =@      D@      >@     �]@     8�@      ;@     �@      (@       @      Q@     �L@      �@     �~@      :@     0q@     �e@      3@      ?@      9@     �X@     �z@      5@     X�@      &@      @      O@      H@     �@     �w@      8@      l@     �K@      @      @      .@      :@     �c@       @     �t@      �?              0@      .@     �i@      ]@       @     �L@      F@      @      @      $@      2@     @`@      @      n@                      &@      $@     @f@     �Y@      @      H@      F@      @      @      $@      2@     @`@      @     @l@                      &@      $@     �e@      X@      @      H@                                                              .@                                      @      @                      &@       @              @       @      :@       @     @V@      �?              @      @      =@      *@      @      "@      �?                              @      �?              @                      @               @      @              @      $@       @              @      @      9@       @     �T@      �?               @      @      ;@      "@      @      @     @]@      *@      8@      $@     @R@      q@      *@     z@      $@      @      G@     �@@     @s@     �p@      0@     �d@     @]@      *@      6@      $@     �P@      p@      $@     pv@      "@      @      D@      ?@     �q@     `n@      0@      c@      =@      @      $@      �?      $@      K@       @      H@      �?       @      ,@       @      G@     �N@      @      A@      V@      $@      (@      "@      L@     @i@       @     ps@       @      @      :@      7@     @m@     �f@      $@     �]@                       @              @      2@      @      M@      �?              @       @      <@      6@              ,@                                              @              @                                      @                                               @              @      (@      @      K@      �?              @       @      6@      6@              ,@      I@      $@      "@      @      4@      g@      @     �y@      �?       @      @      "@     �k@      \@       @     �I@      4@      �?       @      @      $@      M@      �?     �g@               @       @      �?     �\@     �N@              A@      .@      �?      @       @      @      E@      �?      ]@                      �?      �?      R@      G@              :@       @              @       @              $@             �H@                                      B@      $@              @      *@      �?                      @      @@      �?     �P@                      �?      �?      B@      B@              7@      @              @       @      @      0@             �R@               @      �?              E@      .@               @      �?              �?       @      @      ,@             �B@                      �?              ?@      @              @      @               @              �?       @             �B@               @                      &@       @               @      >@      "@      �?      �?      $@     �_@      @     `k@      �?              @       @     �Z@     �I@       @      1@      9@      "@      �?      �?      $@     @^@      @     �j@      �?              @       @     �X@     �I@       @      .@      (@      @                      @     �K@       @      S@                      @      @      ?@      3@       @      @      *@       @      �?      �?      @     �P@      @     `a@      �?                      @      Q@      @@              $@      @                                      @              @                                       @                       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJl��PhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @���D|�?�	           ��@       	                   �<@��)����?�           ��@                            �?�����?H           $�@                           �?�\w����?�           0�@������������������������       �����=�?"           Ћ@������������������������       �n�L����?�           H�@                           �?$=���?           0�@������������������������       �)��<3�?�            �n@������������������������       ��j�=F��?�             u@
                            �?�1ɁA	�?}            �g@                          �@@Nta���?4            �S@������������������������       ��1�^���?-             Q@������������������������       ��G�z��?             $@                          @A@�a*~��?I            @\@������������������������       �g�v��?B            �Y@������������������������       ����k���?             &@                           �?�(���?�           ��@                           �?O��QX�?�           ؄@                           @������?�            Pr@������������������������       �à��i��?�            �m@������������������������       ��:�;73�?            �L@                           @��َ_��?�            `w@������������������������       �g�"8o�?�             l@������������������������       �u�����?Y            �b@                           �?�+�+��?            �}@                           �?贁N��?�             n@������������������������       �{�G�z�?2             T@������������������������       ��Q���?[             d@                           @�U9|H��?�            �m@������������������������       ���.�?p            �f@������������������������       ��0��?#             K@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      D@      B@      5@      X@     �@      >@     ��@      3@       @     @U@     �P@     ��@      �@      3@     0p@     �e@      :@      =@      3@      T@     �|@      7@     h�@      0@      @     �R@     �I@     P|@     �w@      2@     �j@      e@      9@      8@      3@      T@      {@      6@     �@      &@      @     �P@     �I@     pz@     �v@      2@     �g@     �a@      2@      0@      ,@     �J@     pu@      .@     ��@      @             �B@      ?@     �u@     p@      ,@     �`@     �S@      @      .@      @      @@     �c@      "@     �k@      @              4@      4@     �a@     @Z@       @     �Q@      P@      &@      �?      $@      5@     @g@      @     v@                      1@      &@     �i@      c@      @      P@      ;@      @       @      @      ;@     �V@      @     �X@       @      @      >@      4@     �S@     �Z@      @     �L@       @      @      @      @      *@     �B@      @      >@      @      @       @      *@     �@@      J@      @      7@      3@       @      @       @      ,@      K@       @     @Q@       @      @      6@      @      G@      K@      �?      A@      @      �?      @                      9@      �?     �R@      @               @              >@      ,@              5@      �?                                       @             �E@      @                              (@      @              @      �?                                      @              E@      @                              &@       @              @                                               @              �?                                      �?      @               @      @      �?      @                      1@      �?      @@       @               @              2@       @              0@      @      �?      @                      .@      �?      >@       @               @              &@       @              0@                                               @               @                                      @                              H@      ,@      @       @      0@     �f@      @      y@      @      �?      $@      .@      o@     `a@      �?     �G@      A@      @      @      �?      $@      X@      @     �m@      @      �?      @      &@     �_@     �W@      �?      >@      6@      @      @              @     �E@      @     �S@       @      �?      @      @     �N@     �G@      �?      *@      1@      �?      @              @     �E@      @     �H@      �?              @      @     �K@      C@      �?      (@      @       @      �?               @                      =@      �?      �?                      @      "@              �?      (@      �?      �?      �?      @     �J@      @     �c@      �?               @      @     @P@     �G@              1@      "@      �?              �?      @      2@             �[@      �?               @      �?      E@      5@              *@      @              �?                     �A@      @      H@                              @      7@      :@              @      ,@      $@              �?      @     �U@      �?     �d@                      @      @     �^@     �F@              1@      "@       @              �?      @      G@      �?     @R@                      @      @     �H@      :@              0@      "@       @                              $@      �?      2@                       @              5@      $@              @              @              �?      @      B@             �K@                      �?      @      <@      0@              "@      @       @                      �?     �D@              W@                      �?      �?     �R@      3@              �?      @                              �?      :@             �S@                              �?     �L@      0@              �?       @       @                              .@              ,@                      �?              1@      @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�T%FhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @����6��?�	           ��@       	                   �=@sƊP�/�?�           �@                           �?(]o�J�?�           �@                           �?��X����?�           ܒ@������������������������       �ƥ%2�/�?�            �t@������������������������       �5U�~v�?2           p�@                           @�xJ���?�           �@������������������������       �$kLY���?           ��@������������������������       �zoRaj�?            @i@
                           �?~R�q�?_            �`@                           @Z�8��m�?$             I@������������������������       ��0\K5��?            �B@������������������������       �;�;��?
             *@                           @Y�
#)%�?;            �T@������������������������       ����t���?             :@������������������������       ��!��}�?(            �L@                           �?X@Lm�?�           L�@                           �?U}�����?�           (�@                           �?��U�I�?�            �p@������������������������       ����&�?@            @Z@������������������������       ���ݡOH�?m            �c@                           �?�";_��?           �y@������������������������       ���Y�q�?D            �W@������������������������       ���yQ��?�            �s@                           �?������?            �z@                           �?`�pꠝ�?X            @^@������������������������       ��k�n�?9            @U@������������������������       �#e�����?             B@                           @�x�uF�?�            Ps@������������������������       �^s]ev�?H             ]@������������������������       �D�*����?�             h@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @l@      D@     �D@      B@     �Z@     ��@     �C@     ��@      3@      @     �U@     @P@     (�@     @�@      4@     �p@     �e@      ;@      >@     �@@     �T@      |@     �A@     Ѕ@      0@      @      S@     �J@      ~@     �y@      2@     �k@     �e@      8@      >@     �@@     �S@     �z@     �A@     ��@      .@      @     �R@      J@     �|@     �x@      1@      k@      U@      (@      7@      2@     �H@     `h@      5@     @o@      (@      @      B@      9@     �h@     �c@       @     �\@      :@      @      ,@      "@      ,@     �G@      @     �O@      @              2@      @      :@     �D@             �J@      M@      @      "@      "@     �A@     �b@      1@     `g@       @      @      2@      5@     @e@     @]@       @      O@      V@      (@      @      .@      >@      m@      ,@     @x@      @       @      C@      ;@     `p@     �m@      "@     @Y@      T@      (@      @      *@      ;@     �j@      (@     ps@      @       @      =@      6@     �l@      k@      @     �U@       @              �?       @      @      5@       @     @S@                      "@      @      A@      5@      @      .@      �?      @                      @      4@              N@      �?               @      �?      6@      ,@      �?      @      �?                              @      @              <@                                      @      "@               @      �?                              @      @              7@                                      @      @                                                                              @                                              @               @              @                              0@              @@      �?               @      �?      3@      @      �?      @              @                              @              @      �?               @              @      �?      �?       @                                              &@              <@                              �?      (@      @              �?     �J@      *@      &@      @      8@     �f@      @     `w@      @              &@      (@     �l@     �a@       @     �E@      E@      @      $@      @      0@     �X@       @     �m@      �?              @      &@     �[@     @Y@       @     �@@      <@      @      @              $@      F@       @      P@                      @      @     �B@      H@      �?      (@      @               @              @      :@              <@                       @       @      ,@      2@              @      7@      @      @              @      2@       @      B@                       @      �?      7@      >@      �?      @      ,@              @      @      @     �K@             �e@      �?              �?       @     �R@     �J@      �?      5@      @              @              @      $@             �@@                                      7@      *@              @      &@                      @      �?     �F@             �a@      �?              �?       @     �I@      D@      �?      0@      &@      "@      �?               @     �T@       @      a@       @              @      �?     �]@      E@              $@      "@      @                       @      0@             �@@                      @             �A@      .@              @      @      @                       @      *@              .@                      @              9@      (@              @       @                                      @              2@                                      $@      @                       @      @      �?              @     �P@       @      Z@       @               @      �?     �T@      ;@              @       @      @      �?              �?      9@       @      >@                              �?     �C@      $@               @              @                      @      E@             �R@       @               @              F@      1@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�X^hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @���N�_�?�	           ��@       	                     �?yd�0��?�           �@                           �?�C��G��?�           ��@                           �?�:�ߤ�?           �{@������������������������       ��A����?t             g@������������������������       ��j(�?�            0p@                           @�ވF?�?�           ��@������������������������       �0Σ��)�?�           �@������������������������       ��X�%��?
             .@
                           @��[�4�?[           \�@                           �?�3��7H�?�            �@������������������������       �iv��=�?�            �g@������������������������       �����9�?u           �@                          �;@:w5g��?e            �b@������������������������       �paRC4%�?[             a@������������������������       ����Q��?
             .@                           �?h�����?�           �@                          �2@����?�           ؄@                           �?�1X4Y��?[            �c@������������������������       �!{�/���?'             Q@������������������������       �ޏ��k��?4             V@                           @����&�?B           �@������������������������       �֤E�?�            �l@������������������������       ��v���o�?�            �q@                           @� `��?           �z@                           @�n? ���?�            �p@������������������������       �Ҹ�蘗�?|             h@������������������������       �}��\��?2            �R@                          �5@~��ơ�?k            �c@������������������������       ������?;            @U@������������������������       �HR�F��?0            �R@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      <@     �F@      9@      W@     ��@     �C@     ��@      $@      @      Q@      I@     ��@     ��@      1@     pp@     `b@      8@      >@      4@     @S@     P~@     �A@      �@      @      @      M@      F@     �@     �x@      ,@     �k@      L@      &@      (@      @      4@     `f@      0@     �t@      @              *@      $@     �k@      a@      @      F@      6@      @      "@       @      ,@      R@      @     @^@      �?              @       @      W@     �I@      @      @@      @       @      "@      �?      @      7@      @      K@                      @      @      =@      2@       @      7@      0@      �?              �?      &@     �H@      @     �P@      �?              �?      @     �O@     �@@      �?      "@      A@       @      @      @      @     �Z@      $@     �j@       @              @       @     @`@     �U@       @      (@      @@      @      @      @      @     @Y@      $@     `j@       @              @       @      `@     @U@       @      (@       @      �?                      �?      @               @                                       @      �?                     �V@      *@      2@      *@     �L@      s@      3@     `y@      @      @     �F@      A@     @r@     Pp@      "@     @f@      V@      *@      1@      *@      K@     �q@      ,@     v@      @      @     �D@      >@     q@     @m@      "@     �d@      $@               @      @      &@      ?@              =@      �?               @      @     �G@      7@       @      5@     �S@      *@      .@      "@     �E@     �o@      ,@     @t@      @      @     �C@      9@     @l@     `j@      @      b@      @              �?              @      4@      @     �J@                      @      @      3@      ;@              (@      @              �?              @      3@      @     �E@                      @      @      .@      ;@              (@                                              �?              $@                                      @                              E@      @      .@      @      .@     @f@      @      x@      @       @      $@      @     `n@      a@      @     �D@      =@      @      ,@       @       @      [@      �?      o@      �?       @      @       @     �\@     �V@      @     �A@      @               @      �?      @      8@              C@                      @              =@      :@              1@                      @              @      0@              ,@                      @               @      "@              $@      @              @      �?      �?       @              8@                                      5@      1@              @      8@      @      @      �?      @      U@      �?     `j@      �?       @       @       @     �U@      P@      @      2@       @              @      �?       @      9@             �Z@              �?       @      �?     �C@      4@              1@      0@      @                      �?     �M@      �?     @Z@      �?      �?              �?     �G@      F@      @      �?      *@      �?      �?      @      @     �Q@      @      a@       @              @      @      `@      G@              @      "@              �?      @      @      >@      �?     �T@                      @      �?     �X@      ;@              @      @              �?              @      0@      �?     �P@                      @             @S@      ,@              @      @                      @      �?      ,@              0@                       @      �?      5@      *@                      @      �?                      �?      D@       @      K@       @                      @      >@      3@              @      @      �?                      �?      &@      �?      @@                              @      0@      *@              @                                              =@      �?      6@       @                              ,@      @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJoN+hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@"`����?�	           ��@       	                     @K�e!"��?�           @�@                          �5@tB�1��?.           ��@                            �?m�����?�           @�@������������������������       �l����?�           �@������������������������       �+_��'��?           �x@                            �?@�n?���?Q           x�@������������������������       �s�"#k��?�           ��@������������������������       �v&�[r�?�            �o@
                           �?;y#��z�?j           �@                          �2@/
kg�?            {@������������������������       ��=�9�?W             a@������������������������       �!�;M��?�            pr@                           @6OD1��?P           ��@������������������������       ��iA��?           �y@������������������������       ��2�
��?J             ]@                           @5�e����?           �z@                          @A@f3�����?�            �r@                           @WH�,�?�            pq@������������������������       ��]u�X��?�            �k@������������������������       ��)x9/�?'             L@������������������������       ��z�G��?             4@                          �@@ll@�?O            �_@                            �?��	���?D            @[@������������������������       �g\�5�?             :@������������������������       ��G?`��?4            �T@������������������������       ��F����?             1@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@     �@@     �A@      @@     @V@     ��@      B@     (�@      *@      @      T@     �Q@     ��@      �@      4@     �p@     �g@      =@     �@@      @@      U@     p�@      A@     0�@      $@      @     @R@     @P@     (�@     �@      .@     @m@      d@      1@      4@      <@      P@     �y@      >@     �@      "@      @     �M@      L@     �}@     �w@      ,@      g@      [@      &@      (@      ,@      E@     �n@      4@     0y@      @             �B@      C@     �p@     �k@      &@     �]@     @R@      @      "@      &@      @@     `g@      .@     u@      @              .@      2@     �j@     `b@      @      T@     �A@      @      @      @      $@      N@      @     �P@                      6@      4@      K@     @R@      @      C@     �J@      @       @      ,@      6@     �d@      $@      j@      @      @      6@      2@     `j@      d@      @     �P@      A@      @      @      &@      &@      a@      "@     `d@       @              0@      *@     �c@      [@      @      H@      3@       @      @      @      &@      <@      �?     �F@       @      @      @      @      J@      J@              3@      >@      (@      *@      @      4@     @b@      @     0t@      �?              ,@      "@      i@     �`@      �?     �H@      1@      @       @       @      *@      S@      @     �]@                      &@      @     @V@     �M@              8@       @              @       @      @      4@      �?      J@                      @       @      8@      &@              $@      .@      @      @              "@      L@       @     �P@                      @       @     @P@      H@              ,@      *@      @      @       @      @     �Q@      �?     �i@      �?              @      @     �[@      S@      �?      9@      "@      �?      @       @      @     �G@      �?     @f@      �?              @      @      U@      J@              5@      @      @                      �?      7@              :@                               @      ;@      8@      �?      @      0@      @       @              @     �Q@       @     �d@      @      �?      @      @      S@     �@@      @      ?@      *@      @       @              @     �G@       @     �X@       @      �?      @      @     @P@      1@      @      <@      *@      @       @              @      G@       @     @V@       @      �?      @      @      L@      1@      @      ;@      $@      @      �?              @      A@       @      S@      �?      �?      @       @      C@      0@      @      8@      @              �?              �?      (@              *@      �?                      @      2@      �?              @                                              �?              "@                                      "@                      �?      @                                      8@             �P@      �?               @              &@      0@              @       @                                      5@              O@      �?               @              $@       @              @                                                              5@                      �?              @                      �?       @                                      5@             �D@      �?              �?              @       @               @      �?                                      @              @                                      �?       @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJC�\hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @��w��?�	           ��@       	                     �?�����?�           �@                           @.��?N           ��@                          �?@&�:Ƃ��?           Й@������������������������       �(�u���?�           D�@������������������������       �|L�Sw�?            �A@                           @�p�9�i�?@           �~@������������������������       �p�%ΦD�?o            �d@������������������������       ���#���?�            @t@
                           �?pN�����?�           �@                          �6@4� Uz�?�            �m@������������������������       ��g���%�?q             f@������������������������       ��!-�5p�?"            �N@                           @��/�ژ�?           `{@������������������������       ������?�            �n@������������������������       ��$}_��?w             h@                           �?u�9@4�?�           �@                           @b֍g��?o            @g@                           @����P?�?Y            @b@������������������������       �l�(�|�?K            �^@������������������������       ��q�q�?             8@                           �?��Q���?             D@������������������������       �؂-؂-�?             .@������������������������       ��������?             9@                           �?�)[���?R           h�@                           �?�XO5�?&           �|@������������������������       ���;{���?i            @e@������������������������       �x�mQ��?�            @r@                          �2@�JK�5�?,           �{@������������������������       �߉[po�?a            �a@������������������������       ��ԍx&�?�             s@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@     �A@     �B@      7@     @^@     ��@      =@     l�@      2@       @      W@     @P@     0�@     �@      :@     �p@     �a@      8@      9@      2@     �W@     �|@      9@     ؆@      ,@      @      T@      L@     p}@     `z@      :@      l@      [@      0@      4@      .@      K@     �v@      2@     (�@      &@       @      J@     �@@     �w@      r@      .@     �b@     �W@      $@      *@      ,@      A@     �p@      *@     �|@       @              F@      9@     �s@     �m@       @      Z@     �W@      $@      *@      ,@      A@     �p@      *@     0{@       @              F@      9@     �s@     `m@       @     �Y@                                              @              9@                                      �?      @              �?      *@      @      @      �?      4@     �V@      @      c@      @       @       @       @      Q@      J@      @     �G@      �?      @      @              @      3@             @P@      @               @      �?      8@      1@      @      2@      (@       @      @      �?      ,@      R@      @      V@               @      @      @      F@     �A@      @      =@     �@@       @      @      @      D@     �X@      @     �]@      @      @      <@      7@      V@     �`@      &@     @R@      ,@      @       @       @      3@     �A@      �?      8@      �?              @      (@     �B@      G@      @      =@      $@      @       @              1@      ?@              2@      �?              @      (@      =@      6@      �?      7@      @      �?               @       @      @      �?      @                                       @      8@      @      @      3@      @      @      �?      5@      P@      @     �W@       @      @      6@      &@     �I@     �U@      @      F@      &@       @      @      �?      $@      E@      @     �E@       @       @      @      @      C@      F@      @      =@       @      �?                      &@      6@      @     �I@               @      .@       @      *@      E@       @      .@     �H@      &@      (@      @      ;@     `e@      @      x@      @       @      (@      "@     �m@      _@              E@      &@              @              @      9@       @     �G@                      @             �D@      =@              (@      @              @              �?      2@       @      D@                      @             �B@      0@              (@      @              @              �?      1@              ;@                      @             �@@      .@              &@       @                                      �?       @      *@                                      @      �?              �?      @                              @      @              @                                      @      *@                                                      �?      @              @                                       @      @                      @                              @      @              @                                       @       @                      C@      &@      @      @      5@     @b@       @     u@      @       @      @      "@     �h@     �W@              >@      8@      @      @       @       @     �Q@       @     �g@       @       @              @      V@      H@              .@      2@      @      @              @      3@      �?     �P@              �?              �?      ;@      3@              @      @      �?               @       @     �I@      �?     �^@       @      �?               @     �N@      =@              &@      ,@      @      @      @      *@      S@             `b@       @              @      @     �[@     �G@              .@      "@                      @      �?      1@             �D@                      @       @     �I@      (@              @      @      @      @              (@     �M@             �Z@       @               @      @     �M@     �A@              &@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�>hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx                             �?T%�i��?�	           ��@       	                     �?Ô�6�?S           �@                           �?$7���N�?           @{@                          �:@Du�W��?l            �d@������������������������       �VQ&�N�?W            �`@������������������������       �     `�?             @@                           �?P�n#X�?�             q@������������������������       ���
O�?G            @\@������������������������       ������?^            �c@
                          �;@���J�?B           4�@                            @B8�h�\�?�           �@������������������������       ������?�           �@������������������������       ��5�&	�?           �z@                           @{������?S            �`@������������������������       �V4�ͫ�?M             ^@������������������������       �d}h���?             ,@                           !@`_J�)��?n           �@                          �;@�[�-��?c           �@                            @����?�           ��@������������������������       ��R���?]           �@������������������������       ��ȯ	�~�?b           ��@                           �?9��i3�?�             o@������������������������       �Y7Ҍ�A�?#            �K@������������������������       ����xr��?�             h@������������������������       ��8��8��?             8@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@      6@      C@      7@      ]@      �@      B@     d�@      5@      (@     �R@     �L@     �@      �@      3@      o@     @Y@      0@      :@      $@     �N@     �r@      8@     �z@      ,@       @      A@      ?@     �r@     �n@      "@      ^@      4@      @       @      @      1@     �N@       @     @a@       @              @      $@     �R@     �N@       @      <@       @      @       @       @      @      0@      @      N@                       @       @      <@      ,@       @      1@       @      @       @       @      �?      *@       @      E@                       @       @      ;@      ,@       @      (@                                       @      @      @      2@                                      �?                      @      (@      �?              �?      ,@     �F@      @     �S@       @              @       @     �G@     �G@              &@      @                      �?      @      :@      @      ?@                               @      3@      &@               @      @      �?                      "@      3@             �G@       @              @      @      <@      B@              @     @T@      (@      8@      @      F@     �m@      0@      r@      (@       @      =@      5@     �l@      g@      @      W@     �Q@      "@      7@      @      E@     �k@      0@     �n@      "@       @      <@      5@      j@     �d@      @     �T@     �H@      @      1@      @      @@     �a@      (@     �_@      "@      @      7@      2@     �\@     �Y@      @     @P@      6@      @      @              $@     �S@      @     �]@               @      @      @     �W@      O@              1@      $@      @      �?               @      0@              G@      @              �?              4@      4@       @      $@      $@      @      �?               @      0@             �A@      @              �?              1@      4@       @      $@                                                              &@                                      @                             �[@      @      (@      *@     �K@     `w@      (@     h�@      @      @      D@      :@     �z@     �p@      $@      `@     �[@      @      (@      *@     �K@     �v@      (@     @�@      @      @      D@      :@     �z@     �p@      $@      `@     @Y@      @      (@      &@      J@     �s@      &@     �@      @      @     �B@      9@     �w@     `n@      "@     @^@      U@       @      "@      @      G@     @m@      $@      w@       @      @     �A@      0@     �n@     �f@       @      X@      1@       @      @      @      @      U@      �?     `j@       @               @      "@      a@     �N@      �?      9@      $@       @               @      @      F@      �?     @Y@      @      �?      @      �?     �G@      5@      �?       @      @       @                      @      $@              &@                                      .@       @               @      @                       @              A@      �?     �V@      @      �?      @      �?      @@      *@      �?      @                                              (@              @                                      �?      @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJC=9qhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�
��s�?�	           ��@       	                   �=@��]%�?G           ��@                          �7@�5�4B �?           ,�@                           @��,�L�?            �@������������������������       ��7��>�?�           0�@������������������������       �@���4�?{            �f@                          �:@-��S�?            �x@������������������������       �ҌJW�?�            p@������������������������       �n��E�?[            @a@
                            @6Ql����?3            @U@                           @�>4և��?!             L@������������������������       �F]t�E�?             F@������������������������       �9��8���?             (@                          �>@>���Rp�?             =@������������������������       �b���i��?             &@������������������������       ���Hx��?             2@                          �7@�P���?�           R�@                            @+?���0�?�           ��@                           @B�����?�           ��@������������������������       ��@�t��?c            �@������������������������       �n,�Ra�?n             f@                          �2@D��{�?           �x@������������������������       �,V�����?i            @e@������������������������       �}ݕ2޼�?�            �l@                          �;@��V��?�           X�@                          �8@V��b&��?
           �z@������������������������       �R5��\�?S            @`@������������������������       ���X��7�?�            pr@                           @n=g����?�             p@������������������������       �(��/n��?�            �k@������������������������       ��Xp��?             C@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        k@      ;@      D@      =@      X@     ��@      7@     ��@      ,@      @     @T@      Q@     x�@     ��@      .@     `o@     @W@      4@      =@      *@      I@     �s@      (@     �x@      "@      @     �A@     �A@     �s@     @n@      @     �_@     @U@      4@      =@      *@     �F@     @s@      (@     �v@       @      @     �A@     �A@      r@     �l@      @      _@      O@      1@      8@      "@      D@      j@      &@     �q@       @      @      =@      @@     �i@     �f@      @      W@      H@      1@      4@      @      :@     �e@      "@     �m@       @      @      :@      >@     �g@     �c@      @     �S@      ,@              @      @      ,@      B@       @     �F@                      @       @      1@      9@              *@      7@      @      @      @      @      Y@      �?     �T@                      @      @     �T@     �G@              @@      0@                      @      @     �R@             �E@                      �?      @      J@     �C@              6@      @      @      @      �?      �?      :@      �?      D@                      @              ?@       @              $@       @                              @      @              >@      �?                              6@      (@      �?       @      @                              @       @              7@                                      $@      (@               @       @                              @       @              4@                                       @      @               @      �?                                                      @                                       @      @                      @                              �?       @              @      �?                              (@              �?              @                              �?      �?              �?                                      @                              �?                                      �?              @      �?                               @              �?              _@      @      &@      0@      G@     `t@      &@     Ȇ@      @      @      G@     �@@     p{@      r@       @     @_@     �W@      @      $@      "@      ;@     �l@      @     @}@      @       @      @@      <@      r@     @l@      @     �X@     �Q@      @      @      @      7@     �f@      @     Ps@       @       @      ?@      5@     �i@     `g@      @     �S@     @Q@      @      @      @      4@     �b@      @     �n@       @       @      6@      1@     �e@     �d@      @     �Q@      �?      �?                      @      @@      �?      O@                      "@      @      >@      5@      @      "@      9@              @      @      @     �G@      �?     �c@      �?              �?      @      U@     �C@              4@      ,@              @      @      @      (@             �M@                               @     �F@      3@              "@      &@               @      �?      �?     �A@      �?      Y@      �?              �?      @     �C@      4@              &@      =@       @      �?      @      3@     @X@      @     Pp@       @      �?      ,@      @     �b@      O@       @      :@      6@       @      �?      @      0@      H@      @      c@              �?       @       @      Z@     �G@              ,@      @              �?              @      3@      �?      O@                      @      �?      2@      &@               @      1@       @              @      *@      =@       @     �V@              �?      �?      �?     �U@      B@              (@      @                      @      @     �H@      �?      [@       @              @      @     �G@      .@       @      (@      @                      @      @      F@      �?     @T@       @              @      �?      F@      .@       @      (@                                              @              ;@                      �?       @      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�e�phG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �0@! �!d�?�	           ��@       	                    @ƈ��4g�?�            �i@                           �?� ����?X            �^@                           @��6�/�?)             O@������������������������       ��q�q��?              H@������������������������       ����>4��?	             ,@                           @��\�U �?/            �N@������������������������       �vb'vb'�?'             J@������������������������       �VUUUUU�?             "@
                           @eģ���?6            �T@������������������������       �     ��?             0@                           @f������?+            �P@������������������������       �@˜��H�?             G@������������������������       ���&%���?             5@                            @�2�J�?"	           ��@                           @�_<V���?o           `�@                            �?'2,��?�           @�@������������������������       ��eM�gN�?>           x�@������������������������       �PC)j��?�            p@                            �?3��'$��?�           ��@������������������������       �Ԓ6�Um�?�           �@������������������������       ���A�t��?�            @v@                           �?�Œ����?�           ,�@                           @Z�1NU��?A           �@������������������������       �Ah���?           P{@������������������������       �H�ϵ�?&            �Q@                          �;@�MwR���?r           ��@������������������������       �n8�ށ��?F           8�@������������������������       �������?,            @R@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        g@      C@      C@      4@     @Z@     ��@      <@     `�@      "@      @     �T@     @P@      �@     �~@      ,@      o@      "@                              "@      B@      "@      C@       @      �?      @      @      =@      F@      �?      0@      @                              @      6@      @      ,@                      @      @      6@      7@      �?      *@      @                              @      @      @      @                      @      �?      &@      $@      �?      "@       @                              @      @      @      @                      @      �?      "@      $@      �?      @       @                               @                      �?                      �?               @                      @       @                                      0@              $@                      �?      @      &@      *@              @       @                                      (@              @                              @      &@      (@              @                                              @              @                      �?                      �?                      @                              @      ,@      @      8@       @      �?      �?              @      5@              @       @                              �?      �?              "@                                       @      �?                      �?                               @      *@      @      .@       @      �?      �?              @      4@              @                                       @      &@      @      *@       @      �?      �?              @      @               @      �?                                       @      �?       @                                      �?      *@              �?     �e@      C@      C@      4@      X@     ��@      3@     Ȑ@      @      @      S@      N@     �@     0|@      *@      m@      a@      <@      :@      2@      T@      }@      0@     (�@      @      @     �P@      K@     P@     �t@      (@      h@      S@      *@      $@      $@     �B@     `k@       @     `s@      �?       @      2@      :@     �l@     @[@      @      Y@      K@       @      $@       @      7@      f@       @     �p@      �?              1@      .@     �e@     �T@      @     �Q@      6@      @               @      ,@     �E@             �F@               @      �?      &@     �J@      ;@       @      >@      N@      .@      0@       @     �E@     �n@      ,@     �v@      @       @      H@      <@     q@     �k@      @     @W@     �E@      &@      "@       @      =@     �h@      (@     �q@      �?              :@      ,@     �k@      e@      @     �L@      1@      @      @              ,@     �H@       @      T@       @       @      6@      ,@     �J@      J@       @      B@     �C@      $@      (@       @      0@      i@      @     �x@      @              $@      @     �m@     �^@      �?      D@      ;@      $@      $@              "@     �[@       @     `c@      @              @      �?      W@     �L@              7@      ;@      @       @              @      W@       @     �a@      @               @      �?      T@     �H@              2@              @       @              @      3@              *@                      @              (@       @              @      (@               @       @      @     @V@      �?     @n@                      @      @     @b@     @P@      �?      1@      &@               @       @      @     �Q@      �?     �i@                      @      @      a@      O@      �?      .@      �?                              �?      3@             �B@                                      $@      @               @�t�bub�     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�8�'hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?sk����?�	           ��@       	                     @�ΩI�?�           ��@                            �?��&:��?M           ��@                           @�v4��?           �|@������������������������       �'c�E!�?�            �u@������������������������       ���_'y�?J            �[@                           @�x�9!��?1           `~@������������������������       ���z·�?�            v@������������������������       �Ƃ�DL��?W            �`@
                          �0@��BX��?�           ��@������������������������       �����H�?
             2@                           @����5��?�           `�@������������������������       �k�a��?�            �r@������������������������       �:��$^�?�            0t@                           �?~�f���?�           6�@                            @o���9�?�           t�@                          �>@pRT�U�?T           �@������������������������       �7DmS�?F           �@������������������������       �s
^N���?             <@                          �;@�Cc}h��?�             l@������������������������       �� �f���?�            �i@������������������������       �VUUUUU�?             2@                          �0@�8_���?�           ��@                           @���	߬�?.            @Q@������������������������       �     ��?             @@������������������������       ����{z�?            �B@                           @V~��&��?�           �@������������������������       �y1�K��?�            �q@������������������������       �s��O��?�           ��@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `l@      A@     �C@      5@     @Y@     `�@      A@     d�@      7@      @     �U@     �Q@     ��@     �@      4@     @p@     �U@      ,@      5@      @      F@      l@       @     p@      $@      �?      A@      9@     pq@     �h@      $@      ]@     �M@      *@      ,@      @      <@      a@      @     0p@      @              :@      .@     �c@     @_@      @     �V@      <@       @       @      @      *@     �P@      @     @c@      �?              ,@       @     �S@     �G@             �B@      9@                      �?      $@     �K@       @     �[@                      &@      @     @P@      ?@              ?@      @       @       @      @      @      &@      �?     �E@      �?              @      @      ,@      0@              @      ?@      &@      (@      �?      .@     �Q@      �?     @Z@      @              (@      @     �S@     �S@      @     �J@      6@      &@      &@              ,@      B@             �P@      @              $@      @     @P@     �O@      @      D@      "@              �?      �?      �?     �A@      �?      C@       @               @              *@      .@       @      *@      <@      �?      @      �?      0@      V@      @     �n@      @      �?       @      $@     �^@     �R@      @      :@                                       @      �?              @                              �?      @      @                      <@      �?      @      �?      ,@     �U@      @      n@      @      �?       @      "@     �]@     �P@      @      :@      "@              @      �?       @     �A@       @      `@      �?              @      @      I@      ?@              2@      3@      �?      @              @      J@       @     �[@      @      �?       @      @     @Q@      B@      @       @     �a@      4@      2@      .@     �L@     �x@      :@     �@      *@      @     �J@      G@     �}@     s@      $@      b@      W@      "@       @       @      D@     �i@      .@     �o@      @       @      7@      :@     �l@     �d@      @     @V@     �T@       @       @      @     �A@     @e@      &@     �h@      @       @      .@      6@     `f@     �a@      @     @Q@     �S@       @       @      @     �@@     @e@      &@     �g@      @       @      .@      6@     `f@     �_@      @     �P@      @                               @                       @                                              *@               @      $@      �?              �?      @      B@      @     �L@                       @      @      J@      :@              4@      $@      �?              �?      @      B@      @      K@                       @      @     �E@      9@              0@                                      �?                      @                                      "@      �?              @      H@      &@      $@      @      1@     �g@      &@     0v@       @      �?      >@      4@     �n@     `a@      @     �K@                              �?              *@              *@                              @      (@      4@              @                                              @              @                              @      @      ,@               @                              �?              $@              "@                                      @      @              @      H@      &@      $@      @      1@      f@      &@     `u@       @      �?      >@      1@      m@     �]@      @      H@      1@      @      @       @      �?      D@      @     �T@                      @      �?     �V@      :@              @      ?@       @      @      @      0@      a@      @     0p@       @      �?      :@      0@     �a@     @W@      @      E@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJϩ�~hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @c[�[ ��?�	           ��@       	                    �?����a�?           �@                           @/���y��?)           ��@                           �?i�NI��?�           @�@������������������������       �+sI�v�?X            �`@������������������������       ���6�n�?�           $�@                           �?F3Ԟ(��?=            �U@������������������������       ��X�C�?
             ,@������������������������       ��� �3�?3            @R@
                            �?���݅�?�           |�@                           @�rC�?�           |�@������������������������       ���{�6M�?F           �@������������������������       ���ы*��?�           �@                          �4@��8���?�             x@������������������������       �__+F��?v            �f@������������������������       �ie�^�6�?y            @i@                           �?�c���?�           �@                           @T�8�~�??            @                           @"�X���?            {@������������������������       ��q�`B�?�            �v@������������������������       ��yB����?%            �Q@                           @     ��?-             P@������������������������       �IPolg��?"            �H@������������������������       �
ףp=
�?             .@                          @@@>"��?q           ��@                           @�c�^s��?c           Ё@������������������������       �)Ң���?I           x�@������������������������       ��iQT�?            �E@                          �@@�Ҍ���?             7@������������������������       �<+	���?             .@������������������������       �      �?              @�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      F@      B@      ?@     @X@     P�@      ?@     �@      0@      &@     �U@     �N@     8�@      @      2@     �p@     �d@      ?@      =@      8@     �S@     P}@      6@     @�@      (@       @     �R@      H@     @�@      x@      2@     �k@      T@      ,@      8@      $@     �I@      k@      "@      q@      $@      @      A@      6@     �j@     �e@      (@     �[@     �S@      ,@      6@      $@      E@     �i@       @     @o@       @      @      A@      5@      i@      d@      (@     @X@      @       @      @      �?      @      .@       @      B@       @              "@              2@      &@              4@     �Q@      (@      1@      "@     �A@      h@      @     �j@      @      @      9@      5@     �f@     �b@      (@     @S@       @               @              "@      "@      �?      8@       @                      �?      (@      &@              ,@                                               @              @                                      @                               @               @              "@      @      �?      1@       @                      �?      @      &@              ,@     �U@      1@      @      ,@      <@     �o@      *@     `{@       @      @     �D@      :@     @s@     �j@      @     �[@     �O@      0@      @      (@      *@     �i@      &@     0v@       @              0@      ,@     �n@     `c@      @     �Q@     �E@      @      �?       @      @     �X@      @      b@       @              @      @     �^@     �L@             �B@      4@      $@       @      @      @     �Z@      @     `j@                      (@      @     �^@     �X@      @     �@@      8@      �?       @       @      .@     �G@       @     �T@              @      9@      (@      P@     �M@      @     �D@      $@              �?       @       @      4@       @      C@                      &@      @      2@      A@      �?      >@      ,@      �?      �?              @      ;@             �F@              @      ,@      @      G@      9@       @      &@     �C@      *@      @      @      2@     �f@      "@     �w@      @      @      (@      *@     �o@     �[@              E@      :@       @      @       @      "@     @W@      @      b@              �?      $@      @     �[@      J@              9@      9@      @      @              @     �R@      @     @`@              �?      @      @     �Y@      E@              8@      9@      @      @              @     @Q@      @     @Y@              �?       @      @      S@      D@              7@                                      �?      @              =@                      @              ;@       @              �?      �?       @      @       @       @      2@      �?      ,@                      @              @      $@              �?      �?              @       @       @      0@              @                       @              @      $@              �?               @                               @      �?      @                      �?               @                              *@      @      �?      @      "@      V@       @     @m@      @       @       @       @      b@      M@              1@      *@      @      �?      @       @     �U@       @      l@      @               @       @     �a@      M@              1@      *@      @      �?      @       @     �R@       @      k@      @               @       @     @_@      J@              1@              �?                              (@               @                                      0@      @                                                      @      �?              "@               @                      @                                                              @      �?              @               @                      �?                                                                                      @                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?Yj��ߔ�?�	           ��@       	                   �;@N0��$�?A           ؚ@                          �1@Ur�s/�?�           ��@                           @�m�S���?�            �r@������������������������       ���t���?�             r@������������������������       ��]�`��?	             *@                           �?��3d��?           ܒ@������������������������       ��-t��?q            �e@������������������������       �p����?�           $�@
                           @IPS!�0�?{             j@                            �?�T�}���?a            �d@������������������������       ���FP=c�?            �F@������������������������       �ƒ_,���?F             ^@                          �=@h�1aR�?            �E@������������������������       �m��1G��?             :@������������������������       �@�0�!��?
             1@                            @����?u           &�@                            �?��*���?�           ��@                           !@46�E��?�           ܒ@������������������������       ����%��?�           ��@������������������������       �B{	�%��?             "@                           �?ƛ+�4��?�            �x@������������������������       �      �?             @@������������������������       ��<n�Ь�?�            �v@                          �=@���.]g�?z           ��@                           @N� ��j�?Y           �@������������������������       ��++KE��?�            @n@������������������������       ����`ͺ�?�            s@                           @HXD���?!            �H@������������������������       ��d��0�?             >@������������������������       �$����%�?
             3@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        l@      :@     �E@      6@     @]@     @�@      >@     �@      3@      @     �R@      K@     @�@      �@      7@     �n@     �\@      .@      =@      .@     �Q@     �s@      5@     �y@      "@      @     �@@      9@     s@     `k@       @     @^@      V@      &@      8@      .@      O@     r@      5@     �u@      "@      @      @@      9@     0q@     �h@      @     @Z@      0@       @      @       @      6@      M@      "@      I@       @      �?      "@       @     �G@     �B@      @      @@      0@       @      @       @      4@     �L@      "@      I@       @      �?      "@       @     �G@      @@      @      <@                      �?               @      �?                                                              @              @      R@      "@      3@      *@      D@     �l@      (@     �r@      @      @      7@      1@     �l@     �c@      @     @R@      $@      �?      @      �?      @      6@              M@      �?              @      �?      @@      4@              .@      O@       @      .@      (@      B@      j@      (@     �m@      @      @      2@      0@     �h@     `a@      @      M@      :@      @      @               @      9@             @Q@                      �?              >@      7@      �?      0@      :@      @      @               @      2@              H@                      �?              9@      0@      �?      *@                                      @      (@              2@                                      @                      @      :@      @      @              @      @              >@                      �?              3@      0@      �?       @                                              @              5@                                      @      @              @                                              @              &@                                      @      @               @                                                              $@                                       @      @              �?     �[@      &@      ,@      @     �G@     �v@      "@     �@      $@       @     �D@      =@     py@     �t@      .@     �^@     �W@      &@       @      @     �D@     �p@      "@     |@      @       @     �A@      9@     @q@     �o@      (@      Z@     �Q@      $@      @      @      3@      j@       @     �w@      @              1@      ,@      k@     �e@      @     @Q@     �Q@      $@      @      @      3@     @i@       @     �w@      @              1@      ,@      k@     �e@      @     @Q@                                              @              �?                                      �?                              9@      �?      @       @      6@     �L@      �?     �Q@      �?       @      2@      &@     �M@     �S@      @     �A@       @              �?               @      @              @                      �?              *@      @      �?      �?      7@      �?      @       @      4@      K@      �?      Q@      �?       @      1@      &@      G@     @R@      @      A@      0@              @      �?      @      Y@              l@      @              @      @     ``@      S@      @      3@      .@              @      �?      @      V@              j@      @              @      @     �\@      S@      @      3@      @              @      �?      �?      8@             �Y@                      @      �?     �M@      ;@              &@       @               @               @      P@             �Z@      @              �?      @     �K@     �H@      @       @      �?                              @      (@              0@                                      1@                              �?                              @       @              *@                                      &@                                                                      $@              @                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ(]A*hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�{�y�?�	           ��@       	                    �?Xz���?�           t�@                          �=@Uz�k��?           ��@                           �?>����?�           D�@������������������������       ��7=�A�?�            �q@������������������������       ����q[�?6           ��@                           @��ۚ�R�?             G@������������������������       �L�p.0�?             5@������������������������       ��N@a��?             9@
                          �0@v/$��e�?�           �@                           �?` ���t�?5            @Y@������������������������       ��8��8��?             (@������������������������       �#���?.            @V@                            �?�e���@�?�           X�@������������������������       �ȞMT%�?e           ��@������������������������       �!�Y�h��?,           �@                           �?�͠�6�?�           <�@                          �6@�Q�����?t            �g@                           @:m���?I             ^@������������������������       ��(\����?)            �Q@������������������������       ��(��0�?              I@                           @�a2o��?+            @Q@������������������������       �������?              I@������������������������       ��$�_�?             3@                          �<@&�ҷ�?U           ��@                           �?��y��?           Њ@������������������������       �=[6` �?�            �w@������������������������       �:�/���?           �}@                           �?|�j�Y��?I             ^@������������������������       ��q�q��?             H@������������������������       ��n���?.             R@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@     �@@      C@      =@     @[@     Ѓ@     �A@     ��@      <@      "@     �Q@     �N@     H�@     �}@      2@     �p@     �d@      =@      <@      5@     �U@     �z@      :@     �@      4@      @     �O@     �J@     �~@      v@      .@     `l@      Q@      ,@      5@      "@     �M@     �h@      (@     �p@      $@      @      <@      A@      k@     @d@       @      Z@     �P@      ,@      5@      "@     �K@     �h@      (@     �n@      $@      @      <@      A@     �j@      c@       @     �Y@      &@      @      ,@       @      @     �F@       @     �M@      @              0@      @     �A@     �C@      �?      A@     �K@      "@      @      �?      H@      c@      $@      g@      @      @      (@      ;@      f@     �\@      @      Q@       @                              @                      8@                                      @      "@               @      �?                              @                      &@                                      @      �?              �?      �?                                                      *@                                       @       @              �?      X@      .@      @      (@      <@     �l@      ,@     }@      $@      �?     �A@      3@     `q@     �g@      @     �^@      "@                      �?              <@              (@                       @       @      0@      2@              *@      @                                      �?                                                      @      �?               @      @                      �?              ;@              (@                       @       @      (@      1@              &@     �U@      .@      @      &@      <@     `i@      ,@     P|@      $@      �?     �@@      1@     `p@     �e@      @     �[@      >@      $@      @      @      @      W@      @     �i@      @              "@       @      \@      L@      �?      1@     �L@      @      @      @      6@     �[@       @     �n@      @      �?      8@      .@     �b@      ]@      @     @W@     �I@      @      $@       @      6@     �i@      "@      z@       @      @      @       @     @o@     @^@      @      D@      2@               @              �?      C@      �?      L@                       @      �?      ;@      A@              "@      1@              �?              �?      5@      �?      C@                       @      �?      0@      *@              "@      @              �?                      3@              6@                       @              *@      @              @      (@                              �?       @      �?      0@                              �?      @      $@              @      �?              �?                      1@              2@                                      &@      5@                      �?              �?                      @              2@                                      $@      *@                                                              $@                                                      �?       @                     �@@      @       @       @      5@     �d@       @     �v@       @      @      @      @     �k@     �U@      @      ?@      8@      @       @       @      4@     �b@       @     �r@      @      �?      @      @     �i@     �U@       @      =@      0@       @      @      @      0@     @R@      @     �Z@      �?      �?       @      �?     �T@     �D@              4@       @       @      �?      @      @     �R@       @     �g@      @              @      @      _@     �F@       @      "@      "@                              �?      3@              O@      @      @              �?      0@      �?      �?       @       @                              �?      @              7@      @                      �?      @      �?      �?              �?                                      *@             �C@      �?      @                      (@                       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJt�;hhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx         
                    �?���P��?�	           ��@       	                    !@�͝�6b�?U           ��@                          �:@�S�kZ�?O           ��@                           �?�����`�?�           �@������������������������       ��q���?<           �~@������������������������       �mMN1C�?�           h�@                           �?Ʌ�5��?�            `n@������������������������       �[�>��?             ?@������������������������       �j�����?{            �j@������������������������       ��zv��?             &@                           @�����?z           "�@                           �?����X��?L           Ȍ@                           �?�����?W            �a@������������������������       ��J#��P�?>            �X@������������������������       ��|���?             F@                          �2@���U��?�           X�@������������������������       ���]�`��?�             j@������������������������       �r�� ��?j           ؁@                           @dd�x���?.           ��@                           @�H�pkn�?9           ��@������������������������       �� ��w��?D           x�@������������������������       ���O�s��?�            �v@                            �?�������?�            �w@������������������������       �9��8���?�             h@������������������������       �ߗ���?r            @g@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@     �@@      D@      ?@      X@     X�@      B@      �@      .@      (@     �R@     �Q@     �@     �@      8@     �q@     @Y@      1@      @@      *@      I@      s@      7@     0x@      &@      @      B@      C@     r@     �m@      (@      d@      Y@      1@      @@      *@     �H@     s@      3@     0x@      &@      @      B@      C@     r@     `m@      (@     �c@     �U@      (@      =@      *@     �F@     `q@      *@      t@      $@      @      ?@     �B@     �n@     �i@      &@     �^@      4@      @      3@      �?      (@     �W@      �?     �\@      @      �?      &@      @     �R@     �U@       @      F@     �P@      "@      $@      (@     �@@     �f@      (@     �i@      @      @      4@     �@@     @e@     @^@      "@     �S@      *@      @      @              @      ;@      @     �P@      �?              @      �?     �F@      <@      �?     �B@      �?              �?                       @              (@                      @              @      @               @      (@      @       @              @      9@      @     �K@      �?              �?      �?      E@      6@      �?     �A@      �?                              �?      �?      @                                                       @               @      Z@      0@       @      2@      G@     �u@      *@     (�@      @      @     �C@      @@      |@      q@      (@     �^@      H@       @      @      "@      9@     �]@      @     �q@      @      �?      &@      2@     �j@     �Y@      @      O@      @                       @      @      0@              ?@                      �?      @      H@      @              4@      @                       @      @      ,@              4@                      �?      @      =@      @              *@      �?                               @       @              &@                                      3@       @              @      E@       @      @      @      4@     �Y@      @      p@      @      �?      $@      (@     �d@     �W@      @      E@      1@              @      �?      @     �@@              L@                       @      @     �M@      1@       @      &@      9@       @      @      @      1@     @Q@      @      i@      @      �?       @       @     �Z@     �S@       @      ?@      L@       @      �?      "@      5@     `l@      "@     `z@              @      <@      ,@     `m@     @e@       @      N@      @@      @      �?      @      *@     �c@      @     Pr@              @      0@      "@     `g@      _@      @     �A@      ;@      �?      �?      @      $@     �V@      @     @d@              �?      @      @     @^@     �O@      @      :@      @       @              @      @      Q@       @     ``@              @      "@       @     �P@     �N@      @      "@      8@      @               @       @     @Q@      @      `@                      (@      @      H@      G@       @      9@      @      @                      @      A@              S@                       @       @      @@      ,@      �?      0@      1@      �?               @      @     �A@      @     �J@                      $@      @      0@      @@      �?      "@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJI	hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?LW~�'��?�	           ��@       	                    @tsk��?9           �@                           @~��5a�??           �@                          �0@��i|��?�           \�@������������������������       ��C�kRy�?+            �Q@������������������������       ���B����?�           @�@                           �?%������?�            �l@������������������������       ��A��_�?M             a@������������������������       ���� ��?6             W@
                           @�
i��?�            `x@                            @�K���?�             w@������������������������       ���k���?�            Pq@������������������������       ����-�?:            @W@                          �5@�������?             4@������������������������       �4և����?             @������������������������       ��q-��?             *@                           �?�M����?^           �@                           @<����9�?�            �u@                          �=@�����?�            @l@������������������������       �P�vz"�?�             k@������������������������       �X�<ݚ�?             "@                            �?�	�.,4�?I            �]@������������������������       ��P^Cy�?.             S@������������������������       ���0��=�?            �E@                            @'�_����?�           ��@                          �@@�BE�)��?4           �@������������������������       �%���1��?.           ē@������������������������       �      �?              @                           @��2@l��?R           ��@������������������������       �DGX�܁�?I           8�@������������������������       �
ףp=
�?	             .@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@     �E@     �B@      4@     @X@      �@      C@     ��@      &@       @     @Y@     �O@     ��@     `@      6@     �o@      V@      :@      :@      &@     �J@     �r@      4@     �z@      @      @     �H@      <@     0t@     `n@      $@     �]@      O@      3@      6@      $@      I@     @l@      "@      t@      @      @      G@      5@     �p@     �f@      @     �W@      H@      3@      4@       @     �D@     `h@      @     �q@      @      @      C@      3@     @j@     �a@      @     �R@       @       @       @      �?      "@      @      @      @              �?       @      �?      2@      ,@              @      G@      1@      2@      @      @@     �g@      @     @q@      @       @      B@      2@      h@     �_@      @     @Q@      ,@               @       @      "@      ?@       @      E@                       @       @     �K@     �D@              4@      $@               @      �?      @      *@       @      0@                       @              @@      ?@              .@      @                      �?      @      2@              :@                               @      7@      $@              @      :@      @      @      �?      @     @R@      &@      Z@      �?              @      @      M@      O@      @      8@      :@      @      @      �?       @     �Q@      "@     @Y@      �?              @      @      L@     �K@      @      6@      0@      @      @      �?      �?     �L@       @     �P@      �?              �?      @     �D@     �E@      @      6@      $@       @                      �?      *@      �?     �A@                       @       @      .@      (@                                                      �?      @       @      @                                       @      @               @                                              �?       @      �?                                       @                      �?                                      �?       @               @                                              @              �?      Z@      1@      &@      "@      F@     �u@      2@     ��@      @      @      J@     �A@     0{@     0p@      (@      a@      6@      �?      @              .@     �I@      �?      [@                       @             �K@     �H@      @      @@      (@      �?      @              @     �B@             �Q@                       @              D@      9@              <@      &@      �?      @              @     �B@             @P@                       @              C@      9@              <@      �?                                                      @                                       @                              $@              @               @      ,@      �?     �B@                                      .@      8@      @      @      @                              @       @              <@                                      (@      ,@       @      �?      @              @               @      @      �?      "@                                      @      $@      �?      @     �T@      0@      @      "@      =@     `r@      1@     `�@      @      @      I@     �A@     �w@     @j@      "@     @Z@     �P@      (@      @      @      8@     �i@      1@     0v@       @      @      F@      8@     @n@     �d@       @     �V@     �P@      (@      @      @      8@     @i@      1@     0v@       @      @      F@      6@      n@     �d@       @     �V@                                              @                                               @      �?                              0@      @               @      @     �U@              m@      @      �?      @      &@     @a@     �F@      �?      ,@      0@      @               @      @     �T@             �l@      @      �?      @      &@     �`@      D@      �?      ,@                                              @               @                                      @      @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�RyhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @d�N ��?�	           ��@       	                    �?gڼ����?�           �@                           �? 7�'{�?�            �x@                          �0@f)�(�e�?`            �c@������������������������       ��zv��?             &@������������������������       ��h���?Z            @b@                           @r���*�?�            �m@������������������������       �¦	^_�?`            `c@������������������������       ��!�Mq�?9            �T@
                          �;@�?є��?�           ��@                            �?�K�x�?j           &�@������������������������       ������L�?�           @�@������������������������       �&����o�?�           ,�@                           �?�Z���E�?�            `m@������������������������       ��5`��_�?6            �T@������������������������       �D�n�3�?\             c@                           @5Gv��@�?�           �@                           �?z{���?*           p|@                           �?���j��?�            �o@������������������������       ��o�h��?K            �[@������������������������       �r��:�j�?]            �a@                           �?ey�F���?�            `i@������������������������       ���/2��?T            �_@������������������������       �6�80\��?.             S@                           @3\Yc�K�?�           Ѓ@                          �8@��@=aP�?|           ��@������������������������       ��5p`S�?            {@������������������������       ��J���?m            �e@������������������������       ���zۧ��?             ;@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        g@     �@@      C@      8@      [@     ��@      F@     ��@      <@      @      S@      Q@     �@     �@      1@      r@     @b@      :@      =@      2@     �T@     �|@      C@     8�@      6@      @     @P@     �L@     �~@     �w@      .@     `n@      6@       @      @      @      *@     �B@             �\@      @              *@      @     @U@     �I@              C@      "@      �?      @       @      @      @              J@      @              &@      @      =@      .@              .@                      @                                      �?                               @      @       @                      "@      �?      �?       @      @      @             �I@      @              &@       @      :@      *@              .@      *@      �?               @      @     �@@             �O@                       @       @      L@      B@              7@      "@      �?              �?      @      :@             �@@                       @       @      E@      0@              2@      @                      �?      �?      @              >@                                      ,@      4@              @      _@      8@      9@      ,@     �Q@     �z@      C@     ��@      2@      @      J@     �I@     py@     �t@      .@     �i@     �\@      1@      8@      *@     �N@      x@      A@     ��@      1@      @      G@      H@     �w@     0s@      *@     @h@      @@      &@      @      "@      *@     �e@      $@     �j@      @              $@      $@     �`@     �Z@      @     �D@     �T@      @      4@      @      H@     �j@      8@     @t@      $@      @      B@      C@     �n@      i@       @      c@      $@      @      �?      �?      "@      C@      @      W@      �?              @      @      =@      5@       @      &@       @      @      �?              @      $@              ;@                      �?               @      *@              @       @      @              �?       @      <@      @     @P@      �?              @      @      5@       @       @      @      C@      @      "@      @      9@      i@      @     �w@      @              &@      &@     �j@      `@       @     �G@      0@       @       @      @      @     �N@      �?     �d@       @              $@       @     @[@     �G@              7@      @              @      @      �?     �A@             @Y@       @              @       @      H@      <@              ,@      @              @                      1@              C@       @              @       @      7@      $@              @                              @      �?      2@             �O@                      @              9@      2@              @      &@       @      @      �?       @      :@      �?      P@                      @             �N@      3@              "@      &@       @                       @      2@      �?      ;@                      @              E@      ,@              @                      @      �?               @             �B@                                      3@      @               @      6@      @      �?              6@     �a@      @     �j@      @              �?      "@      Z@     �T@       @      8@      6@      @      �?              6@     �_@      @     �i@      @              �?      "@      Y@      T@       @      6@      0@       @      �?              0@     @V@      @     @c@      @              �?      "@     �L@      M@       @      4@      @      @                      @      C@             �J@                                     �E@      6@               @                                              *@              @                                      @       @               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�fRKhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @���m%|�?�	           ��@       	                     �?V�5v��?�           ��@                            �?-f�D)��?.           :�@                           @3H�u(�?t           8�@������������������������       ����K��?�           ��@������������������������       ����\�?�            �p@                           @�`݉6��?�           X�@������������������������       �M��>��?�            �@������������������������       �F]t�E�?             6@
                           �?�f�����?�           ��@                          �7@8�xsr��?�            t@������������������������       ��
�;���?�            �n@������������������������       ��Q,K��?-            �R@                           @�p^���?�            �w@������������������������       �ü�i�?{            �h@������������������������       �4� �^��?o            �f@                           @�̔�?�           ��@                           �?P�,�I�?G           p�@                           �?�E9l9�?�           8�@������������������������       �f�% �
�?{            @i@������������������������       �6�`�B��?7           �}@                           �?��%х;�?�            �l@������������������������       ���0q��?G            �Z@������������������������       �������?N            @_@                           �?���>4��?�             l@                          �7@t��B�u�?G            �\@������������������������       ��@�ܠ�?8            �W@������������������������       �H�z�G�?             4@                           @F���/�?D            @[@������������������������       �>4և���?&             L@������������������������       ��84�a��?            �J@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      A@      A@      9@     �X@     ��@      ?@     ܐ@      ,@      @      Q@      Q@     p�@      �@      1@     p@     �b@      >@      =@      7@     �S@     ��@      <@     h�@      "@       @     �N@      L@     p@      w@      1@      j@     �[@      7@      3@      1@      J@     @z@      6@     ��@      @             �A@      =@     �x@     �o@      &@     `a@      J@      @       @      "@      8@     �f@      "@     r@       @              @      $@     �g@      `@      @      K@     �E@      �?       @      @      0@     �a@      @      k@       @              @       @     @b@     @R@      @      D@      "@      @              @       @      E@      @      R@                      @       @      E@      L@      �?      ,@      M@      0@      1@       @      <@     �m@      *@     �o@      @              =@      3@      j@     @_@      @     @U@      M@      0@      1@       @      <@     �m@      (@     @o@      @              =@      3@      i@     �]@      @     �T@                                                      �?      @                                       @      @              @     �C@      @      $@      @      :@     �[@      @     �a@       @       @      :@      ;@     �Z@      ]@      @     �Q@      3@      @      @       @      $@     �J@      @     @R@      �?       @      @      1@      A@      M@      @      <@      ,@      @      @       @      @     �F@      @     �E@      �?      �?      @      ,@      <@     �E@      @      :@      @                              @       @      �?      >@              �?              @      @      .@               @      4@       @      @      @      0@     �L@      �?     �Q@      �?              5@      $@      R@      M@      @      E@      "@       @       @      �?      @      4@             �C@      �?              (@      @     �I@      ;@       @      9@      &@               @      @      (@     �B@      �?      ?@                      "@      @      5@      ?@      �?      1@     �H@      @      @       @      5@      h@      @     �x@      @      @      @      (@     �n@     �a@              H@     �H@       @      @      �?      2@     @c@       @     �r@      @      @      �?      &@     �i@     @\@             �D@     �B@       @      @      �?      .@     �Y@      �?     `m@      @      @      �?      @     `b@     �U@             �@@      &@               @              @      B@      �?     �M@                              @      C@      @@              *@      :@       @      �?      �?       @     �P@              f@      @      @      �?      @     @[@      K@              4@      (@              �?              @     �I@      �?     �P@                              @      M@      ;@               @      @                               @      ?@      �?      3@                              @      6@      *@               @      @              �?              �?      4@             �G@                                      B@      ,@                               @      �?      �?      @      C@      �?     @W@                      @      �?      E@      =@              @               @      �?      �?      @      3@      �?      B@                      @              ;@      0@              @              �?              �?       @      2@      �?      =@                      @              2@      0@              @              �?      �?              �?      �?              @                                      "@                                                                      3@             �L@                      @      �?      .@      *@              �?                                              @              ?@                              �?      (@      @                                                              *@              :@                      @              @      @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���%hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�v�3#��?�	           ��@       	                    �?޸'�?�           ��@                          �=@&F�|�?           ��@                            �?�#�:���?�           ؒ@������������������������       �OTT��H�?B           X�@������������������������       �2�5����?�            �r@                           @���WV�?             J@������������������������       �9��8���?             8@������������������������       �      �?             <@
                           @E2|�v��?�           ��@                           @������?�           \�@������������������������       ��/��f��?�           ��@������������������������       ��������?�            �y@                          �0@
ףp=
�?            y@������������������������       �46<�R�?             9@������������������������       �v8�Jw��?�            pw@                           �?&���Z,�?�           ��@                           @�[���?            @h@                           @�:˛��?c            �b@������������������������       �sp��P��?4            �T@������������������������       ��]�l�?/             Q@                           @� ��H��?            �E@������������������������       �dh����?            �A@������������������������       �      �?              @                          �:@A�ww���?J           ��@                           �?�/,� �?�           0�@������������������������       ����|O�?�             x@������������������������       �h(�׿��?�            @x@                           �?,�Ra���?a             f@������������������������       ��"���?9            �Y@������������������������       �B����k�?(            �R@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@     �@@      G@      @@     @^@     ��@      =@     d�@      .@      $@     �X@      R@     @�@     P~@      4@     �n@     �e@      :@     �C@      =@      W@     �}@      9@     P�@      &@      @     @T@      K@     �|@     Pv@      .@     �i@     @V@      &@      =@      .@     �K@      n@      1@     0r@       @      @     �C@      ;@      h@     �a@      @     �W@     �T@      &@      =@      .@     �H@     �m@      1@     �p@       @      @     �C@      ;@      h@     @`@      @     @W@     �P@      @      8@      &@      ;@      g@      (@     �j@      @      �?     �B@      4@     �b@     �U@       @     �N@      .@      @      @      @      6@      J@      @      K@      @      @       @      @     �E@      F@      @      @@      @                              @      @              7@                                      �?      $@              �?       @                              @      @              .@                                                                      @                               @      �?               @                                      �?      $@              �?      U@      .@      $@      ,@     �B@     �m@       @     pz@      @       @      E@      ;@     �p@      k@      $@      \@     @R@      $@       @      *@      >@     �g@      @     �r@      @              @@      1@     `i@     �a@      @     �T@     �G@      $@      @      @      4@     @^@      @      e@                      2@      $@      c@     �V@       @     �I@      :@              @       @      $@     �Q@      @      `@      @              ,@      @     �I@     �I@      @      ?@      &@      @       @      �?      @     �G@      �?     �_@               @      $@      $@     �P@      S@      @      >@      @                                      @              �?                                      @      (@              �?      @      @       @      �?      @      F@      �?     �_@               @      $@      $@     �O@      P@      @      =@     �C@      @      @      @      =@     �g@      @     �x@      @      @      2@      2@     @o@      `@      @      C@       @               @               @      H@      �?      I@                      @              C@      7@              (@      @               @              @      C@      �?     �D@                      @              >@      *@              (@      �?              �?               @      6@              8@                       @              3@      "@              @      @              �?              �?      0@      �?      1@                       @              &@      @              "@      �?                              @      $@              "@                                       @      $@                      �?                               @      "@              @                                      @      $@                                                      @      �?              @                                      �?                              ?@      @      @      @      5@     �a@      @     �u@      @      @      ,@      2@     �j@     @Z@      @      :@      :@      @      @      @      ,@     �\@      @     �p@      @      �?      ,@      .@     �f@      X@              8@      0@      @      @       @      @     @P@      �?     �`@      @      �?      @      @      R@     �L@              *@      $@      �?      �?      �?      &@      I@       @     �`@                      $@      "@     �[@     �C@              &@      @       @                      @      <@             �T@              @              @      =@      "@      @       @      @                              �?      (@             �J@              @              @      *@      @      @       @               @                      @      0@              >@                                      0@      @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJr^hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?+������?�	           ��@       	                    �?1U�#�<�?�           ��@                            @��W��I�?k           p�@                           @ԻK	��?�            �s@������������������������       �譎���?�            �r@������������������������       �ֳC��2�?             6@                          �1@t�F�Y�?�             q@������������������������       �5��g�?            �A@������������������������       ��?����?�            �m@
                            @{��m�?f           ��@                          �4@m��d�t�?l            �@������������������������       ���v�P��?s            �g@������������������������       �L�1�j�?�            px@                           @����O�?�            �x@������������������������       ��W�?�            �r@������������������������       ��i�d��?9            @X@                            @����հ�?�           R�@                           �?����5�?�           `�@                           @t�чj�?A           X�@������������������������       ���r��?�           ؅@������������������������       ��n_Y���?�             j@                          �1@Vk��Ś�?q           h�@������������������������       �JeΚV�?z            `g@������������������������       �������?�           ��@                           �?�8����?4           }@                           �?��%��?T            @^@������������������������       �YE�t�?-            �P@������������������������       ��*���?'            �K@                           @>@�?��?�            �u@������������������������       �     ��?S             `@������������������������       �@�9S˅�?�             k@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@      A@      ?@      6@      ^@     ��@      F@     T�@      0@      ,@     �Q@     @Q@     P�@     �@      :@      n@     �V@      ,@      *@      $@     �F@      n@      *@      @      @      @      >@      4@     pq@     �h@      *@      X@      C@      "@      &@      @      ;@      X@      @     @b@       @      @      (@      "@      Y@     @S@      @      G@      1@      @      @      @      5@      M@      @      Q@      �?              $@      @      E@      C@      @     �B@      (@      @      @      @      5@     �K@      @      P@      �?              $@      @      A@      C@      @     �A@      @                                      @              @                                       @                       @      5@      @      @              @      C@      �?     �S@      �?      @       @      @      M@     �C@      @      "@       @              �?               @       @              @                      �?       @      @      @               @      3@      @      @              @      >@      �?     �R@      �?      @      �?      �?     �I@      @@      @      @     �J@      @       @      @      2@      b@      "@     �u@      @              2@      &@     `f@     @^@      @      I@     �E@       @              @      (@     @U@      "@      e@       @              0@      @     @\@     @S@      @     �B@      *@                       @             �A@      @     �F@                       @              J@      5@      �?      (@      >@       @               @      (@      I@      @      _@       @              ,@      @     �N@      L@      @      9@      $@      @       @      @      @      N@             �f@       @               @      @     �P@      F@       @      *@      "@      @       @      @      @      B@             �b@       @               @       @      I@      <@              &@      �?                              �?      8@             �@@                               @      0@      0@       @       @     @[@      4@      2@      (@     �R@     Pz@      ?@     (�@      $@      &@     �D@     �H@     0}@     ps@      *@      b@     @Y@      *@      1@      (@     �P@     pu@      :@     �{@       @      &@      B@     �E@     0v@     `p@      *@     @`@     �K@      "@      "@      @      D@      f@      $@     �f@      @      $@      (@      4@      d@     �^@      "@     @T@      E@      "@      @      @      9@     @_@      "@     @b@      @       @      (@      3@      _@     �V@      "@     �P@      *@               @       @      .@      J@      �?     �B@               @              �?     �B@      ?@              .@      G@      @       @      @      :@     �d@      0@     Pp@      @      �?      8@      7@     @h@     �a@      @     �H@      ,@      �?      �?      @              D@       @      J@                      �?      "@      7@      ?@              $@      @@      @      @      @      :@     �_@      ,@      j@      @      �?      7@      ,@     `e@     @[@      @     �C@       @      @      �?              "@     �S@      @      e@       @              @      @      \@     �H@              ,@      @      �?                              5@              ?@                      @              C@      .@              @      @      �?                              .@              $@                      @              3@       @              @      �?                                      @              5@                                      3@      @              �?      @      @      �?              "@     �L@      @     @a@       @              �?      @     �R@      A@               @       @       @                      @      5@      @     �A@                              @      B@      ,@              @      �?      @      �?              @      B@      �?     �Y@       @              �?              C@      4@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?>?����?�	           ��@       	                    @��B��?E           ��@                           �?<:ț0
�?E           x�@                          �0@�{�q��?s            `f@������������������������       �s
^N���?	             ,@������������������������       ��qg_�S�?j            �d@                           @��d���?�           ��@������������������������       ��ٳ���?M           ��@������������������������       ��8%���?�            �j@
                          @@@�q7����?            �x@                           @'��c���?�            pw@������������������������       ��h^����?�            �p@������������������������       ��E��Y�?K            �[@������������������������       �ҳ�wY;�?             1@                            @9q��(�?X           F�@                          �;@?��6���?�           d�@                           @�����?h           l�@������������������������       �@$�U��?�           @�@������������������������       �s��o��?�           ��@                           @v�R���?w            �g@������������������������       �؋�Ð(�?b            �c@������������������������       �>��R	�?             ?@                           �?^D��h�?y           P�@                           @�Ѥs%�?�            0w@������������������������       ������?�            @q@������������������������       ��\4Jȫ�?7            �W@                          �2@�$ێ���?�            �j@������������������������       ���V��?.            �Q@������������������������       �h/���v�?`             b@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �l@      @@     �C@      6@     �]@     @�@      ?@     ,�@      &@      $@      U@     �I@     ��@      �@      ;@      q@     �]@      1@      @@      &@      O@     @r@      ,@     z@      @      @      @@      <@     Ps@     @k@       @     �`@     @V@      (@      :@      &@      M@     �m@      @     �t@      @      @      <@      7@     �n@      `@      @     @[@      0@              @      �?      "@      0@              L@                      "@      @      7@      9@              0@                      �?              �?                      �?                      @      @      �?      @                      0@               @      �?       @      0@             �K@                      @       @      6@      5@              0@     @R@      (@      7@      $@     �H@     �k@      @      q@      @      @      3@      2@     �k@     �Y@      @     @W@      K@      &@      2@      @      C@     �g@      @     `l@      @      @      1@      2@      e@     �S@      @      S@      3@      �?      @      @      &@      ?@             �G@                       @             �J@      9@              1@      >@      @      @              @      L@       @     �U@      @              @      @     @P@     �V@      @      9@      <@      @      @              @      L@       @      U@      @              @      @     @P@     �S@      @      9@      6@      @      @              �?     �E@      @     @P@      @              @      @     �B@      K@      @      &@      @               @              @      *@      �?      3@                                      <@      8@              ,@       @                                                      @                                              (@                     @[@      .@      @      &@     �L@     @v@      1@     P�@      @      @      J@      7@     0z@     `r@      3@     @a@     @W@      (@      @      "@      H@     @q@      *@     �z@      @      @     �G@      4@     �q@      n@      1@      _@     @U@      &@      @      "@      G@     �l@      &@     w@       @      @     �E@      0@     �o@     @l@      *@     �[@     �H@      @       @      @      7@     �]@       @     �e@      �?              (@      @     �]@      S@      @     �I@      B@      @      @      @      7@     �[@      "@     @h@      �?      @      ?@      "@     �`@     �b@      "@      N@       @      �?                       @     �G@       @     �N@      �?              @      @      =@      ,@      @      *@       @      �?                       @      E@       @     �E@      �?              @      @      7@      ,@      @      *@                                              @              2@                      �?      �?      @                              0@      @       @       @      "@      T@      @     �o@       @      �?      @      @      a@      K@       @      ,@      (@       @       @       @      @      L@      @      c@       @      �?      @      @      S@      @@       @      ,@       @       @       @       @      @     �@@      @     �^@       @      �?      @      @     �L@      0@              *@      @                                      7@              >@                                      3@      0@       @      �?      @      �?                      @      8@             �X@                                     �N@      6@                       @                                      @              :@                                      ?@      @                       @      �?                      @      1@             @R@                                      >@      1@                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�`HhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @���l�?�	           ��@       	                   �<@NR����?�           "�@                            �?C�#��?a           l�@                           �?��KJ��?T           �@������������������������       ������?a             e@������������������������       �`���}�?�           Ј@                            �?�� ��?           ̙@������������������������       ��TI��?           ؏@������������������������       �:�!i�?�           ��@
                            �?�|���?�            `k@                           �?z������?B            �Y@������������������������       �������?	             *@������������������������       �Y�JV���?9            @V@                           �?�x��?G            @]@������������������������       ���8��8�?             8@������������������������       �����Bx�?:            @W@                           �?F�U��?�           ��@                          �2@��k���?t             f@                          �1@UUUUU�?             H@������������������������       �`������?             7@������������������������       �U���N@�?             9@                           @     ��?U             `@������������������������       �����?A            �W@������������������������       �xC�Ҁ��?            �@@                          �2@`YV;3�?=           @�@                           @N�jo�?�             o@������������������������       ���lL��?r            @g@������������������������       �^�/��#�?)            �O@                          �3@M�����?�           x�@������������������������       �j�@u��?9            @V@������������������������       ��=�]@�?i           ��@�t�b�[     h�h4h7K ��h9��R�(KKKK��h��B�       �i@      ;@      D@      6@      [@     ��@      A@     Б@      7@      @      T@     �P@     ��@     0~@      .@      o@     �d@      3@      ;@      2@      X@     0~@      >@     ��@      1@      @     @Q@      L@     ��@     �v@      *@     �j@      d@      2@      ;@      2@     @W@     �{@      ;@     �@      0@      @     �M@     �H@     �~@     �u@      (@     �h@     �I@      @      @      "@      3@      f@      (@     �r@      @              "@      $@     @g@     @[@      @      M@      @       @               @      @      3@      @      N@                       @              E@      ,@              ,@      F@      @      @      @      .@     �c@      "@     `n@      @              @      $@      b@     �W@      @      F@     @[@      *@      8@      "@     �R@     �p@      .@     @u@      "@      @      I@     �C@     Ps@     �m@      @     �a@      P@      @      .@      @     �E@     �f@      "@     `l@      @       @      2@      7@     �j@     �a@      @     �P@     �F@      $@      "@      @      ?@     �U@      @     @\@      @      @      @@      0@     @X@      X@       @     �R@      @      �?                      @     �B@      @      U@      �?              $@      @      A@      2@      �?      ,@                                       @      .@       @     �H@      �?                       @      0@      &@              @                                              @               @                                      @       @              �?                                       @      $@       @     �G@      �?                       @      *@      "@              @      @      �?                      �?      6@      �?     �A@                      $@      @      2@      @      �?      $@      @                                      @               @                      @      @      @      �?                       @      �?                      �?      3@      �?     �@@                      @      �?      &@      @      �?      $@      D@       @      *@      @      (@      f@      @     �y@      @              &@      &@     @l@     @]@       @     �B@       @              @              @     �@@             �I@                      @       @      @@      <@              (@      �?              �?              @      "@              5@                      @       @      @       @               @      �?                              �?      @              @                       @       @      @       @              �?                      �?               @      @              .@                      �?              �?                      �?      @              @                      8@              >@                                      <@      :@              $@      @              @                      4@              8@                                      7@      &@              $@      @                                      @              @                                      @      .@                      @@       @      "@      @      "@     �a@      @     �v@      @               @      "@     @h@     @V@       @      9@      @              @       @      �?     �F@      @     �S@                      �?      @     �R@      :@              @      @              @       @      �?     �A@             �J@                               @     @P@      1@              @       @                                      $@      @      :@                      �?       @      $@      "@                      ;@       @      @       @       @     �X@      �?     �q@      @              @      @     �]@     �O@       @      6@      @      @                              @              J@                                      $@       @               @      4@      @      @       @       @     �V@      �?     �l@      @              @      @     @[@     �K@       @      4@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�$�LhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @��!s�?�	           ��@       	                    @B�����?�           إ@                           �?�A�9��?           (�@                            �?Ҝ%�y�?s           �@������������������������       ����
<��?           `y@������������������������       �ϸ�����?f            �e@                            �?�$M�N�?�           8�@������������������������       ���xp	��?9           `@������������������������       ��8���!�?c             b@
                            �?^^���?�           ��@                           @̗�P��?d           8�@������������������������       ��ZR[q�?           �{@������������������������       �&�;Y-o�?R            �a@                           �?t�v(;�?t           ؎@������������������������       ����]��?P            �\@������������������������       ����M.�?$           @�@                           @��p��?�           t�@                           @@G����/�?7           P}@                           �?���ҝ=�?/           �|@������������������������       ���λ�Z�?�            �k@������������������������       �H��.��?�            @m@������������������������       ��؉�؉�?             *@                          �5@�7�N��?�           @�@                          �3@U2�5T�?�            �s@������������������������       ��0jB��?y             g@������������������������       ��,�F.�?K            �`@                          �;@�A*�\|�?�            �t@������������������������       ��\	ͭ��?�            @l@������������������������       �E�V�.{�?A            @Z@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @e@     �@@      C@      5@     @[@     ��@     �B@     ȑ@      8@       @      Q@     �Q@     ��@     8�@      5@     �p@     ``@      9@      ?@      .@     �V@     }@      ?@     �@      3@      @     �N@      J@     �}@     �y@      4@      m@      P@      1@      3@      (@     �F@     �j@      @     `s@      $@       @      5@      8@     @n@     �`@      @      Y@      >@      $@      *@      $@      ;@      \@      @      `@      @       @      &@      (@      W@     @P@      �?     �L@      6@      @      &@      @      ,@     �T@      @     �X@      @              &@      @     �S@     �A@              >@       @      @       @      @      *@      >@              >@       @       @              @      *@      >@      �?      ;@      A@      @      @       @      2@     �Y@       @     �f@      @              $@      (@     �b@     �Q@      @     �E@      :@      @               @      &@     �T@       @      c@      @              @      $@     �\@      I@      @      @@       @      �?      @              @      5@              =@                      @       @     �A@      4@      �?      &@     �P@       @      (@      @     �F@     @o@      :@     pz@      "@      @      D@      <@      m@      q@      .@     �`@      2@      @      @       @      (@     �U@      *@     @h@      @              @      "@     @V@     �X@      @      C@      (@       @      @       @      @     �R@      &@     �`@      @              @      @     �Q@     @T@              ?@      @      @                      @      &@       @     �N@                              @      2@      1@      @      @     �H@      @       @      �?     �@@     �d@      *@     �l@      @      @      A@      3@     �a@      f@      "@     �W@      @                      �?      @      3@              5@      @              �?             �B@      *@       @      @      E@      @       @              <@      b@      *@      j@       @      @     �@@      3@     �Z@     `d@      @     �V@     �C@       @      @      @      3@     �h@      @     Py@      @      �?      @      2@      o@     �[@      �?      C@      1@      �?      @      @      @     @P@       @      g@              �?      @      @      \@     �F@              0@      1@      �?      @      @      @     @P@       @      f@                      @      @      \@     �F@              0@      &@      �?      @              @     �D@       @      S@                      @      �?     �E@      9@              (@      @               @      @      �?      8@              Y@                      �?      @     @Q@      4@              @                                      @                      "@              �?                                                      6@      @      �?       @      (@     �`@      @     �k@      @              @      ,@      a@     @P@      �?      6@      *@       @      �?       @      "@      E@      @     �\@       @              @       @     �P@      @@              2@      "@       @      �?       @      @      ;@       @      L@                      @       @     �H@      2@              $@      @                              @      .@       @      M@       @                      @      2@      ,@               @      "@      @                      @      W@             �Z@      @                      @     @Q@     �@@      �?      @       @      @                       @     �P@              O@                              @      J@      =@              �?      @                              �?      9@              F@      @                              1@      @      �?      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��jhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?t,�Փ�?�	           ��@       	                     �?����5=�?=           8�@                           �?��:O �?           �x@                           �?h3F��(�?^            �b@������������������������       ��"w����?%            �L@������������������������       �"*w�?9             W@                           ?@�f����?�             o@������������������������       �l;�z��?�            �m@������������������������       �.y0��k�?             *@
                           @ףp=Jx�?8            �@                           @Wb��q�?�           ��@������������������������       �>q9]�?�           h�@������������������������       ����4�h�?�            �w@                            �?�5yb[�?�            �j@������������������������       �K�=�U�?=             Y@������������������������       ����ٓ�?E            �\@                            @SJs���?|           v�@                          �0@S�3�%}�?�           �@                           @[�vuT�?6            �R@������������������������       ��f���?)            �K@������������������������       �333333�?             4@                            �?b�{*�f�?�           ؗ@������������������������       �����g��?�           ��@������������������������       �"\Ź�O�?�            �w@                          �3@ch)�w-�?~           Ѓ@                           �?��.GA�?{            �h@������������������������       �֭pw���?H            �]@������������������������       �^�^��?3            �S@                           @hO�ll��?           P{@������������������������       �@��+�?�            �n@������������������������       �r�q?�?m             h@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @i@      ?@      G@      >@     �Z@     ��@      >@      �@      7@      @      R@     @P@     8�@     ��@      4@      p@     @Z@      *@      =@      "@     @R@     �q@      .@     y@      (@      @     �C@      =@     @s@     �i@      @     `b@      7@      �?       @      @      $@     @P@      @      `@      �?              (@      @      P@      I@      �?      <@      *@              �?       @       @      ?@      @     �A@                      @      @      6@      .@              .@      �?              �?              �?      @              0@                      @      @      $@      @              $@      (@                       @      �?      9@      @      3@                                      (@      (@              @      $@      �?      �?       @       @      A@      �?     �W@      �?              @              E@     �A@      �?      *@      $@      �?      �?       @       @     �@@      �?     �T@      �?              @              E@      A@      �?      *@                                              �?              &@                                              �?                     �T@      (@      ;@      @     �O@      k@      $@      q@      &@      @      ;@      :@     �n@     �c@      @     �]@     �P@      (@      :@      @     �D@     �e@      @     �l@      &@      @      6@      :@      j@      `@      @     �Y@      C@      "@      5@       @     �A@      ]@      �?     �a@      @      @      0@      &@     @b@     �Q@       @      P@      =@      @      @      �?      @      L@      @     �U@      @              @      .@     �O@      M@      @      C@      .@              �?       @      6@      F@      @      E@                      @             �A@      ;@              1@      $@              �?              0@      1@      @      .@                      @              6@      @              @      @                       @      @      ;@       @      ;@                       @              *@      5@              $@     @X@      2@      1@      5@      A@     �u@      .@     x�@      &@      @     �@@      B@     0}@     `t@      *@     �[@     �S@      *@      0@      2@      :@     �o@      (@     {@      "@             �@@      =@     �t@     �n@      &@     �V@      @                      @              $@              @                       @      @      2@      5@              @      @                      @              "@              @                       @      @      .@      "@              @       @                                      �?              �?                                      @      (@              �?     @R@      *@      0@      .@      :@     @n@      (@     �z@      "@              ?@      :@     �s@     @l@      &@     �T@      M@      $@      @      *@      ,@      h@      "@     pv@      "@              3@      0@     �m@     �b@      @      J@      .@      @      $@       @      (@      I@      @      Q@                      (@      $@     �S@      S@      @      ?@      3@      @      �?      @       @     �W@      @     �o@       @      @              @     �`@     �S@       @      5@      *@              �?       @      @      6@      �?     @R@                                     �I@      <@               @      &@              �?       @      @      (@      �?      F@                                      4@      8@              �?       @                              �?      $@              =@                                      ?@      @              �?      @      @              �?      @      R@       @     �f@       @      @              @     �T@     �I@       @      3@      @      �?              �?      @      =@             �^@       @      @              @     �E@      4@              *@      @      @                             �E@       @      M@                              @     �C@      ?@       @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��#6hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @fU=��?�	           ��@       	                    �?dI��?�           �@                          �=@�Rpl�?+           ,�@                            �?���2v�?           t�@������������������������       �P%�
��?M           ��@������������������������       ���Qn�,�?�            �r@                           @�fl ��?             G@������������������������       �r`�����?             C@������������������������       �      �?              @
                            �?
�*HΠ�?�           �@                           @8�U��?�           �@������������������������       ����	�?           ؉@������������������������       �ܴ�L��?�            �t@                           @]��έ�?�            �w@������������������������       �{�	d�?�            0t@������������������������       ��>4և��?#             L@                           �?/c.��?�           �@                           �?�<�(�5�?,           �~@                           @�Ӝ)��?�            `l@������������������������       ����l�?i            `e@������������������������       ���)x9�?             L@                           @����?�            �p@������������������������       �ء�wN��?L            �`@������������������������       ��X��(�?X            �`@                          �2@���2�?o           h�@                           �?� {�/��?Y             a@������������������������       �/k��\�?-             Q@������������������������       ��paRC4�?,             Q@                           @���i��?           P|@������������������������       �������?c             d@������������������������       ���J���?�            @r@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      :@     �E@      =@     @^@     Ȅ@     �B@     \�@      2@       @     �T@     �N@      �@     �@      4@     p@      b@      3@     �B@      <@      Y@     �@      =@     �@      .@       @     �Q@     �I@     �@     �w@      4@      j@      T@      @      =@      (@      I@     @o@      ,@     �q@      $@      @      >@      ;@     �j@     @d@      @     �\@      S@      @      =@      (@      G@      o@      ,@     Pp@      $@      @      >@      ;@      j@     �b@      @     �\@      J@      @      5@      &@     �A@     `i@      $@      k@      @       @      4@      *@     �c@     �Z@      @     @T@      8@      �?       @      �?      &@     �F@      @      F@      @      @      $@      ,@     �I@      F@       @      A@      @                              @       @              5@                                      @      &@                      @                              @       @              2@                                      @      @                                                                              @                                              @                     @P@      (@       @      0@      I@     �o@      .@     pz@      @      @     �D@      8@     `r@     `k@      ,@     �W@     �F@      (@      @      ,@      <@     `h@      (@     �v@      @              3@      (@      n@     @c@      @      I@      C@      @      @       @      0@      c@      @     @m@      @              ,@       @     �f@     �[@      @     �C@      @      @              @      (@      E@      @     ``@                      @      @      M@      F@              &@      4@              @       @      6@      N@      @      M@      �?      @      6@      (@     �J@     @P@      "@      F@      1@              @       @      ,@     �K@      @     �H@      �?      @      4@      (@     �D@     �N@      "@      ?@      @                               @      @              "@                       @              (@      @              *@     �F@      @      @      �?      5@      d@       @     `y@      @              (@      $@     @m@     �^@              H@      ;@       @      @              0@      U@      @     �a@       @               @      @     �Y@     �P@              <@      ,@      �?      �?              @     �@@       @      M@                      @             �O@      >@              ,@      (@      �?      �?              @      6@       @     �D@                      �?              L@      5@              $@       @                              �?      &@              1@                      @              @      "@              @      *@      �?      @              &@     �I@      @     @U@       @               @      @     �C@     �B@              ,@      @               @              &@      =@             �F@                      �?      @      1@      (@              @      @      �?       @                      6@      @      D@       @              �?      �?      6@      9@              @      2@      @      �?      �?      @      S@      �?     pp@      �?              @      @     �`@      L@              4@      @                      �?              .@             �H@                       @              F@      1@              @      @                      �?               @              :@                                      *@      *@              @      �?                                      @              7@                       @              ?@      @                      *@      @      �?              @     �N@      �?     �j@      �?               @      @      V@     �C@              1@       @              �?              @      *@              U@                       @      @      >@       @              *@      &@      @                              H@      �?     @`@      �?                      @      M@      ?@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJHa�^hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @3j0�hy�?�	           ��@       	                    @���_7��?           &�@                           �?��+��?#            �@                          �?@�}R�݆�?O           ؍@������������������������       �t�����?A           �@������������������������       �VUUUUU�?             8@                           �?�{�ƹ��?�           T�@������������������������       ��rE���?           �z@������������������������       ��}@VT�?�           h�@
                          �;@@�H�Q�?�           �@                           @������?�           h�@������������������������       �:��:�?B           �@������������������������       �"P7��?o            `e@                           @K�z���?7            �U@������������������������       �ZQl�R�?            �G@������������������������       �?;���x�?            �C@                           �?��x�<��?�           ؐ@                          �2@�#qW��?�            ps@                           �?�Ks�g��?D            �Y@������������������������       �ͯ�
��?"            �J@������������������������       �4��7���?"             I@                           �?ֻ�����?�             j@������������������������       �gr��
�?Q            �[@������������������������       ��b��P��?<            @X@                          �2@�������?�           ��@                           @�O�2���?q             f@������������������������       �x�$!]�?O            @`@������������������������       ��яǆ�?"            �G@                           @r;!�4��?k           p�@������������������������       �̻��)��?B           `�@������������������������       ���;�JB�?)            �P@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@      ?@     �E@      =@     @[@     p�@      B@     ��@      ,@      $@      T@      N@     ��@     P�@      3@     �o@     �b@      5@     �A@      7@     @W@     P~@      <@     8�@      *@       @     @Q@      H@     p~@     �x@      0@      k@      _@      .@      8@      3@     @S@     �u@      .@     X�@      $@      @     �K@      D@     �w@     �p@      (@     �b@     �N@      @      5@      &@      K@     @d@       @     @k@      "@      @      <@      .@     �d@     �Z@      @     @S@      N@      @      5@      &@      K@      c@       @     �i@      "@      @      <@      .@     �d@     �Z@      @     @S@      �?                                      $@              (@                                              �?                     �O@       @      @       @      7@     `g@      @     s@      �?              ;@      9@      j@      d@       @     �R@      :@      @              �?      @      S@      �?     �W@                      $@      (@     @X@      N@      @      @@     �B@      @      @      @      0@     �[@      @     @j@      �?              1@      *@      \@     @Y@      @      E@      ;@      @      &@      @      0@      a@      *@     �k@      @       @      ,@       @     �[@     ``@      @     @P@      ;@      @      &@      @      0@      ^@      *@     �e@      @       @      *@       @     �Y@     �]@      @     �O@      7@      @      "@      @      $@      X@      *@     �^@      @       @      &@      @     @U@     �U@      @      B@      @      �?       @              @      8@              J@                       @      @      2@      @@              ;@                                              0@              G@                      �?               @      *@               @                                              $@              6@                                      @      (@                                                              @              8@                      �?              @      �?               @     �D@      $@       @      @      0@      e@       @     px@      �?       @      &@      (@      n@     �^@      @      B@      ,@      @      �?       @      @      D@              X@                      @      @     �T@      B@              6@      @              �?       @              &@              =@                                     �D@      $@              @       @              �?       @              @              0@                                      .@       @               @      @                                      @              *@                                      :@       @               @      "@      @                      @      =@             �P@                      @      @     �D@      :@              2@      @      @                      @      1@              8@                      @      @      9@      0@               @       @                               @      (@             �E@                       @              0@      $@              $@      ;@      @      @      @      &@      `@       @     pr@      �?       @      @       @     �c@     �U@      @      ,@      @               @      @      @     �A@       @      H@                      @       @     �E@      5@              @      @               @      @      @      8@              9@                      @       @     �A@      3@              @                                              &@       @      7@                      �?               @       @                      5@      @      @      �?      @     �W@      @     �n@      �?       @              @      ]@     �P@      @      "@      5@      @      @      �?      @     �V@      @     �k@      �?       @              @      Y@      H@      @      "@              �?                              @              ;@                                      0@      2@                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ7]jXhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?,ia�j�?�	           ��@       	                    �?�B?���?           ��@                            �?��(\�Y�?�            �@                          �1@q=
ף0�?�             t@������������������������       �h+�v:�?-             Q@������������������������       �k���?�            �o@                           @�����U�?�             t@������������������������       �D˩�m��?`            �b@������������������������       �������?e            �e@
                          �2@̬.o�)�?t           @�@                          �1@���i��?y            `j@������������������������       ���`��?G            �\@������������������������       �r�qw�?2             X@                           @~�K��?�            Py@������������������������       �����
��?�            Pu@������������������������       �     ��?)             P@                           �?�铤'�?�           ¤@                            @�Z�	�?�           L�@                          �=@>�C�uV�?�           P�@������������������������       ����Zg�?�           �@������������������������       ���RT��?            �C@                           @OA���?�            �r@������������������������       �%!ɧ�a�?�            �h@������������������������       �C４�$�?B            �X@                            @J�%�ci�?�           8�@                            �?ci�5�?�           @�@������������������������       ���2� �?           ��@������������������������       �wona��?�            @q@                          �2@$ܔM��?7           �@������������������������       � �j���?E             ]@������������������������       ���f݄"�?�            �x@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @i@      5@     �H@      8@     �Z@     0�@      :@     ��@      0@      "@      R@      O@     �@      �@      0@     �o@     @T@      @      (@      (@      E@      i@      @     �s@      &@              7@      >@      p@     �e@      @     �U@     �A@      @      "@      $@      :@     @^@      @     �a@       @              1@      *@     @\@     @T@      @     �K@      2@              @      @      *@      O@       @     �T@      @              &@      @     �G@     �A@      �?      9@       @               @              �?      .@              @       @              �?      @      1@      0@              @      0@              @      @      (@     �G@       @     �S@      @              $@      @      >@      3@      �?      4@      1@      @      @      @      *@     �M@       @     �M@       @              @      @     �P@      G@       @      >@      @               @              @      A@      �?     �@@      �?              �?      �?      7@      6@              2@      &@      @       @      @      @      9@      �?      :@      �?              @      @     �E@      8@       @      (@      G@      �?      @       @      0@     �S@       @     �e@      @              @      1@      b@     �V@              @@      8@              �?      �?      �?      <@              D@                       @      @     �Q@      @@              @      .@              �?                      *@              ?@                       @      @      @@      ,@              @      "@                      �?      �?      .@              "@                               @      C@      2@              @      6@      �?       @      �?      .@     �I@       @     �`@      @              @      (@     �R@     �M@              9@      5@      �?       @      �?      (@      A@       @     �]@      @              @      $@      P@      K@              .@      �?                              @      1@              .@                               @      &@      @              $@     @^@      0@     �B@      (@     @P@     �{@      4@     p�@      @      "@     �H@      @@     �@     �u@      *@     �d@     �M@      &@      8@      �?      E@     @h@       @     0p@      @      @      ,@      .@     �e@      b@      @     �T@     �E@       @      2@      �?      <@     �a@       @     @d@      @      @      (@      &@     �^@     �Z@      @      R@     �D@       @      2@      �?      9@      a@       @     `b@      @      @      (@      &@      ^@     �W@      @      R@       @                              @      @              .@                                      @      &@                      0@      @      @              ,@     �J@             @X@               @       @      @      I@     �C@      �?      $@      0@       @      @              @     �C@              M@               @       @      @      <@      >@      �?      @              �?      �?              @      ,@             �C@                                      6@      "@              @      O@      @      *@      &@      7@     �o@      (@     X�@              @     �A@      1@     �t@     �h@       @     @U@      K@      @      "@      "@      1@     �b@      (@     v@              @      >@      (@     @k@     �c@       @     �Q@     �A@       @      @      "@       @     �\@      $@     `r@                      $@      @     `f@     �[@      @     �E@      3@      �?      @              "@      A@       @     �M@              @      4@      @     �C@      G@      @      <@       @       @      @       @      @     �Y@             @i@                      @      @      ]@     �E@              ,@      �?              �?                      6@             �@@                      @       @     �@@      .@              @      @       @      @       @      @     @T@              e@                              @     �T@      <@              $@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��?*hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �1@ԋ"s��?�	           ��@       	                     �?���(�?�           ��@                          �0@��� ���?e             e@                           @&1����?&            �O@������������������������       ���~1���?            �D@������������������������       �袋.���?             6@                           �?�sl����??            �Z@������������������������       �
"����?             ?@������������������������       ��۱�5�?-            �R@
                            @�5 
��?*           �~@                            �?������?�            �v@������������������������       ��0��>�?            �i@������������������������       �.c�R��?[            @c@                           @D>�Q�?P            @`@������������������������       �K����?8             W@������������������������       �^.��?             C@                           !@	�E�c�?           j�@                          �;@Q�ژb�?           H�@                           �?�kb����?           J�@������������������������       ��Q$�Cg�?           �{@������������������������       �D0k؆}�?�           Ң@                          �>@��?�72�?�            �w@������������������������       �G�)��\�?�            �p@������������������������       �n ��X�?J            �]@                          �9@|�l�]�?             1@������������������������       ����(\��?             $@������������������������       �����>4�?             @�t�bh�h4h7K ��h9��R�(KKKK��h��B�        j@     �@@      E@      1@     �Z@     H�@      ?@     4�@      ,@      @      U@      R@     ��@     �@      5@     0p@     �F@      @      (@      @      .@     �]@      $@      d@      �?       @      ,@      ,@     @V@      \@      @      J@      @              @       @      @      <@      @     �P@                      �?      �?      6@      7@              @                               @      �?      (@       @      ,@                      �?              *@      .@              @                               @      �?      (@       @       @                                      *@       @              �?                                                              (@                      �?                      @               @      @              @              @      0@      @      J@                              �?      "@       @              @       @              @                      @      @      ,@                                      �?                              �?                              @      &@      �?      C@                              �?       @       @              @      E@      @      @      �?      &@     �V@      @     �W@      �?       @      *@      *@     �P@     @V@      @     �F@      A@      @      @      �?      &@     �Q@       @      M@      �?       @      &@      $@     �E@     �P@      @      A@      1@       @      @              @     �D@             �D@      �?      �?      @      �?      >@      C@      �?      0@      1@      @              �?      @      =@       @      1@              �?      @      "@      *@      =@      @      2@       @      �?                              5@       @      B@                       @      @      8@      6@              &@      @      �?                              .@              3@                       @      @      3@      3@              "@      @                                      @       @      1@                                      @      @               @     �d@      ;@      >@      ,@      W@     ��@      5@     h�@      *@      @     �Q@      M@     ��@     �x@      .@     �i@     �d@      ;@      >@      ,@     �V@     P�@      5@     X�@      *@      @     �Q@      M@     �@     �x@      .@     �i@      b@      5@      :@      *@      T@     P~@      4@     ��@      (@      @     @P@      L@     ��@     �v@      &@     �g@      ,@      �?      @              5@     �M@             �^@      @              $@             @W@     �P@       @      F@     @`@      4@      4@      *@     �M@     �z@      4@      �@       @      @     �K@      L@     �}@     �r@      "@      b@      4@      @      @      �?      &@     @Q@      �?     �a@      �?      �?      @       @     �Q@      =@      @      2@      &@      @      @      �?      @     �D@             @[@      �?              @              I@      2@       @      (@      "@                              @      <@      �?      ?@              �?      �?       @      5@      &@       @      @                                      �?       @               @                                      �?      @              �?                                      �?      @                                                              @                                                              @               @                                      �?                      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ?�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �1@�s�:�z�?�	           ��@       	                   �0@њ}?|(�?�           x�@                           @*St�ó�?�            �h@                           @�64k0�??            �V@������������������������       ��D�M��?4            �Q@������������������������       �u#����?             3@                           �?N���9�?A            �Z@������������������������       ��ĳ����?#             N@������������������������       ��TA�>��?             G@
                           �?B~��%�?           �z@                            �?IV�A��?�            @j@������������������������       �U�x?r��?!             F@������������������������       �P�?i            �d@                           @������?�             k@������������������������       ���x0Ta�?p             f@������������������������       �R���Q�?             D@                            @z�8I�?           ��@                            �?K�"���?�           ,�@                          �;@�Ӱ���?3           ��@������������������������       ��V�� �?�           p�@������������������������       �+ʤ��I�?T            �`@                           @�iL�?�           �@������������������������       �/l;�c�?.           4�@������������������������       ��[�E�h�?S            �]@                           @�2����?a            �@                           �?:?I�q��?
           �y@������������������������       ���"�/p�?�            pp@������������������������       ����Y�?d            �b@                           @P&:�.w�?W           0�@������������������������       �齁�ne�?o            �e@������������������������       �������?�            �w@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `h@      A@      G@      :@     @]@     ��@     �@@     p�@      8@      @     �P@     �I@     �@     ��@      0@     @o@     �L@              (@       @      &@     @^@      "@     @`@      �?      �?      ,@      &@     @\@     �V@      @     �G@      &@                       @      @      G@      @      >@      �?      �?      �?      @     �B@      D@      �?      ,@      @                      �?       @      >@       @       @      �?              �?      �?      5@      1@              @      @                      �?       @      8@       @      @      �?              �?      �?      *@      *@              @                                              @              �?                                       @      @                       @                      �?      �?      0@      @      6@              �?              @      0@      7@      �?      &@      @                              �?      @      @       @              �?               @      "@      ,@      �?       @       @                      �?              "@              ,@                              �?      @      "@              @      G@              (@               @     �R@      @      Y@                      *@      @      S@     �I@       @     �@@      :@              $@              @      E@      @      =@                      @      @      ?@      ;@       @      6@      @               @               @      @      �?      $@                              @      @      @              @      7@               @              @     �A@       @      3@                      @      @      ;@      4@       @      1@      4@               @              �?     �@@      �?     �Q@                       @      �?     �F@      8@              &@      4@               @              �?      ?@              M@                      @      �?      A@      8@              @                                               @      �?      *@                      @              &@                       @     @a@      A@      A@      8@     �Z@     ��@      8@     Ў@      7@      @      J@      D@     ��@     �{@      *@     `i@      Z@      ;@      8@      6@      V@     y@      3@     ��@      2@       @     �E@     �A@     0y@     Pt@      (@     �e@      8@      (@       @      *@      ;@     `d@      @     r@       @              &@      @     `e@     `a@      @     �B@      7@      (@       @      *@      3@     �b@      @      l@      @              $@      @     @b@      `@      @      @@      �?                               @      .@             @P@      �?              �?              9@      &@              @      T@      .@      6@      "@     �N@     �m@      *@     Pu@      $@       @      @@      =@      m@     @g@      @      a@     �S@      .@      4@      "@     �M@     �l@      (@     �r@      "@       @      ;@      <@     �i@      e@      @     �^@      �?               @               @      "@      �?     �D@      �?              @      �?      9@      2@              *@      A@      @      $@       @      2@     `a@      @     @v@      @      �?      "@      @     �k@     �]@      �?      >@      2@      @      "@       @       @     �A@      @     @c@                      @      @     �Y@     �I@              1@      *@               @      �?      @      3@      @     @[@                      �?      @     �I@      ?@              .@      @      @      �?      �?      �?      0@             �F@                      @              J@      4@               @      0@      @      �?              $@      Z@      �?     @i@      @      �?      @      �?      ^@      Q@      �?      *@      @      �?                       @     �D@              K@       @               @              A@      2@              @      "@      @      �?               @     �O@      �?     �b@      @      �?      �?      �?     �U@      I@      �?      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ/	hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�G��W��?�	           ��@       	                     @Ic(�<�?^           8�@                            �?(���y�?1           ��@                           @+#��'<�?d            �@������������������������       ��L����?�           ��@������������������������       �[�9���?�            @u@                           �?ų8ֵ�?�            �t@������������������������       �~�Q���?             3@������������������������       �����T��?�            �s@
                           @w�r�?-           �}@                          �<@���}���?�            �t@������������������������       �
߬:���?�            �q@������������������������       �ҽ��?            �E@                           @ʖî,E�?`            �b@������������������������       �>F?�!��?             E@������������������������       �XB1B&�?E            �Z@                          �;@,C�V���?l           ��@                           @��#��?�           ĝ@                            @�b>��?(           (�@������������������������       �W���Y��?�           ��@������������������������       �ì�~?�?�            �n@                            �?� �X�	�?�           0�@������������������������       ��
���?d           `�@������������������������       ���|s�?6            ~@                           @���.u�?�            �p@                           �?��@!���?�            `j@������������������������       �C)��,��?            �H@������������������������       ��4�/�j�?h            @d@                          �=@�4#`�v�?#            �K@������������������������       �ҳ�wY;�?             1@������������������������       ��k(����?             C@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `l@      @@     �C@      <@     �Z@     ��@      =@     $�@      4@      $@     �O@     �R@     �@     P�@      .@      p@     �^@      1@      <@      *@      N@     �s@      3@     �y@      *@      @      9@      D@     �r@      n@      "@     @`@     �U@      $@      1@      (@      H@      m@      2@      q@      (@      @      5@      A@     �i@     �f@      "@      Y@     @P@      @      ,@      &@     �@@     �f@      &@     �k@       @      �?      3@      5@     �c@     �[@      @     @P@      D@       @      &@       @      7@     @[@       @     @c@      @              &@      *@     @Z@      P@      @      D@      9@      @      @      @      $@     �Q@      "@     �P@      @      �?       @       @      K@     �G@      �?      9@      6@      @      @      �?      .@     �J@      @      J@      @      @       @      *@     �G@     @Q@       @     �A@                      �?              �?                      @       @                              @                      @      6@      @       @      �?      ,@     �J@      @      H@       @      @       @      *@     �D@     @Q@       @      >@     �A@      @      &@      �?      (@     @T@      �?      a@      �?      �?      @      @     �V@     �N@              >@      ?@      @      $@               @      L@      �?     �V@      �?      �?       @      @      J@      G@              2@      ,@      @      $@               @     �J@      �?     @T@              �?       @      @     �F@     �E@              0@      1@                                      @              $@      �?                              @      @               @      @              �?      �?      @      9@              G@                       @             �C@      .@              (@       @                              �?      @              .@                                      "@      @              @       @              �?      �?      @      5@              ?@                       @              >@      "@              @     @Z@      .@      &@      .@     �G@     �u@      $@     ��@      @      @      C@     �A@     @{@     �q@      @     �_@     �W@      ,@      &@      .@     �F@     pr@      "@     ��@      �?      @     �A@      >@      y@     �p@      @     �\@     �F@      @      @       @      5@     �_@      �?     �n@                      ,@      .@      k@     �W@       @     �P@     �B@      @      @      @      5@     �Y@      �?     �c@                      &@      $@      b@     �Q@       @     �K@       @              @      @              9@              V@                      @      @     @R@      8@              (@      I@      $@      @      @      8@      e@       @     t@      �?      @      5@      .@     �f@     @e@      @      H@      3@      @      @      @      (@     @W@      @     �f@                      "@      @     @\@     �S@      �?      9@      ?@      @      �?       @      (@     �R@      @     @a@      �?      @      (@      "@     �Q@      W@       @      7@      $@      �?                       @     �I@      �?      ^@      @       @      @      @      B@      1@      �?      &@      $@      �?                       @      A@      �?      Z@               @      @      @      5@      1@      �?      &@      @      �?                      �?      $@              (@                               @      @      "@              @      @                              �?      8@      �?      W@               @      @       @      2@       @      �?      @                                              1@              0@      @                      �?      .@                                                                      @              (@                                       @                                                                      ,@              @      @                      �?      *@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJU�$hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@�"�2�e�?�	           ��@                           �?�$����?g           �@                           @ELI�+�?�           �@                            @O��,�?�           ��@������������������������       �����Fw�?�           �@������������������������       �)i)�D/�?           �z@������������������������       �l�l��?	             .@                            @1w)�>��?�           Н@	       
                    @�R�~1m�?W           0�@������������������������       �����+�?�           (�@������������������������       ���ށ��?�           8�@                           @�ځ�v�?Q           @�@������������������������       ��t��7��?�            `o@������������������������       ��v��?�            �r@                           @����T��?$           �}@                           @�Uj>�?�            `y@                           @����̍�?�            �t@������������������������       ��8�QF%�?�             p@������������������������       ��"e����?)             R@                          �=@q9W��S�?3             S@������������������������       �"sLj�'�?            �D@������������������������       ����:��?            �A@                           �?J�q"���?'            �P@                            �?��$�<u�?            �A@������������������������       �T#G�h�?             7@������������������������       ��8��8��?             (@                           @     ��?             @@������������������������       �      �?             8@������������������������       �      �?              @�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      8@     �B@      8@     �Y@     Ȅ@     �A@     \�@      .@       @      T@     �F@     ��@     �@      .@     �m@      i@      4@     �@@      8@     �W@     (�@      @@     Ќ@      (@      @     �Q@      E@     �@     0}@      ,@     �j@     @X@      &@      8@      "@     �L@     �q@      0@     �u@      "@      @      =@      6@     @r@     �h@       @     �_@     @X@      &@      8@      "@     �L@     Pq@      *@     pu@      "@      @      =@      6@      r@     �h@       @     �_@     @S@      @      .@      @      E@     �h@      &@      l@       @      @      8@      2@     @h@     �a@       @     @[@      4@      @      "@       @      .@      T@       @     �]@      �?              @      @     �W@     �K@              2@                                              @      @       @                                      @                             �Y@      "@      "@      .@     �B@     �r@      0@     �@      @              E@      4@     �y@     �p@      @      V@      T@      @      @      ,@     �@@     �k@      &@     �w@      @             �C@      2@     q@      i@      @     �Q@      E@      @      @      &@      "@      [@      @     �g@      @              *@      &@     �f@     �W@       @      ?@      C@       @      �?      @      8@      \@       @     `g@                      :@      @     �V@     �Z@      �?      D@      7@      @       @      �?      @     �S@      @      i@                      @       @     �a@     �Q@      @      1@      .@                      �?      �?      9@              W@                       @      �?     �R@      =@              $@       @      @       @              @     �J@      @      [@                      �?      �?     �P@     �D@      @      @      4@      @      @               @      U@      @     �g@      @      �?      "@      @     �T@      C@      �?      8@      4@      @      @               @     �S@      @     @b@      @      �?       @      �?     �Q@      B@      �?      6@      (@      @       @              @     �O@      @     �`@      �?      �?       @      �?      I@      ?@      �?      ,@      "@      @       @              @     �G@      @     �W@      �?      �?       @      �?      H@      2@      �?      *@      @                                      0@             �B@                                       @      *@              �?       @               @              �?      .@              ,@       @                              5@      @               @      @               @                      @               @                                      $@      �?               @      �?                              �?      $@              @       @                              &@      @                                                              @             �E@                      �?       @      &@       @               @                                              @              .@                      �?       @       @       @               @                                              @              @                      �?       @       @       @               @                                              �?              &@                                                                                                              �?              <@                                      @                                                                      �?              6@                                      �?                                                                                      @                                       @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�.�VhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?,7��|~�?�	           ��@       	                   �;@NU��E�?           0�@                           �?rnlQ�?�           ��@                          �6@���o��?�            �j@������������������������       �#W��{�?a             c@������������������������       �������?!            �M@                          �8@�P啣S�?5           <�@������������������������       ��3`�h�?�           ��@������������������������       ��֟�g�?h            �d@
                           @���9Q��?g             e@                            �?d>j����?S            �`@������������������������       ��7x,�?            �D@������������������������       ��3�U�?9            @W@                          �<@K��o!`�?            �A@������������������������       ���!pc�?             &@������������������������       ��q�q�?             8@                          �;@���)��?�           z�@                           !@�8�[��?�           <�@                            @�cb���?�           �@������������������������       ���A�h�?}           ĕ@������������������������       ��x0��?F           ��@������������������������       ��5��?             *@                          �<@K:8p�a�?�            �r@                           @     ��?)             P@������������������������       ��g�`�|�?            �B@������������������������       ���ͦ-��?             ;@                           @6�ɿ��?�            �m@������������������������       �b@�ܻ�?6            @U@������������������������       ���l��?Y             c@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      C@     �B@      7@     �]@     ��@      A@     �@      .@      @     �W@      P@     ȅ@     �~@      4@     �p@     @S@      7@      8@      &@      Q@     �r@      1@     Px@      *@      @      A@     �C@      r@      m@      *@     @a@     �O@      5@      7@      &@     �N@     �q@      1@     �t@      (@      @      7@     �C@     0p@     `k@      *@     �_@      @      @       @      @      $@      9@       @      N@       @               @      @     �C@      >@              0@      @      @                      "@      .@       @      I@       @               @      @      <@      &@              *@                       @      @      �?      $@              $@                                      &@      3@              @      L@      2@      5@       @     �I@      p@      .@     �p@      $@      @      .@      A@     �k@     �g@      *@     �[@     �H@      .@      5@      @      I@     �i@      $@     �n@       @      @      .@      @@     �h@     @d@      *@      X@      @      @              �?      �?      K@      @      ;@       @                       @      7@      ;@              .@      ,@       @      �?              @      3@              M@      �?              &@              ?@      ,@              &@      &@       @      �?              @      2@             �C@      �?              &@              8@      "@              &@                                      @      @              3@                                      @       @              @      &@       @      �?              @      *@              4@      �?              &@              3@      @              @      @                                      �?              3@                                      @      @                      �?                                      �?              "@                                                                       @                                                      $@                                      @      @                     �\@      .@      *@      (@     �I@     pv@      1@     ��@       @      �?     �N@      9@     py@      p@      @     ``@     @Z@      *@      *@      (@      H@     �r@      *@     ��@      �?      �?      J@      4@     �v@     �n@      @     @]@     @Z@      *@      *@      (@      H@     Pr@      *@     ��@      �?      �?      J@      4@     pv@     `n@      @     @]@     �T@      (@       @      $@     �C@     �j@      $@     �z@      �?      �?      H@      2@      o@      f@      @     �W@      6@      �?      @       @      "@     @T@      @      i@                      @       @     �[@     �P@              6@                                              "@               @                                      �?      �?                      "@       @                      @     �L@      @      a@      �?              "@      @     �G@      ,@      �?      ,@       @                                       @              A@                       @              *@      @              �?       @                                      @              0@                                      &@      @              �?                                              @              2@                       @               @      �?                      @       @                      @     �H@      @     �Y@      �?              @      @      A@      $@      �?      *@      @       @                      @      2@      @      9@      �?              @      @      "@       @      �?      "@       @                                      ?@      �?     @S@                      @      �?      9@       @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJE�chG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@_��>��?�	           ��@       	                     @1(ah��?�           ��@                            �?�}��)�?           j�@                           @W�.h���?�           8�@������������������������       ����7��?D           ،@������������������������       ����I��?I           ��@                           @9	����?�           8�@������������������������       �,�<��~�?w            �g@������������������������       ��>����?           �z@
                          �2@���#�?l           H�@                           @Ӝ��� �?�            `q@������������������������       ���s���?z             i@������������������������       �#l^��?4            �S@                           �?jR��c�?�           ��@������������������������       ���+e`�?�            �s@������������������������       �G�����?�            pw@                           �?b�U�x��?!           �|@                          @@@�Q�ߧ��?o            `e@                           �?���� �?c             c@������������������������       ��K~���?             >@������������������������       �l>/���?T            �^@                           @��[��"�?             2@������������������������       �      �?              @������������������������       ���Q��?             $@                           �?uk~X��?�             r@                            @�W���?m            `f@������������������������       ��X�N��?G            @[@������������������������       �����S�?&            �Q@                           @���w˕�?E            @[@������������������������       �Stvn|�?9            @W@������������������������       �     ��?             0@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `j@      ?@      D@      >@     @[@     P�@      G@     ,�@      0@      "@     �U@     �Q@     �@     0�@      &@     �k@     �g@      :@      C@      >@     �Y@     �@      E@     ��@      &@      @     �Q@      O@     ��@     �@      "@     `i@     �a@      1@      >@      :@     �U@     �{@      C@     ��@      $@      @     �O@      K@     �z@     �v@       @      f@     @X@      (@      4@      6@     �J@     0v@      <@     �~@      @             �E@      D@      t@     Pp@      @     �\@     �P@      @      (@      &@      5@      e@       @     �k@      @              3@      .@     �g@      `@      @      J@      >@      @       @      &@      @@     @g@      4@     �p@      @              8@      9@     �`@     �`@      @     �O@     �F@      @      $@      @      A@      V@      $@      Z@      @      @      4@      ,@     @Z@     @Z@       @     �N@       @      @      @               @      8@       @      5@                      $@      @      D@      D@              9@     �B@      �?      @      @      :@      P@       @     �T@      @      @      $@       @     @P@     @P@       @      B@      G@      "@       @      @      0@     �`@      @     Pt@      �?       @      @       @     �l@     `b@      �?      ;@      "@      �?      @      @      @      9@      �?     �Y@                      �?      @     �T@      @@              "@       @              @      @              *@              S@                      �?      �?     �Q@      1@              @      �?      �?                      @      (@      �?      :@                               @      (@      .@               @     �B@       @      @              $@     �[@      @     �k@      �?       @      @      @     `b@     �\@      �?      2@      <@      @      @              @      J@      �?     �S@               @      @      @      L@     �P@              "@      "@      @       @              @      M@       @      b@      �?               @       @     �V@      H@      �?      "@      7@      @       @              @      R@      @     �f@      @       @      1@       @     @S@     �B@       @      2@      3@      @       @               @      0@             �N@       @              "@       @      <@      0@              $@      0@      @       @               @      .@             �J@       @              "@       @      <@      $@              $@       @                                      �?               @                      @              &@      �?              �?      ,@      @       @               @      ,@             �F@       @              @       @      1@      "@              "@      @                                      �?               @                                              @                                                              �?              @                                               @                      @                                                      @                                              @                      @      �?                      @      L@      @      ^@      @       @       @      @     �H@      5@       @       @      @      �?                      @     �A@      @      T@               @      �?      @      9@      *@       @      @      @      �?                      �?      6@      @     �@@                      �?      @      6@      &@       @      @                                       @      *@             �G@               @                      @       @              �?                                      �?      5@              D@      @              @       @      8@       @              @                                      �?      4@              <@      @              @       @      5@       @              @                                              �?              (@                                      @                        �t�bub�"     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���PhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @4il���?�	           ��@       	                    @r<�9	�?           &�@                           �?
 �:P�?*           0�@                            �?e��\��?N           ȍ@������������������������       �wZ����?�            Pt@������������������������       ��/��?�           ��@                            �?�q?̌�?�           |�@������������������������       �Ղp��?,           ؊@������������������������       �Hfh�Fp�?�            @p@
                          �0@� ����?�           ؇@                           �?r�q��?             H@������������������������       ��ˠT�?             6@������������������������       �G���ջ�?             :@                            �?<�G_��?�           X�@������������������������       ��Ŝ�?�            @m@������������������������       �IE�8�?&           ~@                           �?�	\�v��?�           ؐ@                           �?��;�f�?�           Ȃ@                           @�m��v�?�             m@������������������������       �MƻL��?z            �f@������������������������       ���+e��?              I@                           @:��]��?�             w@������������������������       �,�2aȽ�?f             c@������������������������       ���Q0�x�?�            �j@                          �5@w��ޝ��?+           �}@                           @Pf��r��?�            �q@������������������������       ��a�fG�?�             l@������������������������       ��.���S�?(             O@                           @�4���.�?{            �g@������������������������       �0�
K�z�?5            �U@������������������������       �	j*D�?F             Z@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �f@      B@      B@      @@     @X@     8�@     �F@     �@      (@      @     �S@      Q@     ��@     �@      6@     �q@     @b@      3@      >@      ;@     �S@     p~@     �C@     �@      $@      @     @Q@     �L@     P�@      x@      4@     �m@     @\@      0@      9@      8@      P@     �u@      5@     H�@      @      @     �M@     �E@     �w@     �m@      *@     �h@     �K@      "@      1@      1@      D@     �d@      $@     @i@      @      @      <@      5@     �d@     �\@       @     �V@      5@      �?               @       @      P@       @     @[@       @              "@       @     �J@      8@      �?      5@      A@       @      1@      .@      @@     �Y@       @     @W@       @      @      3@      *@      \@     �V@      @     �Q@      M@      @       @      @      8@     �f@      &@     �s@      �?              ?@      6@     �j@     @^@      @     �Z@      G@      @       @      @      *@     �b@      "@     0p@      �?              3@      0@     �e@     �V@      @     �O@      (@      �?      @      @      &@      @@       @      N@                      (@      @     �D@      >@              F@     �@@      @      @      @      .@      a@      2@     �f@      @              $@      ,@     �a@     �b@      @     �D@       @              �?              �?      &@              @                                      @      6@      �?                              �?              �?      @               @                                      @       @      �?               @                                      @               @                                      @      ,@                      ?@      @      @      @      ,@     �_@      2@      f@      @              $@      ,@      a@      `@      @     �D@      @       @      @      @       @     �A@      @     �P@                      @       @      J@     �H@       @      @      <@      �?      �?              (@     �V@      ,@     @[@      @              @      (@      U@     �S@      @     �A@     �B@      1@      @      @      2@      d@      @     Px@       @       @      "@      &@     @n@      `@       @     �E@      :@      $@      @      @      @     �T@      �?     �k@      �?       @      @      @      ^@     �R@       @      @@      2@      @      @              @      ?@             @P@      �?      �?      @      �?     �I@      @@      �?      (@      ,@       @      @              @      ;@              G@      �?              @      �?      E@      8@      �?      &@      @      @                              @              3@              �?                      "@       @              �?       @      @      �?      @              J@      �?     �c@              �?      @      @     @Q@      E@      �?      4@      @              �?       @              1@             @R@              �?      @              =@      *@              &@      @      @               @             �A@      �?      U@                              @      D@      =@      �?      "@      &@      @       @      �?      &@     @S@      @     �d@      �?               @      @     �^@     �K@              &@      @      @       @      �?      @      A@      �?     �\@                      �?      @      S@      :@              @      @      @       @      �?      @      ?@      �?     @T@                      �?       @      P@      6@              @      �?      @                       @      @             �@@                              @      (@      @              �?      @                              @     �E@      @     �J@      �?              �?              G@      =@              @      @                               @      @              :@                      �?              <@      ,@              @                                       @     �B@      @      ;@      �?                              2@      .@                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJٞzWhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @���Co�?�	           ��@       	                    �?x�����?�           ��@                           @t�b���?           l�@                          �1@�����?�           �@������������������������       � ��~٢�?�            @m@������������������������       �F0$��?           ؈@                          �;@�^C�v�?~            �j@������������������������       ���"B<�?u            �h@������������������������       �     ��?	             0@
                           @y3�W03�?�           ��@                          �=@jp4\J�?�           ��@������������������������       ���%3h��?r           H�@������������������������       ��w����?            �D@                          �;@w/�>o�?.           ��@������������������������       �$� �/S�?�           x�@������������������������       ��v:����?P             a@                           @����?�           �@                           �?8�9#5�?R           �@                          �0@{��,��?�            0x@������������������������       �9��8���?             (@������������������������       �ľ(��a�?�            pw@                           @J!���?Y           ��@������������������������       �	�%���?<           �~@������������������������       ��8��8��?             H@                           �?������?�            �l@                          �4@�1�g
�?L            @\@������������������������       �v�*� ��?*            �O@������������������������       ����Mb�?"             I@                           @*���ت�?D            �\@������������������������       ��@*���?            �A@������������������������       ���(\���?/             T@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@      ?@      K@      4@     @U@     ؄@     �@@     ��@      2@      *@     �S@      L@     ��@     p~@      :@     �o@     �c@      :@     �C@      2@      O@     P}@      :@     `�@      *@      $@     �P@     �H@      �@     �v@      8@      i@      X@      &@      >@      &@      G@     @l@      &@      q@      &@      "@      ?@      <@     �i@      c@      $@      W@     �P@      &@      <@      @     �@@     �f@      &@     �k@      &@       @      =@      8@     `f@      _@      $@     �T@      5@      @      2@      �?      $@      <@      @      :@      @      @      @      @     �D@      >@      @      :@      G@       @      $@      @      7@     `c@      @     �h@      @      @      6@      3@     @a@     �W@      @     �L@      =@               @      @      *@     �E@              I@              �?       @      @      <@      <@              "@      5@               @      @      *@     �E@             �F@              �?       @      @      <@      9@              "@       @                                                      @                                              @                     �N@      .@      "@      @      0@     `n@      .@     �{@       @      �?     �A@      5@     Ps@     �j@      ,@     @[@      :@      &@      @      @      @     �\@      @      d@      �?              "@       @     �d@     �O@      @      H@      :@      @      @      @      @      Y@       @      c@                      "@       @     �c@      O@       @     �F@              @                              ,@       @      @      �?                              @      �?      @      @     �A@      @      @      @      (@      `@      &@     �q@      �?      �?      :@      *@      b@     �b@      "@     �N@     �A@      @      @      @      (@     �[@      @     �k@              �?      4@      *@      ^@      a@       @      J@                                              2@      @     �N@      �?              @              8@      (@      �?      "@     �E@      @      .@       @      7@     �h@      @     �y@      @      @      (@      @     `o@     �^@       @      J@     �B@      @      .@      �?      2@     �b@      @     �s@      @      @      @      @     `k@      Y@       @     �F@      8@       @      $@              *@     �P@      @     �Y@       @       @      @       @     @T@     �F@      �?      :@                                      �?                                               @                      @              @      8@       @      $@              (@     �P@      @     �Y@       @       @       @       @     @T@      E@      �?      4@      *@       @      @      �?      @     @T@             �j@      �?      �?      @      @     @a@     �K@      �?      3@      &@       @      @      �?      @      Q@             `h@      �?      �?      @      @      _@     �J@      �?      3@       @                                      *@              1@                                      ,@       @                      @      �?              �?      @      I@       @     �W@       @              @              @@      7@              @      �?      �?              �?      @      9@       @     �D@                      @              .@      *@              @      �?                      �?      @      1@       @      6@                      @              @       @              @              �?                               @              3@                                       @      &@              @      @                                      9@             �J@       @               @              1@      $@              �?      @                                      @              2@                       @              @      @                       @                                      6@             �A@       @                              (@      @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�8�mhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �0@Eby�1��?�	           ��@                           @ڦ�^�?�            `j@                           @	խ�9�?S            �a@                           �?��*;�?H             ^@������������������������       ��Z�����?*             S@������������������������       ��Ra����?             F@������������������������       �d�
��?             6@                            �?M���3��?.            @Q@	       
                    @�qǱ�?!             H@������������������������       �3�R�f�?             3@������������������������       �(��&y��?             =@                           �?�E�_���?             5@������������������������       ��q-��?             *@������������������������       �      �?              @                          �>@��Vۤo�?)	           �@                            @�5���?�           ��@                            �?�5��5��?H           �@������������������������       �#�t��?�           ��@������������������������       �5��F�?�           @�@                           �?b���R�?u           ��@������������������������       �_D��o�?           �z@������������������������       ��f��.�?a           @�@                           @r�[wGO�?l            �e@                          @@@���l5d�?c            �c@������������������������       �8��d�`�?;             Y@������������������������       ��t�� �?(            �M@������������������������       �ƒ_,���?	             .@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        g@      C@     �E@      ?@     �Y@     h�@      A@     ��@      *@      @      S@      G@     (�@     H�@      0@      o@      @      �?      �?      @      @     �F@      @      ?@              �?      @      @      A@     �B@              ;@       @      �?              @      @      B@      @      6@              �?      @      @      7@      2@              0@       @      �?              @       @      =@      @      4@              �?      @      @      5@      &@              0@       @      �?              @      �?      5@      @      "@                       @      @      .@      $@              @                                      �?       @       @      &@              �?       @              @      �?              (@                                      @      @               @                                       @      @                      @              �?       @              "@              "@                       @              &@      3@              &@      @              �?                      @              "@                       @              $@      "@              "@       @                                      @                                                      @       @               @      �?              �?                      �?              "@                       @              @      �?              @       @                       @              @                                                      �?      $@               @       @                                      �?                                                      �?      @               @                               @              @                                                              @                      f@     �B@      E@      9@     @X@      �@      <@      �@      *@      @     �Q@     �E@     �@      �@      0@     �k@      e@     �B@      E@      9@      X@     P�@      9@     �@      &@      @     �P@      D@     Ѕ@     ��@      ,@      k@     @`@      <@      ?@      4@      S@      z@      3@     �@      $@      @     �O@      A@     ~@      y@      *@     �f@     �U@      5@      3@      3@     �L@     �s@      &@     8�@      @              D@      8@     �w@     �p@      &@     �]@      F@      @      (@      �?      3@     �X@       @     �^@      @      @      7@      $@     �X@     �`@       @     �N@     �C@      "@      &@      @      4@      e@      @     t@      �?              @      @      k@     �`@      �?     �B@      9@      @      @      @      .@      U@      @      Z@                       @       @     @U@     �Q@              6@      ,@      @      @       @      @      U@      @      k@      �?               @      @     �`@      O@      �?      .@       @                              �?      6@      @     @Q@       @              @      @     �D@      .@       @      @       @                              �?      6@      @      P@       @              @      �?     �@@      .@       @      @       @                                      .@      @      B@      �?              @      �?      <@      @      �?      @      @                              �?      @              <@      �?                              @      "@      �?      �?                                                              @                               @       @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���FhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?^���W�?�	           ��@       	                     @�Ȭl�?1           ��@                          �7@���z6Y�?           ��@                            �?܍'x�r�?L           ��@������������������������       �:��#+�?�           ��@������������������������       ��־a��?�            �k@                           �?��ܕ�?�            �s@������������������������       ��}3���?C            �Z@������������������������       ��%�2��?}            �i@
                           @��;�,�?%            }@                          �5@w�Xj��?�             n@������������������������       ��5YYP�?S             `@������������������������       ���S�r��?I             \@                           @Rs�O�1�?�             l@������������������������       ���G�A�?.            �S@������������������������       ���f1F��?[            `b@                          �<@�Zȝ��?k           �@                           @X�-���?�           8�@                           �?�{l�v]�?2            �@������������������������       �����,�?�           `�@������������������������       �0���?�             k@                            @Ƕ�����?�           (�@������������������������       �:m��O�?�           ��@������������������������       �#P�! T�?�            ps@                            @�	��
�?|            �g@                           @��#a�?R            �_@������������������������       �j�V���?:             V@������������������������       �����6��?             C@                           @     ��?*             P@������������������������       �rmhc^Y�?#            �I@������������������������       ���WV��?             *@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@     �K@     �F@      4@     �Y@     p�@      @@     |�@      .@      "@     �R@      L@     ��@      }@      4@     �p@     �U@      >@      :@      (@     �K@     ps@      1@      {@      "@      @     �@@      =@     Pr@     �l@      &@     �b@      N@      1@      5@      (@     �F@     @k@      ,@     �r@       @      @      :@      ;@     �i@      e@      &@      _@      G@      .@      3@      @      B@      f@      (@     �j@      @      �?      2@      ;@     �`@     �a@      &@      U@     �C@      @      .@      @      9@     �a@      &@     `f@      �?      �?      0@      1@      [@     �W@      @      O@      @      "@      @      �?      &@      B@      �?      B@      @               @      $@      9@     �F@      @      6@      ,@       @       @      @      "@     �D@       @     �T@       @      @       @             @R@      =@              D@               @       @      @      @      .@              ?@                      @              *@      @              2@      ,@                              @      :@       @     �I@       @      @      �?              N@      6@              6@      :@      *@      @              $@     @W@      @     �`@      �?      �?      @       @     �U@     �M@              8@      (@      @      @              @      D@      @     �R@      �?              @      �?     �L@      5@              ,@      @      @       @              @     �@@      �?     �E@                      @              3@      @              @      @              @                      @       @      @@      �?                      �?      C@      ,@              @      ,@      "@                      @     �J@              N@              �?       @      �?      >@      C@              $@      @                               @      <@              4@                                      @      .@              @      "@      "@                      @      9@              D@              �?       @      �?      9@      7@              @     �Z@      9@      3@       @     �G@     ps@      .@     x�@      @      @     �D@      ;@     �|@     �m@      "@      ^@      Z@      9@      3@       @     �F@     �q@      .@     �@       @      �?     �@@      7@      z@     �l@       @      \@      O@      $@      "@      @      6@      ^@      @     `s@                      @      @      j@      T@              L@     �H@      �?       @      @      1@     �V@      @     �n@                      @      @     �b@      O@              C@      *@      "@      �?              @      >@             �O@                      �?              M@      2@              2@      E@      .@      $@       @      7@     @d@      &@     �v@       @      �?      ;@      0@     @j@     �b@       @      L@     �A@       @       @       @      1@     �Z@      "@     �m@      �?      �?      :@      &@      c@     @]@      @     �H@      @      @       @              @      L@       @      _@      �?              �?      @      M@     �@@       @      @       @                               @      =@             �S@      @      @       @      @     �E@       @      �?       @       @                                      3@              F@       @               @      @      >@       @      �?       @      �?                                      .@             �@@                              @      3@       @      �?       @      �?                                      @              &@       @               @      �?      &@                                                               @      $@              A@       @      @                      *@                                                               @      @              ;@              @                      *@                                                                      @              @       @                                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ<_hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @D�3 �k�?�	           ��@       	                     �?������?�           L�@                            �?=�8��?@           �@                          �<@[��s���?�           �@������������������������       ��l���	�?\           8�@������������������������       �*J���V�?;            �V@                           @�-�}��?�           Ȑ@������������������������       ��Ѩ�E�?h           8�@������������������������       �4�0���?A            �Z@
                           �?������?�           ��@                           @���Jʸ�?�             n@������������������������       �֔5eMY�?f            �e@������������������������       �4����?.            @Q@                          �0@��4|k�?           |@������������������������       ��9����?            �@@������������������������       ���B��C�?            z@                           �?�b�)��?�           ��@                           @S3��+�?-           �{@                           @���.c�?�            �u@������������������������       ���q��p�?�            @k@������������������������       ���x
��?P            ``@                           @��m��?I            @X@������������������������       ��m����?-             M@������������������������       �~C_j��?            �C@                          �2@k�N�y�?�           (�@                           @zj�ì?�?`            �a@������������������������       ���n�)��?Y            @`@������������������������       �Y�����?             &@                          �8@F,��T�?'           �}@������������������������       ����h/��?�            @s@������������������������       �i�uZ���?k            �d@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @j@      .@     �F@      9@      ]@     H�@      ?@     ȑ@      >@      @      R@     �P@      �@     @~@      3@     �m@     `d@      &@      C@      8@     @W@     �}@      8@     `�@      8@      @     �P@     �H@     Ȁ@     Pw@      3@      i@     @_@       @      :@      2@     �I@     x@      0@     ��@      2@      �?      H@      A@     p{@     �o@      ,@      `@      L@      @      @       @      3@     �i@      @     0u@      "@              0@      *@     `l@     �]@      @     �J@      K@      @      @       @      1@      h@      @     @r@       @              0@      (@     @j@     �\@      @     �J@       @                               @      .@      �?     �G@      �?                      �?      1@      @                     @Q@      @      3@      $@      @@     @f@      "@     @p@      "@      �?      @@      5@     �j@     �`@      @     �R@      Q@      @      3@      $@      ?@     �d@      @     �k@      "@      �?      ?@      2@     �g@     �]@      @     �P@      �?                              �?      ,@       @     �B@                      �?      @      8@      0@               @      C@      @      (@      @      E@     @W@       @     �b@      @      @      3@      .@     �X@     �]@      @     @R@      3@       @      @      @      6@      6@       @     �C@       @      �?      @      @     �A@     �K@      �?      8@      &@       @              @      .@      .@       @      @@       @              @      @      3@      F@      �?      3@       @              @      �?      @      @              @              �?              �?      0@      &@              @      3@      �?      @       @      4@     �Q@      @     �[@      @      @      0@      $@     �O@      P@      @     �H@      �?                       @      �?      &@      �?      �?               @      �?              @      @      �?              2@      �?      @              3@      N@      @     @[@      @      �?      .@      $@     �L@      M@      @     �H@     �G@      @      @      �?      7@     `e@      @     `x@      @       @      @      1@     �l@     �[@             �B@      :@      @      @              0@     @T@      @     �_@      @      �?      @      "@     �W@     �M@              ,@      8@      @      @              ,@     @Q@       @      W@      @      �?       @      "@     �P@      J@              @      0@              @              (@      I@       @      H@      �?               @      @     �G@      <@              @       @      @      �?               @      3@              F@       @      �?              @      4@      8@              @       @               @               @      (@       @      A@                      �?              <@      @              @       @               @              �?       @              0@                      �?              3@      @              @                                      �?      @       @      2@                                      "@      �?              @      5@      �?      �?      �?      @     �V@      @     �p@      @      �?       @       @      a@      J@              7@       @              �?              �?      *@              K@                                      G@      &@              @       @              �?              �?      @             �J@                                      E@      &@              @                                              @              �?                                      @                              *@      �?              �?      @     @S@      @     @j@      @      �?       @       @     �V@     �D@              0@      $@      �?              �?              K@      @     @b@      @               @      @     �H@      4@              (@      @                              @      7@              P@              �?              �?     �D@      5@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�@yhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �7@�����?�	           ��@       	                    �?��6���?�           ��@                          �0@������?           �@                           @cT!)��?G            �\@������������������������       �AA�?4             U@������������������������       ��>�>�?             >@                            @X󳶣��?�           P�@������������������������       ��������?           ��@������������������������       ��%��n�?�            �s@
                          �0@j�
%�<�?�           �@                           �?�Ѻ��E�?@             [@������������������������       �(>gj�p�?             ;@������������������������       �x�ĩa�?2            @T@                          �5@����.�?�           T�@������������������������       �,��s-�?�           ��@������������������������       �R�ǅ���?�            Pr@                          �8@�{-��?�           �@                           �?tS]����?�            �p@                           @���!sL�?8            �T@������������������������       �     ��?,             P@������������������������       �<ݚ�?             2@                           @��2ˋF�?w            �f@������������������������       ���^Y��?j            �d@������������������������       ��F����?             1@                           �?h����?7           Ћ@                           �?���%���?�            �s@������������������������       �����?e            �b@������������������������       �T���b�?r            �d@                           �?'���U�?`           ��@������������������������       �܈���H�?=            �[@������������������������       ��yo}���?#           �|@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      B@      I@      ;@      ^@     �@      9@     D�@      5@      @     �V@      N@     �@      @      2@     �o@      e@      7@      H@      4@     �T@     �}@      4@     ��@      1@      @     �P@      G@     `}@     �w@      1@     @h@     �S@      4@     �@@      @      O@     �k@      0@     �q@      *@      @     �B@      >@      k@     �c@      @     �X@      "@      �?      @      �?       @      $@      @      0@      �?       @      @      @      6@      7@              @      @      �?      @      �?      @      "@      �?      *@      �?       @      @       @      3@      &@              @      @              �?              �?      �?       @      @                              �?      @      (@               @     @Q@      3@      =@      @      K@     �j@      *@     �p@      (@      @     �@@      ;@     @h@     �`@      @     �V@     �H@      *@      3@      @     �F@      d@      $@     `f@      (@       @      :@      :@      `@      X@      @     @S@      4@      @      $@              "@     �I@      @     �V@               @      @      �?     �P@     �B@              ,@     �V@      @      .@      ,@      4@     �o@      @     `{@      @      �?      =@      0@     �o@     `l@      $@      X@       @                                     �A@              1@                      �?      @      7@      2@               @      �?                                      $@                                                      @      @              @      �?                                      9@              1@                      �?      @      0@      (@              @      V@      @      .@      ,@      4@      k@      @     Pz@      @      �?      <@      (@     �l@      j@      $@      V@     @P@      �?      *@      $@      ,@     �d@      @     Pu@       @              5@       @      g@     �c@      @     �S@      7@       @       @      @      @     �I@              T@       @      �?      @      @      G@     �J@      @      "@     �K@      *@       @      @      C@      i@      @     �w@      @              8@      ,@     �m@     @\@      �?     �M@      "@       @      �?      �?      @     �C@      @     @\@                      @      @     �I@      0@              (@      @                      �?      @      $@              7@                      @              4@      @              @      @                      �?      @       @              2@                      @              1@      @               @      @                                       @              @                                      @                      @       @       @      �?               @      =@      @     �V@                      @      @      ?@      "@              @       @       @                      �?      =@      @      U@                      @      @      8@      "@              @                      �?              �?                      @                                      @                       @      G@      &@      �?      @      ?@     @d@       @     �p@      @              1@      &@     @g@     @X@      �?     �G@      ;@      @      �?      @      ,@     �L@       @     @T@      �?              @      �?     �I@      E@              9@      2@      @               @       @      6@             �D@                      @              4@      (@              0@      "@      �?      �?      �?      @     �A@       @      D@      �?                      �?      ?@      >@              "@      3@      @              @      1@     @Z@             `g@      @              &@      $@     �`@     �K@      �?      6@      @       @                      @      6@              =@                              �?      3@      4@              @      ,@      @              @      $@     �T@             �c@      @              &@      "@      ]@     �A@      �?      0@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���shG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@/w��Wu�?�	           ��@       	                    �?�U3��?�           <�@                           �?1�v\*�?�           4�@                            �?�?ӈ�7�?}            `g@������������������������       ��.�?��?'             N@������������������������       ��M�F�~�?V            �_@                          �1@�{f�>�?\           H�@������������������������       ��C�1 �?�            �q@������������������������       ��JӞ��?�           ��@
                           @����V��?�           D�@                            @ޢ��ɵ�?	           ��@������������������������       ��j��@�?m           ��@������������������������       ��"���?�            `n@                           �?��Ze���?�           ��@������������������������       ��q��U�?g             e@������������������������       ��:��#��?T           ��@                           @ؿv�"��?
           �z@                           �?|�Pk��?s             i@                           �?��d�7��?             A@������������������������       �3�R�f�?             3@������������������������       ��K~���?             .@                          @@@��N���?`            �d@������������������������       �]ǿ��S�?N            �`@������������������������       ���3���?             ?@                            @����u�?�            `l@                          @@@^*80��?f            `c@������������������������       ��K�H"�?W            �`@������������������������       ��4_�g�?             6@                           @
�%����?1             R@������������������������       �v�"���?             5@������������������������       �R�3�t�?#            �I@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @l@     �B@     �E@      3@     @V@     ��@     �@@     �@      1@      @     �U@      P@     ��@     �@      5@      o@     `i@      =@     �C@      1@     �S@      �@      >@     ��@      ,@      @     @Q@     �N@     H�@     @~@      2@     �l@     �W@      (@      9@      "@      I@     �r@      4@      v@      "@      @      ?@     �A@     �q@     �g@      $@      ^@       @      �?      @              @      ;@      �?      M@       @              @      @      B@      6@              2@      �?      �?                              @      �?      7@                       @      @      *@       @              @      @              @              @      8@             �A@       @              @              7@      ,@              *@     �U@      &@      6@      "@     �G@     @q@      3@     �r@      @      @      :@      @@     �n@      e@      $@     �Y@      5@      @       @              0@     �F@      @      C@              �?       @      "@     �J@     �C@      @      =@     @P@      @      ,@      "@      ?@     �l@      (@      p@      @      @      2@      7@      h@     @`@      @     @R@     @[@      1@      ,@       @      =@     s@      $@     ��@      @       @      C@      :@     �t@     Pr@       @      [@     �O@      @      @       @      "@     @a@      �?     Pp@                      $@      *@     `e@     @V@              I@     �L@      @      @              "@     �W@      �?     �e@                      @      *@     @Z@     �P@              D@      @              �?       @             �E@             @V@                      @             �P@      7@              $@      G@      (@      "@      @      4@     �d@      "@     w@      @       @      <@      *@     �d@     �i@       @      M@      ,@              @              "@      2@      �?     �G@                       @              6@     �D@      @      @      @@      (@      @      @      &@     �b@       @      t@      @       @      :@      *@     �a@     `d@      @      J@      7@       @      @       @      $@      L@      @     @e@      @      �?      2@      @      S@      ;@      @      4@      (@       @      @       @      @      6@      @     �O@       @      �?      $@      @     �D@      &@       @      $@      @      @                              "@              �?                      @       @      @      �?               @                                               @              �?                      �?       @      @      �?              �?      @      @                              �?                                      @              �?                      �?      "@      @      @       @      @      *@      @      O@       @      �?      @      �?     �A@      $@       @       @      @      @      @       @      @      *@      @     �E@                      @      �?      >@      $@               @       @                                                      3@       @      �?                      @               @              &@                              @      A@             �Z@      �?               @             �A@      0@      �?      $@      @                              @      2@             @Q@                       @              :@      ,@      �?      $@      @                              @      0@             �O@                       @              5@      @      �?      $@      �?                                       @              @                                      @       @                      @                              �?      0@              C@      �?                              "@       @                      �?                                      @              (@                                              �?                      @                              �?      "@              :@      �?                              "@      �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @Oni̹y�?�	           ��@       	                    �?������?�           ��@                           @���b�V�?�           �@                           �?��-�%�?�           �@������������������������       ��i&�<�?           |@������������������������       ��wt��?�            v@                          �;@�_UY�o�?           �y@������������������������       ���a�`�?�            @v@������������������������       �eIG��S�?             K@
                            �?�R��s�?�           ��@                           @mR\o�?�           Ē@������������������������       ��j��8&�?9           ��@������������������������       ����Kh�?�             r@                           @m�c��x�?�            0w@������������������������       �}�s���?�            �s@������������������������       �W��_��?$            �K@                           @�$��33�?�           ��@                          �0@������?           @�@                           @V4�ͫ�?             >@������������������������       ����,�?             3@������������������������       �b���i��?             &@                           @{����Z�?�           P�@������������������������       ��Q��'�?<           �}@������������������������       �Z������?�            �r@                          �<@��O��'�?�            t@                          �:@=V���?�            0r@������������������������       ��(��dN�?�             q@������������������������       ����.�?             3@                           �?d��0u��?             >@������������������������       ��IєX�?	             1@������������������������       ��n_Y�K�?             *@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @g@     �C@     �C@      8@     �V@     �@      :@     @�@      .@       @     @U@      P@     ��@     P@      6@     @q@     �`@      <@      ?@      6@     �Q@     @|@      5@     8�@      *@      @     �Q@      K@     H�@     w@      6@      l@     �P@      $@      6@      (@     �I@     �k@      $@     `q@      @      @      >@      <@      j@      c@      @     �Y@      L@      @      .@       @     �F@     �a@      �?      i@      @      @      1@      2@     �a@     �W@      �?      J@     �@@      �?       @       @      2@     �V@      �?      [@       @       @      (@      &@     �O@      M@      �?     �@@      7@      @      @              ;@     �I@             @W@       @      @      @      @     @S@      B@              3@      &@      @      @      @      @     @T@      "@     @S@       @              *@      $@     @Q@     �M@      @     �I@       @      @      @      @      @     @T@      "@     @P@       @              $@      $@      L@      I@      @     �B@      @                                                      (@                      @              *@      "@              ,@      Q@      2@      "@      $@      4@     �l@      &@     {@      @       @      D@      :@     �u@      k@      0@     �^@     �F@      1@      @      "@      ,@     �g@       @     v@      @              5@      *@     �p@      d@      "@     �T@      E@      ,@      @      @      $@     `b@       @     �o@      @              0@      $@     �i@     �`@      @     �J@      @      @      �?       @      @      E@             �X@      @              @      @      P@      :@      @      =@      7@      �?      @      �?      @     �D@      @      T@               @      3@      *@     �R@      L@      @      D@      3@      �?      @      �?      @      B@      @      O@               @      2@      *@      M@      K@      @      ?@      @                                      @              2@                      �?              0@       @              "@     �I@      &@       @       @      4@     �g@      @     �x@       @      �?      .@      $@     �m@     �`@             �I@     �F@       @      @      �?      0@     �a@      @     `p@       @      �?      @      "@     �e@     �W@             �B@       @                              �?      @              @                       @      �?      @      &@               @                                              �?              @                       @      �?      @      @              �?       @                              �?       @                                                              @              �?     �E@       @      @      �?      .@     `a@      @     0p@       @      �?      @       @     @e@     �T@             �A@      7@              @      �?      $@      T@      @     �c@       @      �?      @      @     �]@      G@              8@      4@       @      �?              @     �M@       @     @Y@                              @      J@     �B@              &@      @      @      @      �?      @     �G@             ``@                      "@      �?      P@      C@              ,@      @      @      @      �?      @     �F@             �[@                      "@      �?      M@     �B@              ,@      @       @              �?      @      B@              [@                      "@      �?     �L@      B@              (@              �?      @                      "@               @                                      �?      �?               @                                               @              5@                                      @      �?                                                                              (@                                      @      �?                                                               @              "@                                       @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�rWhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?fYM����?�	           ��@       	                   �:@�,e�%�?D           ܚ@                           @{<	�,�?�           @�@                           �?]���s�?�           x�@������������������������       �P,E���?�            �h@������������������������       ��L}5��?           �|@                           @=��G'�?           �@������������������������       ����G��?s           ��@������������������������       ��	]�!��?�            @m@
                           �?��� �?�            �l@                           �?�<q,���?#             M@������������������������       ��{�ۨ�?            �A@������������������������       ��o����?             7@                            �?�o�p���?u            �e@������������������������       �t��*f��?             E@������������������������       ���g�0��?X            ``@                           @h#�LD��?j           $�@                           �?T1�κ�?C           ��@                            �?Lj�'Z��?e            �d@������������������������       �0�S�v�?"            �I@������������������������       �,��i�?C            @\@                           �?��z\�g�?�           ��@������������������������       �y!'�/�?q           ��@������������������������       ���Q���?m             d@                          �<@�����?'           ��@                            @�2�L�?�           ��@������������������������       �зs`G��?           ؉@������������������������       �6j �N�?�            �r@                          �=@������?W            �b@������������������������       ��Q����?             D@������������������������       ��9S˅��?@             [@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `h@      =@      @@      >@     @\@     ��@      6@     ̐@      1@      @     �S@     �O@     ��@     x�@      6@     �p@     �W@      2@      :@      0@     @P@     �s@      *@     `x@      &@      @      ;@      B@     pt@     �m@      "@     �`@      U@      (@      6@      *@      L@      r@      (@     Ps@      "@      @      3@      A@     �q@      k@       @     �\@      H@      @      &@      "@      2@     �`@      @     �`@       @      �?      @      @     @Z@     @\@      �?     �M@      0@      �?              @      "@     �A@      �?      E@       @              @      �?     �F@      7@              0@      @@      @      &@      @      "@     �X@      @     @W@              �?       @      @      N@     �V@      �?     �E@      B@       @      &@      @      C@     �c@      @     �e@      @       @      ,@      =@     �f@      Z@      @      L@      7@       @      &@      �?      8@     @]@      @     @]@      @       @      &@      9@     �a@      O@      @      C@      *@                      @      ,@     �C@       @     �L@                      @      @     �C@      E@              2@      &@      @      @      @      "@      8@      �?     @T@       @               @       @      E@      4@      �?      1@      @                      @              @              1@                      @       @      0@       @              @                              @               @              ,@                      @       @      @                      @      @                                       @              @                                      (@       @              �?       @      @      @              "@      4@      �?      P@       @               @              :@      2@      �?      (@                                      @      @      �?      ;@                      �?              �?       @              �?       @      @      @              @      ,@             �B@       @              �?              9@      0@      �?      &@      Y@      &@      @      ,@      H@     pw@      "@     h�@      @       @     �I@      ;@     �z@      r@      *@     �`@     �L@       @       @       @      7@      a@       @      r@      �?      �?      .@      "@     `j@     @X@      �?     �N@       @      �?       @       @      @      ;@              B@                      @             �C@      4@              4@      @                              @      .@               @                                      &@      @              @      @      �?       @       @      @      (@              <@                      @              <@      0@              .@     �H@      �?              @      1@     @[@       @     �o@      �?      �?      (@      "@     �e@     @S@      �?     �D@     �C@      �?              @      &@      U@      �?      j@      �?      �?       @       @     �`@     �P@      �?      8@      $@                              @      9@      �?      G@                      @      �?      D@      $@              1@     �E@      "@      @      @      9@     �m@      @     �x@      @      �?      B@      2@     �j@      h@      (@     �Q@      E@      "@      @      @      9@     �i@      @     �t@      �?      �?     �@@      2@     @g@      g@      (@      Q@      C@       @      @      @      3@     �b@      @     �j@      �?      �?      @@      (@     �^@     @b@      $@     �M@      @      �?      �?              @     �K@      �?      ]@                      �?      @     �O@      C@       @      "@      �?                                      A@             �P@      @              @              <@      "@              @                                              *@              3@                       @               @      @                      �?                                      5@             �G@      @              �?              :@      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���1hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �<@�$j�!m�?�	           ��@       	                    �?"�`���?�           :�@                          �1@�����?           |�@                           @�f����?�            �r@������������������������       �ÇՊ~��?�            �l@������������������������       �5�w.�?)            �R@                           @��N��?A           ��@������������������������       ���K���?           8�@������������������������       �{���9��?=            �X@
                           !@�������?�           ��@                           @��0����?�           ��@������������������������       �������?�           �@������������������������       �`�/�VU�?            P�@������������������������       �T�r
^N�?
             ,@                           �?����Mb�?�            �r@                            �?�d:�1�?             �K@                           @ ��$��?            �E@������������������������       ���<b���?             7@������������������������       �H�z�G�?             4@������������������������       �r�q��?             (@                           �?$�>��?�            �n@                           @|�!��?>            @V@������������������������       �:m��:�?*             N@������������������������       ���`���?             =@                          �?@��|�l�?j            �c@������������������������       �w/�Ln��?B            �Y@������������������������       �JS9�I�?(            �J@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `j@      =@      E@      :@     �V@     �@     �A@     ��@      4@      @     �Q@      K@     ��@      @      0@     �p@      i@      ;@     �D@      :@     �U@     P�@     �@@     ��@      .@      @     �P@     �I@     `�@      ~@      0@     `o@     �Z@      &@      ?@      0@      K@     0q@      1@     �y@      *@      @      ;@      8@     pp@      m@       @     �`@      6@      �?       @      �?      2@     �F@      @     �K@      @       @      @      @     �C@      L@      @      =@      2@              @      �?      ,@     �A@       @      @@      @      �?      @      @      @@     �G@       @      9@      @      �?      @              @      $@      @      7@              �?              @      @      "@       @      @      U@      $@      7@      .@      B@     �l@      &@     �v@      "@       @      4@      2@      l@      f@      @     @Z@     @T@      $@      6@      .@      B@     �k@       @     �t@       @       @      4@      1@     `i@     �d@      @     �U@      @              �?                       @      @      =@      �?                      �?      5@      (@              3@     �W@      0@      $@      $@      @@     pu@      0@     ��@       @       @      D@      ;@     Pz@     �n@       @     @]@     �W@      0@      $@      $@      @@     �t@      0@     ��@       @       @      D@      ;@     @z@     �n@       @     �\@     �J@       @      @      @      .@     �h@      @     v@       @      �?      9@      ,@     `q@      a@      @     �M@     �D@       @      @      @      1@     @a@      &@     �n@              �?      .@      *@     �a@      [@      @      L@                                              "@                                                      �?       @               @      &@       @      �?              @     �L@       @     @^@      @              @      @     �I@      2@              4@      @                                      ,@              2@                       @              @      @              "@      @                                      *@              "@                       @              @      @              "@      @                                      $@               @                                                              @                                              @              @                       @              @      @               @                                              �?              "@                                               @                      @       @      �?              @     �E@       @     �Y@      @               @      @      H@      *@              &@      @       @      �?              @       @              B@       @               @              1@      @              @      @       @      �?              @       @              7@       @               @              &@      @              �?      �?                                                      *@                                      @      @              @       @                               @     �A@       @     �P@      @                      @      ?@      @              @      �?                                      ;@       @      H@      �?                              0@      @              @      �?                               @       @              3@       @                      @      .@      @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ13�ohG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?`tб�j�?�	           ��@       	                   �<@��y�h�?`           ��@                           @�)&�)�?           Ș@                          �3@3�i$�?           t�@������������������������       �F}RE&;�?�           ��@������������������������       ��x��*��?g           (�@                           !@ŕ�(�?             5@������������������������       ���!pc�?             &@������������������������       �R���Q�?             $@
                            �?��-T���?P             _@                           @      �?             @@������������������������       �9����!�?             6@������������������������       ����(\��?             $@                          @@@�H�~Z��?<             W@������������������������       �	~�ϰ�?2            @S@������������������������       �<+	���?
             .@                            @naU���?v           6�@                          �2@?m�1?b�?�           ��@                           @:�Jq���?           �y@������������������������       �0�Z�?�            `m@������������������������       ���s�q��?j            �e@                           @�d@9%�?�           X�@������������������������       �c����%�?�           T�@������������������������       ���4��?T             `@                           �?������?�           `�@                          �1@��4	u�??            @W@������������������������       ��h$��W�?             .@������������������������       ��P1���?8            �S@                           �?��w�R��?P           x�@������������������������       ��)�Y7��?�            �r@������������������������       �d*<��?�            �l@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @h@      A@      @@      <@      Z@     �@      >@     ��@      7@      $@      T@      M@     ��@     0�@      1@     �l@     �X@      5@      9@      $@      O@     �q@      ,@     {@      0@      @     �B@     �@@     Ps@     �m@      (@     �\@     @V@      3@      7@      $@      N@      q@      ,@     x@      .@      @     �@@     �@@     �q@     `k@      &@     �[@      V@      3@      7@      $@     �M@     �p@      (@     x@      .@      @     �@@     �@@     �q@      k@      &@      [@      @@      &@      (@      @      :@     �S@      @     �d@      @      @      7@      .@     �]@     @U@      @     �E@      L@       @      &@      @     �@@      g@      @     �k@      (@       @      $@      2@     �d@     ``@      @     @P@      �?                              �?      $@       @                                               @      @               @                                              @                                                       @       @              �?      �?                              �?      @       @                                                      �?              �?      $@       @       @               @      @              H@      �?              @              7@      4@      �?      @                                      �?      @              5@                                      @      �?              �?                                      �?       @              .@                                      @                      �?                                               @              @                                      �?      �?                      $@       @       @              �?       @              ;@      �?              @              3@      3@      �?      @      @       @       @              �?       @              9@      �?              @              2@      (@      �?      @      @                                                       @                                      �?      @              �?     �W@      *@      @      2@      E@     �v@      0@     ��@      @      @     �E@      9@     �{@     ps@      @     �\@     �R@      (@      @      1@     �C@     �p@      ,@     �{@      @      @     �B@      3@     �s@     `m@      @     �V@      9@               @      @      $@     �S@      �?     @X@                      *@      @      P@      S@      @      >@      .@               @               @     �K@      �?     �J@                       @      @     �G@      ?@      �?      6@      $@                      @       @      7@              F@                      &@      �?      1@     �F@      @       @      I@      (@      @      *@      =@     @g@      *@     �u@      @      @      8@      ,@     �o@     �c@      �?     �N@     �G@      "@      @      &@      <@      f@      "@     �r@      @      @      .@      (@     @l@      a@      �?      M@      @      @               @      �?      $@      @      F@                      "@       @      :@      6@              @      4@      �?      �?      �?      @     @X@       @     �o@       @      �?      @      @      `@      S@              8@      @              �?                      "@      �?     �D@                                      *@      2@              @                                                               @                                      @                      @      @              �?                      "@      �?     �@@                                      $@      2@               @      0@      �?              �?      @      V@      �?     `j@       @      �?      @      @     �\@      M@              2@       @      �?              �?      @      H@      �?     �\@      �?      �?      @      @      L@     �A@              0@       @                                      D@              X@      �?               @             �M@      7@               @�t�bub��
     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ �JhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @W�-����?�	           ��@       	                     @ұ�UF��?�           �@                          �0@����2�?6           ��@                           @�\��$�?h            �e@������������������������       ����Kh�?T             b@������������������������       ��QN���?             ?@                          �2@�z(�g�?�           T�@������������������������       �~2�P%�?]            �@������������������������       �x)"��?q           (�@
                           �?dҍV�$�?�           Ȑ@                          �<@�j�Y�?7           ~@������������������������       �y�c��?           0{@������������������������       ���4c�?             G@                          �5@����%�?j           ��@������������������������       ���n�6�?�            Pt@������������������������       ��9��K�?�            �p@                           @��#ʆA�?�            �s@                            �?O��Ez�?�             r@                           �?<��J���?:            @U@������������������������       �r�q��?              H@������������������������       �0.1�r�?            �B@                           !@��eְ��?�            `i@������������������������       ��_��[��?�            @h@������������������������       �B{	�%��?             "@                            �?b�r���?             >@������������������������       ��8��8��?             (@������������������������       �)O���?             2@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �l@     �D@      F@      >@     �Y@     X�@     �A@     ܐ@      8@      @     �Q@      Q@     ��@     @      3@     �l@      k@     �C@     �B@      =@     �X@     �@      ?@     �@      6@      @     �O@     �P@     ��@     @|@      3@     �j@     @e@      <@      >@      6@     �S@     �{@      8@     h�@      2@      @      L@      N@     �}@     pt@      2@     �e@      &@       @      �?      @      @      A@      @      0@      @               @      $@      :@      @@      �?      *@      &@       @              @      @      =@      @      (@      @               @       @      5@      3@              *@                      �?                      @              @                               @      @      *@      �?             �c@      :@      =@      .@     @R@     �y@      5@     �@      *@      @      H@      I@      |@     pr@      1@     @d@     �J@      @      @       @      (@     �U@      @      b@              �?      (@      .@     �R@     �R@       @     �F@     �Z@      7@      7@      *@     �N@     @t@      ,@     �z@      *@      @      B@     �A@     pw@     �k@      "@     @]@     �G@      &@      @      @      4@     �h@      @     `w@      @      �?      @      @     `k@     @_@      �?     �C@      =@      $@      @      �?      &@     �W@      @     �a@      �?              @      @     �U@      P@      �?      7@      4@      $@      @      �?       @     �W@      @     �_@      �?              @       @      T@      L@              7@      "@                              @      �?              0@                              �?      @       @      �?              2@      �?       @      @      "@     �Y@      @      m@      @      �?       @      @     �`@     �N@              0@      ,@               @      @      @      O@      @      Z@      �?               @      �?     �R@      E@              "@      @      �?                      @     �D@              `@       @      �?              @     �L@      3@              @      &@       @      @      �?      @     �D@      @      ]@       @              @      �?      N@     �F@              1@      &@       @      @      �?      @     �B@      @      Y@       @              @             �M@      D@              ,@      @       @      �?      �?              &@      �?      3@       @              �?              :@      (@              @      �?       @      �?      �?              @              "@       @              �?              (@      "@              @      @                                      @      �?      $@                                      ,@      @              �?      @              @              @      :@      @     @T@                      @             �@@      <@              $@      @              @              @      9@             �S@                      @             �@@      ;@              "@                                              �?      @      @                                              �?              �?                                              @              0@                              �?      �?      @              @                                               @              @                                      �?      �?              �?                                               @              "@                              �?              @               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJi�>2hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �0@ꬱo@��?�	           ��@       	                    @�y)[IP�?            �h@                           �?�-'��?c            �b@                           �?�lXP��?9            @V@������������������������       �@�"s�?             =@������������������������       �[�[��?)             N@                           �?���v��?*             O@������������������������       ��?�߾�?             9@������������������������       ��bp���?            �B@
                           �?�X�%��?            �F@                           @��<,��?             9@������������������������       �UUUUUU�?             (@������������������������       ��q-�?             *@                            �?ffffff�?             4@������������������������       �      �?              @������������������������       ��q�q�?             (@                           �?�?�8���?	           
�@                           @n�$��?�           `�@                           @l���?�           ��@������������������������       ���y��8�?P           Ѐ@������������������������       �'6@���?G           h�@                          @@@KO�����?g           ��@������������������������       �g��r��?_           �@������������������������       �:/����?             ,@                           �?l�n����?           Z�@                          �>@B��Vjo�?�            s@������������������������       ������h�?�            r@������������������������       �     ��?	             0@                           @���	���?Y           �@������������������������       �9��8��?Y            �@������������������������       ��ځ�v`�?            ��@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@      A@     �B@      <@     @Z@     ؄@      D@     ��@       @       @     �T@     �P@     x�@     @      7@     �p@      @      �?      @      @       @     �@@      "@      ?@               @      @      @      ;@     �H@              ,@      @      �?       @      @      @      <@      @      ;@               @      @      @      6@      >@              &@      @      �?       @       @      @      2@      @      *@                              @      *@      9@              �?                       @                       @                                               @      @      *@              �?      @      �?               @      @      $@      @      *@                              �?      $@      (@                       @                      �?      �?      $@      @      ,@               @      @      �?      "@      @              $@       @                              �?       @      @      �?               @       @              @      @              @                              �?               @              *@                       @      �?      @                      @                      @              @      @       @      @                              �?      @      3@              @                      @              @      @       @                                      �?       @      @              @                      @              @      �?                                              �?      �?                      @                                              @       @                                              �?      @                                                              �?              @                                      @      (@                                                                              �?                                      @      @                                                              �?              @                                               @                     �h@     �@@      @@      9@     @X@     Ѓ@      ?@     (�@       @      @     �S@      O@     ��@      |@      7@     �o@     �V@      1@      8@      (@     �M@     pt@      .@     @w@      @      @      ?@     �@@     �r@      i@      "@      `@      K@       @      2@      &@     �I@     �k@      @     �l@      @      �?      7@      6@      j@     �[@      @      V@     �@@      @      *@      @      9@     �X@      @      `@       @              3@      @     �X@     �G@      @     �H@      5@      @      @      @      :@      _@       @     �X@      �?      �?      @      3@     @[@      P@      @     �C@      B@      "@      @      �?       @      Z@       @      b@       @       @       @      &@     �V@     @V@       @     �D@     �@@      "@      @      �?       @     @Y@       @     �a@       @       @       @      &@     �V@     �T@       @     �D@      @                                      @              �?                                              @                     �Z@      0@       @      *@      C@     0s@      0@     ��@      @      @      H@      =@     �|@      o@      ,@      _@      .@              @      �?       @     �@@             @S@                      $@      @     �S@     �D@      @      ?@      .@              @      �?       @      @@             �Q@                      $@      @     �S@     �A@      @      <@                                              �?              @                                              @              @     �V@      0@      @      (@      >@      q@      0@     H�@      @      @      C@      :@     �w@     �i@      &@     @W@     �C@      $@       @       @       @      c@       @     0u@              �?      4@      .@      k@     @Y@      @      A@      J@      @      �?      @      6@     �^@       @     �n@      @       @      2@      &@     `d@     �Z@      @     �M@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�C�WhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@2x��i��?�	           ��@       	                   �0@�cߊ���?�           H�@                           @�1�����?y            �g@                           �?&]^z���?7            �U@������������������������       ����ʀ��?/            @R@������������������������       �����>4�?             ,@                           @�`��[k�?B            @Y@������������������������       �-C��6�?"             I@������������������������       �Y�X��?             �I@
                            @��)���?            Щ@                           @)yF��?�           z�@������������������������       ��F�����?�           ��@������������������������       ��a�n�+�?&           X�@                           @X��D5�?Q           X�@������������������������       �ǆ��q�?            {@������������������������       �T|���?;           �@                           @/��"W�?           Pz@                           �?�����
�?�            `w@                            �?<�4�{�?�            �l@������������������������       �(�:/.��?*            �Q@������������������������       ��p=
�3�?f             d@                            @uk~X���?`             b@������������������������       �	�I�N��?B            @W@������������������������       �(Z���"�?            �I@                          �=@��ȼ��?!            �G@                           �?m��:m�?             >@������������������������       ��(\����?             4@������������������������       �                     $@                          �?@�"�O�|�?             1@������������������������       ������H�?             "@������������������������       �      �?              @�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      A@      B@      4@     �]@     ��@     �C@     X�@      (@      @     �T@      N@     h�@     �~@      3@     �p@     @f@      =@      @@      4@     �[@      �@      C@     H�@      $@      @     �S@      M@     ؄@     �|@      2@     �m@      @      �?      �?      �?       @      A@       @     �@@              �?      �?      @      ?@      E@              4@       @      �?      �?      �?      @      4@       @      1@                      �?      @      &@      2@               @              �?      �?      �?      @      0@       @      &@                      �?      @      "@      2@               @       @                                      @              @                                       @                              @                              �?      ,@              0@              �?              @      4@      8@              2@      @                                      @               @              �?              �?      $@      @              ,@                                      �?      @               @                               @      $@      3@              @     �e@      <@      ?@      3@     �Y@     �@      B@     @�@      $@      @     @S@     �I@     ��@      z@      2@     `k@      a@      4@      6@      ,@      T@     z@      =@     �@      "@      @     �P@      E@     �{@     �s@      1@      f@     @R@      @      *@       @      E@     �f@      (@     Pq@      @      @      3@      4@     �k@     �Z@      @     �R@      P@      .@      "@      @      C@     �m@      1@     �r@      @       @     �G@      6@     �k@     �i@      &@     �Y@     �A@       @      "@      @      6@      d@      @     �t@      �?              &@      "@      h@      Z@      �?     �E@      3@      @      "@      @      @     �M@      @      a@                       @       @     �\@      H@              7@      0@      @               @      1@     �Y@      @     `h@      �?              @      @     @S@      L@      �?      4@      3@      @      @              "@     �M@      �?     �e@       @      �?      @       @     �T@      A@      �?      9@      3@      @      @              "@      K@      �?     `a@       @      �?      @      �?     �S@      ?@      �?      9@      $@      @       @              @     �A@      �?      U@              �?      @      �?      B@      8@      �?      5@       @                              �?      @              A@                                      @      "@              &@       @      @       @              @      =@      �?      I@              �?      @      �?      =@      .@      �?      $@      "@               @              @      3@             �K@       @              �?              E@      @              @      "@                              �?      1@              ?@      �?              �?              9@      @              @                       @               @       @              8@      �?                              1@       @              �?                                              @              A@                              �?      @      @                                                              @              4@                                       @      @                                                              @              $@                                       @      @                                                                              $@                                                                                                                              ,@                              �?       @                                                                                       @                                      �?                                                                                      @                              �?      �?                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJSulMhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B(                             !@�	�̇�?�	           ��@       	                     @��GT���?�	           X�@                           �?�<�`���?�           T�@                           @a���tM�?           Ȓ@������������������������       ���)�[�?�           h�@������������������������       ��������?9             V@                            �?��g(���?�           ��@������������������������       ��<@~���?�           �@������������������������       ��|�N�?�            Pw@
                           �?�c�[)�?�           �@                          �;@(����"�?C           �@������������������������       �m̖C�?            |@������������������������       ���F9���?'            �O@                           @p
�dx1�?�           �@������������������������       ��/>��?�            @w@������������������������       �[?,��?�            �p@                          �8@ �^�@��?             =@������������������������       �x�5?,R�?
             2@������������������������       �b���i��?             &@�t�bh�h4h7K ��h9��R�(KKKK��h��B�	        j@     �@@      C@      >@     �Y@     @�@     �@@     |�@      9@      @     �S@      O@     8�@     p@      3@     �p@      j@     �@@      C@      >@     @Y@     ��@      <@     t�@      9@      @     �S@      O@     (�@     @      3@     `p@      c@      8@      =@      6@     �T@     �{@      9@     X�@      1@      @      P@     �J@     P~@     `x@      0@     `j@     @S@      ,@      5@      @     �G@      l@      &@     �q@      (@      @      1@      <@      g@     �d@      @     �Z@      S@      ,@      .@      @      G@     �j@      &@     �o@      (@      @      1@      <@     �d@     @c@      @      W@      �?              @              �?      &@              ;@                                      1@      &@              ,@     �R@      $@       @      .@     �A@      k@      ,@      {@      @             �G@      9@     �r@      l@      *@     @Z@     �H@      @      @      *@      0@     �e@      $@     �v@      @              7@      ,@      o@     �c@       @     �O@      :@      @      @       @      3@      E@      @      Q@       @              8@      &@     �J@     �P@      @      E@     �L@      "@      "@       @      3@     �h@      @      y@       @      �?      ,@      "@      p@     �Z@      @     �I@      >@      @      @       @      ,@      W@      �?     �b@      @              &@      @     �\@      J@       @      8@      8@      @      @       @      *@     �U@      �?      ^@      @              &@      @      Z@      G@              4@      @                              �?      @              <@                                      &@      @       @      @      ;@      @       @      @      @     �Z@       @     �o@      @      �?      @      @     �a@     �K@      �?      ;@      4@      �?      �?      @      @      C@              c@       @      �?      �?       @     �X@      8@              5@      @       @      �?              �?      Q@       @     �Y@      �?               @      @      E@      ?@      �?      @                                       @      "@      @       @                                       @      @              @                                       @       @      @                                                      �?               @                                              �?               @                                       @      @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�{��8��?�	           ��@       	                    @H��bf�?�           V�@                           �?��x3�?*           f�@                           �?����ΰ�?�           ��@������������������������       ����	`��?�            ps@������������������������       �� ��?           ��@                           �?��V\��?Z           �@������������������������       ��/��U2�?E           ��@������������������������       ��1o���?           ��@
                           @�s�-���?�             o@                          �:@/Fy���?x            �h@������������������������       ��p�]�?\            @c@������������������������       ��ˠT�?             F@                            �?t$���~�?             I@������������������������       �����K�?
             2@������������������������       �     @�?             @@                           @�*�����?�           x�@                           �?�G8�b��?D           �@                           �?��C0�?�             r@������������������������       �|?_���?{            �f@������������������������       ���3S��?I            �Z@                          �2@Dn6mq��?�             k@������������������������       �]t�E�?3             V@������������������������       �     ��?M             `@                          �3@���/��?�            �@                           �?�nג���?w            @h@������������������������       �8	C)��??            @Z@������������������������       ��T&>MJ�?8            @V@                           @���B��?            ~@������������������������       ����P��?^            �c@������������������������       �a
67١�?�            @t@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @k@     �@@     �E@      4@      Y@     p�@      A@     (�@      (@      @      Q@     �V@     `�@     �@      4@     `p@      f@      2@      @@      (@      U@     |@      =@     8�@       @      @     �O@     �T@      ~@     �w@      .@     `k@     @e@      1@      >@      (@     �S@     Pz@      7@     ��@       @      @      M@     �S@     p{@     �u@      .@     �g@     �T@      @      8@      @      G@     �j@      "@     @k@      @      @      =@      F@     �g@      c@      $@      W@      &@      @      *@       @      &@      L@      �?     �L@       @              0@      $@     �C@     �H@       @     �C@      R@      @      &@      @     �A@     �c@       @      d@      @      @      *@      A@     �b@      Z@       @     �J@     �U@      $@      @      @     �@@      j@      ,@     �w@       @      �?      =@     �A@     @o@     �g@      @      X@     �B@      @      @       @      @      T@       @     �d@      �?              @      8@     @Z@     �N@       @     �A@      I@      @      @      @      =@      `@      @     �j@      �?      �?      :@      &@      b@     @`@      @     �N@      @      �?       @              @      <@      @      U@                      @      @     �E@     �@@              ?@      �?               @              �?      4@      @     �R@                      @      @      A@      ;@              9@                       @              �?      0@      @     �F@                      @       @      =@      9@              8@      �?                                      @              >@                              �?      @       @              �?      @      �?                      @       @      �?      "@                                      "@      @              @      @      �?                      @      @                                                                              @      @                                       @      �?      "@                                      "@      @               @     �D@      .@      &@       @      0@     �i@      @     0z@      @       @      @      "@     �p@      `@      @     �E@      0@      @      &@       @      @      P@       @     @g@                      @      �?     @`@     �H@              8@      @              @      @      @      F@      �?     @^@                       @              K@     �A@              (@      �?               @      @              @@      �?     @R@                                      A@      <@              "@      @              @       @      @      (@              H@                       @              4@      @              @      "@      @      @      @      �?      4@      �?     @P@                      @      �?      S@      ,@              (@       @                      @              $@              6@                                     �F@      @              @      @      @      @              �?      $@      �?     �E@                      @      �?      ?@      &@              "@      9@      $@                      &@     �a@      @      m@      @       @               @      a@     �S@      @      3@      *@      @                      @      6@      �?      S@                              @     �B@      4@              &@      *@       @                      @       @      �?      ?@                              @      1@      0@               @               @                              ,@             �F@                              �?      4@      @              @      (@      @                      @     �]@       @     �c@      @       @              @     �X@     �M@      @       @      @                              @      G@              G@                                      >@      3@              @       @      @                             @R@       @     �[@      @       @              @     @Q@      D@      @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�E"VhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�P���?�	           ��@       	                   �1@H3YP���?�           �@                           �?��[��?4           `@                           @�͘DA�?�            �p@������������������������       �s��A�?w             i@������������������������       �lRyӳ�?.            �Q@                            �?�>��W��?�            �l@������������������������       ��in��?i            `e@������������������������       ���Wϊ�?&             N@
                          �=@�g�����?�           �@                            �?���5��?_           �@������������������������       ���[R�W�?           ��@������������������������       �t�Y���?I           H�@                          �@@9,�WT��?[             b@������������������������       ��_,�Œ�?M             ^@������������������������       ���+e��?             9@                           @��(#�#�?�           D�@                           �?��~�?	           ��@                           �?�j:�ٶ�?�            0t@������������������������       �     ��?�             p@������������������������       ��E�6@J�?&            �P@                           @M�s��D�?;           P@������������������������       �������?�            @x@������������������������       �Pql�4�?I            @\@                          �2@|;%dG��?�            �q@                           @R:�&�u�?B            @Y@������������������������       �?�ܵ�?"             I@������������������������       �b�H�/��?             �I@                           @�7V��?~            �f@������������������������       ���1G���?D            �V@������������������������       �UIS�"�?:            @V@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `h@      >@     �E@      3@     �Z@      �@     �D@     |�@      3@      @      Q@     �P@     8�@     �@      6@     `q@     `a@      8@      >@      ,@     @V@     @}@      =@     ��@      0@      @      O@      N@     �~@     @y@      5@      m@     �@@      @      "@      �?      4@      X@      &@     �W@      �?      �?      (@      6@      O@     @U@      @     �E@      1@      @      @              4@      I@      &@     �B@      �?      �?      @      *@     �@@      F@      @      9@      *@      @      @              $@      A@       @      =@                      @      (@      <@      ?@      @      4@      @              �?              $@      0@      @       @      �?      �?      @      �?      @      *@              @      0@       @      @      �?              G@             �L@                      @      "@      =@     �D@       @      2@      *@       @                              ?@             �J@                      �?      @      ;@      8@              .@      @              @      �?              .@              @                      @      @       @      1@       @      @     �Z@      3@      5@      *@     @Q@     @w@      2@     ��@      .@      @      I@      C@     �z@     �s@      ,@     �g@     �Y@      2@      5@      *@     �P@      v@      1@     ��@      *@      @      I@     �@@     �y@     �r@      ,@      f@     �Q@      ,@      ,@      $@      F@     �r@      *@     p}@      @              B@      7@     0t@     �h@      $@      \@      @@      @      @      @      7@      L@      @     @Y@      "@      @      ,@      $@     �U@     �X@      @     @P@      @      �?                       @      4@      �?     �L@       @                      @      5@      5@              (@      @      �?                       @      .@      �?     �K@       @                      @      1@      (@              "@                                              @               @                               @      @      "@              @      L@      @      *@      @      1@      f@      (@     �x@      @      �?      @      @     @k@     �a@      �?      G@      I@      @      (@      @      $@     �`@       @      q@       @      �?      @      @     �d@     �]@      �?      B@      7@       @      @               @      P@       @     �R@       @              �?       @      N@      K@      �?      1@      4@      �?      @               @      I@              O@       @              �?       @     �E@      G@      �?      ,@      @      �?                              ,@       @      *@                                      1@       @              @      ;@      �?      @      @       @     @Q@             �h@              �?       @      @     @Z@      P@              3@      1@      �?      @      @       @     �E@             �d@              �?       @      �?     @U@     �E@              2@      $@                                      :@             �@@                               @      4@      5@              �?      @      @      �?       @      @     �E@      @     �^@      �?              @      �?     �J@      9@              $@       @                       @              &@      @     �F@                      �?              =@      @               @      �?                                      @              4@                                      5@                       @      �?                       @              @      @      9@                      �?               @      @                      @      @      �?              @      @@             @S@      �?               @      �?      8@      4@               @      @      �?                       @      "@             �G@                      �?              *@      $@              @               @      �?              @      7@              >@      �?              �?      �?      &@      $@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @���\��?�	           ��@       	                     �?��| ��?�           �@                           �?��`�%�?�           4�@                           �?���ݡ�?            �|@������������������������       �g�W���?2             Q@������������������������       ��1 .��?�            `x@                           @*kއc��?}           �@������������������������       �ap�&��?           Py@������������������������       ��@���?u            �e@
                            �?`�+h�Y�?Q           ��@                           �?"]s
�?�           ��@������������������������       ����^��?N           ��@������������������������       ����\�?V           ��@                          �;@��џS��?�           0�@������������������������       �[,�~��?�           ��@������������������������       �<�J���?            �I@                           �?0��ďE�?�           D�@                           @��K�lR�?1           �~@                           @H�E7#��?�            Pt@������������������������       �}^���?�            p@������������������������       ��n#،�?)             Q@                           @9���k�?h            �d@������������������������       �EN7W�?X            @a@������������������������       �4և����?             <@                           @���C+�?�           0�@                           �?3�=;���?�            Px@������������������������       �>����?'            �Q@������������������������       �;u�N��?�            �s@                           @zoi^�?�             l@������������������������       �Ȓ�SB�?s            �f@������������������������       �@r��ճ�?             F@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      @@     �I@      7@     �X@     p�@      A@     �@      6@      "@     �M@     �K@     І@     ��@      4@     Pr@     �b@      8@      D@      2@     �T@     P~@      ;@     0�@      3@      @     �H@      E@     �~@     py@      3@     �m@      K@      @      @       @      9@      g@      (@     �r@      @              "@      .@     �i@      b@      @     �M@      <@      �?      @      �?      .@     @T@      @     �^@      @              @      "@      U@     @P@              @@      @                              �?      @      �?      :@                       @      @      1@      @              @      9@      �?      @      �?      ,@      S@      @     @X@      @              @      @     �P@      N@              ;@      :@      @      �?      @      $@      Z@      @     �f@       @              @      @     @^@      T@      @      ;@      2@      �?      �?       @      @     �S@       @      ]@       @               @      @     �W@     �H@      @      8@       @       @              @      @      9@      @      P@                       @              ;@      ?@              @      X@      4@     �A@      $@     �L@     �r@      .@     py@      ,@      @      D@      ;@     �q@     `p@      0@     �f@     �N@      *@      5@      @      ;@     @g@       @     �p@      @              5@      0@      e@      a@      @      ^@      @@      $@      4@       @      4@     �X@      @     @]@      @              &@       @     @U@      M@       @      L@      =@      @      �?       @      @     �U@      �?      c@                      $@       @     �T@     �S@       @      P@     �A@      @      ,@      @      >@     �\@      @      a@       @      @      3@      &@     �]@     �_@      (@      N@      A@      @      ,@      @      >@      Y@      @     �^@       @      @      2@      $@     �[@      _@      @     �L@      �?                                      ,@       @      .@                      �?      �?      @       @      @      @      C@       @      &@      @      1@      i@      @     Pw@      @      @      $@      *@     �m@     �^@      �?      K@      9@      @      @       @      *@     @Y@      @     �`@      �?      �?      @      @     �X@      L@      �?      >@      $@       @      @       @      @     �R@      @     @T@                      @      �?     �S@      A@              3@      $@       @      @              @     �N@      @      M@                       @      �?      Q@      :@              0@                      �?       @       @      ,@              7@                      @              $@       @              @      .@       @                       @      :@      @     �J@      �?      �?              @      4@      6@      �?      &@      ,@       @                       @      5@      @      G@      �?      �?              @      &@      2@      �?      "@      �?                                      @              @                                      "@      @               @      *@      @      @      @      @      Y@             �m@       @       @      @      "@     �a@     �P@              8@       @      @      @      @      @      I@              d@      �?       @      �?      @     @W@     �A@              8@      @                              �?      @              >@                                      ,@      @              (@      @      @      @      @       @     �E@             @`@      �?       @      �?      @     �S@      ?@              (@      @      �?      �?              �?      I@             �S@      �?               @      @      H@      ?@                      @              �?              �?      F@             �N@                              @      E@      5@                              �?                              @              2@      �?               @              @      $@                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ6g� hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx                            �1@��G{\�?�	           ��@       	                    @�H��;�?�           p�@                           �?�����?           `z@                           @B�Z�.w�?�            �l@������������������������       �D��Vl�?y            �g@������������������������       ��w����?            �D@                          �0@r�q�?�             h@������������������������       ��l�l�?*             N@������������������������       �ogH���?Y            �`@
                           �?�(��0�?|             i@������������������������       ��:���?             ;@                           @K�m��?k            �e@������������������������       �zqY���?X            �a@������������������������       ��(�B'�?            �@@                           !@5}��<�?1           ��@                            @�����?$           ��@                           @d^9���?�           ԡ@������������������������       �>	rLm��?E           ��@������������������������       �_B{	�Y�?o            �@                           @C�CV���?p           ��@������������������������       �����=��?            |@������������������������       �w��5�?V           ��@                           @8��d�`�?             9@������������������������       �     ��?             0@������������������������       ��2�tk~�?             "@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      @@      >@      6@     �[@      �@      9@     ̑@      .@      $@      S@      J@     ��@     �~@      5@     @o@     �H@      �?      "@      �?      1@      _@      @      ^@      �?      @      @      .@     �[@     @X@      @     �K@      D@      �?      @      �?      *@     @X@      @     �P@               @      �?      @     �T@     �O@      �?      D@      6@      �?       @      �?      *@      E@       @      @@               @      �?      @      G@     �B@      �?      7@      2@      �?      �?      �?      $@     �A@       @      ;@               @      �?      @      E@      7@      �?      4@      @              �?              @      @              @                                      @      ,@              @      2@              �?                     �K@       @     �A@                               @      B@      :@              1@       @                                      4@              "@                               @      &@      @              "@      0@              �?                     �A@       @      :@                                      9@      3@               @      "@              @              @      ;@      @     �J@      �?      @      @       @      =@      A@       @      .@      @                               @      @       @      "@      �?                               @               @              @              @               @      5@      �?      F@              @      @       @      ;@      A@              .@      @              @               @      (@      �?     �A@                      @       @      4@      @@              ,@                                              "@              "@              @      �?              @       @              �?     `c@      ?@      5@      5@     �W@     @�@      2@     ؏@      ,@      @     �Q@     �B@      �@     �x@      2@     `h@     @c@      ?@      5@      5@     @W@     Ѐ@      .@     ȏ@      ,@      @     �Q@     �B@      �@     �x@      2@     `h@      ^@      8@      1@      2@     �R@      w@      (@     8�@      (@      �?     �M@      A@     �z@     r@      *@     �d@     �Y@      *@      .@      0@     �O@     �q@      @     p~@       @      �?      G@      =@     �r@     �h@       @      `@      2@      &@       @       @      &@      U@       @      d@      @              *@      @     �^@      W@      @      C@      A@      @      @      @      3@      e@      @      w@       @      @      &@      @     @k@     @Z@      @      =@      2@       @      @       @      &@      M@      �?     `c@               @      "@       @     @_@      H@              *@      0@      @              �?       @     �[@       @     �j@       @      �?       @      �?     @W@     �L@      @      0@      �?                              �?      ,@      @       @                                              @                      �?                                      (@                                                              @                                                      �?       @      @       @                                              �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJlt$hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�H�M��?�	           ��@       	                   �>@�(�C��?]           ��@                            @�����?O           Ѐ@                          �:@Z1�ĺ�?�            Pv@������������������������       ������?�            @s@������������������������       ��.P��?            �H@                          �6@���n1�?m            �f@������������������������       �Q������?I            �\@������������������������       ��ˠT�?$            �P@
                          �?@�o����?             7@������������������������       �      �?             (@������������������������       �b���i��?             &@                           �?켨*q�?R           0�@                            �?&��}��?�           Đ@                           @4(�.P�?�            `p@������������������������       �&~�_���?�            �k@������������������������       �̄���?            �D@                            @��&#��?�           X�@������������������������       �ޔ�'$��?Q           ��@������������������������       �d_�r:�?�            @q@                          �6@Hb9�5�?�           Ρ@                            @~|d���?�           0�@������������������������       ���w�%�?�           ؏@������������������������       �s�R�t�?�            y@                           �?F�C�J�?#           ؊@������������������������       �>�����?.            �S@������������������������       �_{S���?�           `�@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@     �A@      F@      ;@      \@     �@     �C@     �@      2@      @      T@     �O@     ��@     `}@      @     p@      >@      @       @      @      1@     �Q@       @     �`@      �?              .@      @     �a@     �S@              J@      =@      @       @      @      1@     @P@       @     �^@      �?              .@      @     @a@      S@              J@      5@      @      @      @      *@      C@              T@      �?              (@      @     @W@      E@              F@      4@      �?      @      @      *@      @@             �R@      �?              &@      �?     �P@      D@              D@      �?       @                              @              @                      �?       @      :@       @              @       @              @              @      ;@       @     �E@                      @       @     �F@      A@               @       @               @              @      .@       @      8@                      @       @      @@      .@               @                      @                      (@              3@                                      *@      3@                      �?                                      @              &@                                      @       @                                                               @               @                                               @                      �?                                      @              @                                      @                              e@      @@      B@      7@     �W@     ��@     �B@     �@      1@      @     @P@      M@     ��@     �x@      @     �i@      O@      @      .@      *@      >@      h@      *@     @p@       @              5@      5@     �l@     �a@      @     �M@      .@               @      @      @      J@      @     �W@      �?               @      @     �F@      2@      �?      "@      .@               @      @      @     �D@      @      S@      �?               @      �?     �E@      .@      �?      @                              �?      �?      &@              2@                              @       @      @               @     �G@      @      *@      @      9@     �a@      @     �d@      @              3@      1@      g@     �^@      @      I@      B@      @      &@      @      7@     @Y@       @      V@      @              *@      ,@     �X@      W@      @      B@      &@       @       @               @     �C@      @     �S@                      @      @     @U@      >@              ,@     �Z@      :@      5@      $@     @P@     `y@      8@     ȅ@      "@      @      F@     �B@     �z@     �o@      @     @b@      T@      ,@      .@       @      E@      o@      *@     0y@       @       @      >@      @@     `n@     @f@       @      [@     �P@      &@      &@      @     �A@     �e@      (@      p@       @       @      :@      <@      e@     ``@       @     �V@      ,@      @      @      @      @     �R@      �?      b@                      @      @     �R@     �G@              2@      :@      (@      @       @      7@     �c@      &@     `r@      @       @      ,@      @     @g@     �R@      �?      C@                              �?              "@      @      F@      @      �?      �?              ,@       @              �?      :@      (@      @      �?      7@     �b@       @     @o@      @      �?      *@      @     �e@      R@      �?     �B@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�;|fhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?)�b�g{�?�	           ��@       	                    �? �h[��?1           ��@                           @Կ�e_�?�             m@                           �?bI5����?m             e@������������������������       ���2���?7            �U@������������������������       �R4���5�?6            �T@                            �?     �?*             P@������������������������       ��G�z��?             D@������������������������       ��8��8��?             8@
                            @���L�?�           ܖ@                           @��_A�?�           ��@������������������������       �8���B�?�           ��@������������������������       �!��wy��?�             w@                           @��ˏ�M�?�            0y@������������������������       �s�����?�            �t@������������������������       �t�@�t�?.            �R@                           @ۍ����?e           R�@                           �?5�@L���?Q           �@                          �3@�p.0��?c             e@������������������������       ������?%            �Q@������������������������       �9*��K��?>            �X@                            @<����?�           ؇@������������������������       �n���d�?U           x�@������������������������       �T$�0��?�            �m@                           @�ۉzp��?           �@                           �?_���?�           h�@������������������������       ��n*ɶ��?�            t@������������������������       �t)e�=��?�            �x@                           @�����?d           ȁ@������������������������       �]���j�?#           �|@������������������������       ��>�x��?A            @[@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `g@      A@     �C@      ;@     �X@     �@     �@@     0�@      3@      @      Q@     �R@     Ȉ@     �@      3@     0p@      [@      .@      >@      *@     �L@     �r@      2@     �z@      (@      @      ?@      ?@     �s@      k@      @     �\@      ,@      �?      @              0@     �@@       @     �S@      @               @      @      A@      4@              0@      (@              @              (@      7@              I@                       @      @      9@      0@              .@      @              @              @      @              @@                      @       @      &@       @              "@       @              �?              @      1@              2@                       @       @      ,@       @              @       @      �?                      @      $@       @      <@      @                              "@      @              �?       @      �?                      @       @       @      ,@      �?                              @       @              �?                                               @              ,@       @                              @       @                     �W@      ,@      :@      *@     �D@     pp@      0@     �u@      "@      @      7@      ;@     �q@     �h@      @     �X@     @P@      &@      5@      $@      @@      h@      (@     �l@      @      @      0@      9@     �i@     `a@      @     @U@     �G@       @      1@      $@      >@     �]@       @      d@      @      @      *@      *@     �a@     �Q@       @      J@      2@      @      @               @     �R@      $@     �Q@      �?              @      (@     �P@     @Q@       @     �@@      =@      @      @      @      "@     �Q@      @      ]@      @      �?      @       @     �S@     �L@      @      *@      ;@      @      @              @     �G@      @     �Y@      @      �?      @       @      Q@      G@      @       @       @               @      @       @      7@      �?      *@                      @              $@      &@              @     �S@      3@      "@      ,@      E@     �u@      .@     �@      @       @     �B@      F@     �}@     �r@      (@      b@     �C@      @      @       @      0@      c@             Pp@                      ,@      *@     �m@     �X@      @     �S@      @      �?              �?      @      6@              B@                      �?      @      E@      2@              <@       @                               @      "@              1@                                      1@       @              5@      @      �?              �?      @      *@              3@                      �?      @      9@      0@              @      @@      @      @      @      &@     ``@              l@                      *@      @     @h@     @T@      @      I@      ;@      @       @      @      $@      Y@             �_@                      (@      @      _@     �P@      @      D@      @              @      @      �?      ?@             �X@                      �?             �Q@      ,@              $@      D@      ,@      @      @      :@      h@      .@     �y@      @       @      7@      ?@     �m@     �h@       @     �P@      9@      @      @       @      .@     �Y@      $@     `n@      @       @      .@      6@      ^@     �Y@      @      E@      4@      @      �?       @      &@      L@      @      U@                      �?      $@      Q@      B@              8@      @               @              @      G@      @     �c@      @       @      ,@      (@      J@     �P@      @      2@      .@      &@      �?      @      &@     �V@      @     `e@      �?               @      "@     �]@      X@      @      9@      *@      @      �?      @       @     �Q@      @     `b@      �?              @      @     �W@     �U@      @      @       @      @                      @      3@              8@                       @      @      8@      $@              2@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�7�fhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @ꑑn�?�	           ��@       	                    @Y|�(���?�           ��@                           �?No�����?�           ��@                           �?۳X;���?9           p�@������������������������       ��,�y���?C            �\@������������������������       �.3z��f�?�           ؈@                           �?ڗ=��\�?�           ��@������������������������       �P`;��?s            @g@������������������������       �_��#�?K           ��@
                           @N`��ҽ�?�            �@                           �?b2U0*��?             I@������������������������       ���:m��?             .@������������������������       �
��-��?            �A@                          �;@>��Ϋ��?�           p�@������������������������       �%� �$?�?�           ��@������������������������       �R����?1             T@                          �=@p?����?�           đ@                           �?�x��p��?�           X�@                           @�(�X ��?,           �|@������������������������       �� ��&�?�             u@������������������������       ���y�{�?K            @^@                          �;@f}T�#��?l           X�@������������������������       �*S$Y1��?V           (�@������������������������       ���)�c{�?             C@                           �?���9^�?6            �V@������������������������       �*D>��?             *@                           �?�G�o,�?0            �S@������������������������       ��m۶m��?             <@������������������������       �rh��|?�?             I@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      9@     �E@      6@     @Z@     8�@      A@     ��@      2@      @     �P@      Q@     `�@      @      6@      m@      e@      2@      A@      0@     �V@     �}@      ;@     P�@      .@      @      L@     �L@     �@     `w@      5@     �h@      b@      ,@      7@      (@      Q@     @v@      ,@     (�@      &@       @     �A@     �D@     x@     �n@      0@     �c@     �P@      $@      3@      @     �C@     `d@       @     �h@      $@       @      0@      8@     �c@      Z@      @     �T@      @      �?      @              @      .@              8@      @              "@      @      3@      @              0@      O@      "@      (@      @      @@     �b@       @     �e@      @       @      @      4@      a@      Y@      @     �P@     �S@      @      @      @      =@      h@      @      t@      �?              3@      1@     �l@     �a@      "@     �R@      ,@      �?              �?      (@      6@             �E@                      �?      @     �B@      <@      @      5@      P@      @      @      @      1@     `e@      @     Pq@      �?              2@      ,@      h@      \@      @     �J@      7@      @      &@      @      6@     �]@      *@     �h@      @       @      5@      0@     @_@     @`@      @     �D@                               @       @       @              =@                      �?      @              $@              �?                                              �?              @                              �?              @                                               @       @      �?              6@                      �?       @              @              �?      7@      @      &@       @      4@      ]@      *@      e@      @       @      4@      *@     @_@      ^@      @      D@      6@      @      &@       @      4@     �Y@      *@      `@      @       @      4@      *@     @\@      [@      @     �C@      �?                                      ,@              D@                                      (@      (@              �?     �K@      @      "@      @      .@     �i@      @     �y@      @      �?      $@      &@     �m@     �^@      �?      A@      G@      @      "@      @      (@     @h@      @     �w@      �?      �?      $@      $@      j@     @^@              >@      9@      @      @              (@     �U@       @      a@      �?      �?       @       @     @X@      O@              .@      6@      @      @              &@      P@       @     @V@      �?      �?       @       @      S@      H@              &@      @      �?      �?              �?      7@             �G@                      @              5@      ,@              @      5@      @       @      @             �Z@      @     �n@                       @       @      \@     �M@              .@      5@      @       @      @             @X@      @      l@                       @       @     �[@      K@              .@                                              $@              6@                                      �?      @                      "@                              @      &@              >@       @                      �?      =@      �?      �?      @      @                              �?      �?               @                                                                      @                               @      $@              6@       @                      �?      =@      �?      �?      @      @                               @      �?              @      �?                      �?      @      �?      �?      @       @                                      "@              .@      �?                              7@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJmc6vhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @9��<|�?�	           ��@       	                     �?�������?�           ޥ@                           @Z���5��?2           ��@                          �0@
O��΀�?j           x�@������������������������       ��q����?#            �J@������������������������       �l)�\�?G           Ќ@                           �?
�4���?�           �@������������������������       �h�Zs>�?,            @������������������������       ��]ޒ���?�           ��@
                          �4@E$Gi��?�           Ȅ@                           �?&7)���?�             u@������������������������       ��b-�I�?             3@������������������������       �X��?��?�            �s@                          �=@���p�F�?�            �t@������������������������       ��s|�f'�?�            Pr@������������������������       ��n����?             B@                          �;@n��)Y��?�           h�@                          �2@��S�%�?n           �@                           @�A� э�?�            q@������������������������       �T���sG�?            �g@������������������������       �dIa�_e�?6            �T@                          �9@��#ט��?�           ��@������������������������       �?���?{           ��@������������������������       �N4̡���?>            �W@                           @���=A�?]             c@                           �?x?I|V��?I            �]@������������������������       ��9J����?              J@������������������������       ��Jr[��?)            �P@                           @��M���?             A@������������������������       �����!p�?             6@������������������������       �      �?             (@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      6@      >@      <@     �[@     �@     �C@     ��@      .@       @      U@     �P@     ؇@     �~@      1@     @o@     �e@      2@      7@      7@     @U@      }@     �@@     p�@      $@      @      P@      N@     X�@     `w@      *@     `j@     �`@      &@      &@      4@     �I@     �w@      ;@     h�@       @      �?      G@      @@     �y@      p@      &@     `b@     @T@       @      @      @      <@      g@      "@     �p@      @              7@      &@     �h@     �U@      �?      P@      �?              �?              @      $@      @      @       @               @              .@      @              @      T@       @      @      @      8@     �e@      @     pp@       @              5@      &@     �f@     �S@      �?      N@     �I@      @      @      ,@      7@      h@      2@      t@      @      �?      7@      5@     @k@     �e@      $@     �T@      9@      @      @      @      ,@      V@      @     �Z@      @      �?      *@      "@     @V@     @T@      @     �G@      :@              �?      "@      "@      Z@      &@      k@      �?              $@      (@      `@     �V@      @      B@      E@      @      (@      @      A@      V@      @      `@       @      @      2@      <@     @[@      ]@       @      P@      .@      @      @      @      0@     �H@              L@              @      $@      4@     �B@     �P@      �?     �G@                      @              �?      �?               @                       @               @                       @      .@      @      @      @      .@      H@              K@              @       @      4@     �A@     �P@      �?     �C@      ;@       @      @              2@     �C@      @     @R@       @       @       @       @      R@     �H@      �?      1@      8@       @      @              2@      @@      @      N@       @       @      @      @     �Q@      G@              *@      @                                      @       @      *@                      �?      �?      �?      @      �?      @      H@      @      @      @      :@     @f@      @     `y@      @       @      4@      @      n@     @]@      @     �C@      E@      @      @      @      4@     �b@      @     �t@       @      �?      4@      @      k@      \@             �A@      $@              @      @       @     �F@       @     �S@                       @       @     �R@      ?@              @      $@               @      @      �?      ?@             �F@                      @       @     �O@      5@              @                      �?              @      ,@       @      A@                      @              &@      $@              �?      @@      @      @      �?      (@     �Z@      @      p@       @      �?      (@      @     �a@     @T@              <@      ;@      �?       @      �?      (@     �W@      @     `l@       @      �?      (@      @     @\@      Q@              8@      @      @      �?                      &@              =@                                      =@      *@              @      @              �?              @      ;@             �Q@      @      �?                      8@      @      @      @      @              �?              @      .@              J@      @      �?                      8@      @      @      �?      @              �?              @      @              .@      @                              &@      @      @      �?                                      @      &@             �B@              �?                      *@      �?                                                              (@              3@                                                              @                                              "@              $@                                                              @                                              @              "@                                                                �t�bub��     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���RhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @$�}8X�?�	           ��@       	                     �?�Z��s��?�           ��@                          �:@WF�o��?�           ��@                           �?:���	F�?,           p�@������������������������       ������#�?b            �d@������������������������       �f6&0%^�?�           P�@                          �@@���rӇ�?g            `f@������������������������       �D�����?_             e@������������������������       ��(\����?             $@
                           �?S��µ�?=           ؚ@                          �<@� 0D�?           �{@������������������������       �@C�E
�?�            �x@������������������������       ��F&K:�?"             K@                            �?�I~&���?%           ܓ@������������������������       ��'o\�?�           ��@������������������������       ��E��[�?i            �@                           @�]���?�           ȑ@                          �4@P�(� �?F           �@                           @�<�
I�?�            �l@������������������������       �]�p�0��?|            �g@������������������������       ���,���?             C@                          @@@EN궍�?�            �q@������������������������       ���BU��?�             q@������������������������       ��q�q�?             (@                          �;@�Mc����?�           ��@                           @�@i!�o�?Z           Ѐ@������������������������       �s��?c�?P           @�@������������������������       �VUUUUU�?
             2@                           @VF$ʬ �?5            �U@������������������������       �����?.            @Q@������������������������       �.k��\�?             1@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@      A@      ;@      4@     �]@     8�@      <@     ��@      .@       @      R@     �J@     8�@     @�@      ,@     �n@      c@      7@      4@      2@      X@      |@      7@     ��@      $@      @     �M@      D@      �@     `y@      "@     �g@     �J@      @      @      "@      B@     �e@      &@     @s@      @              *@      &@     �l@      b@      �?      K@      J@      @      @      @      8@     �c@      $@     �n@      @              &@      $@      f@     @`@      �?     �D@      .@      �?               @      @      5@      @     �O@                      �?       @      <@      0@              @     �B@      @      @      @      4@      a@      @     �f@      @              $@       @     �b@     �\@      �?      A@      �?                       @      (@      0@      �?     �O@      �?               @      �?      J@      .@              *@      �?                       @      (@      *@      �?      O@      �?               @             �I@      (@              (@                                              @              �?                              �?      �?      @              �?      Y@      1@      0@      "@      N@     0q@      (@     @z@      @      @      G@      =@     �s@     Pp@       @      a@      7@      @      @              &@     �N@       @     �U@      @      �?      1@       @     �U@     �U@       @     �G@      5@      @      @              &@      F@      �?     @S@      @      �?      *@      @     @U@     @T@      �?      C@       @       @                              1@      �?      $@                      @      �?       @      @      �?      "@     @S@      &@      $@      "@     �H@     �j@      $@     �t@       @      @      =@      5@     �l@     �e@      @     �V@      D@      �?      @      @      2@     ``@      @     `h@               @      ,@       @     @a@     �S@       @      I@     �B@      $@      @      @      ?@     �T@      @     @a@       @      @      .@      *@     �V@     @X@      @      D@      H@      &@      @       @      6@     �h@      @     �y@      @      �?      *@      *@     �l@     �\@      @      K@      9@      @      @      �?      @     �P@      @     �f@      �?      �?      "@      @     �^@     �H@             �@@      *@      @      @      �?      �?      C@             �P@                      �?              P@      4@              1@       @      @      @      �?      �?      ;@             �K@                                      O@      0@              ,@      @                                      &@              (@                      �?               @      @              @      (@              @              @      =@      @      ]@      �?      �?       @      @      M@      =@              0@      (@              @               @      =@      @      [@      �?               @      @      M@      =@              0@                                      @                       @              �?                                                      7@       @              �?      0@     �`@      �?      l@      @              @      $@     @[@     @P@      @      5@      5@       @              �?      0@     @[@      �?     `f@      @              @      $@      Y@     @P@      @      2@      5@       @              �?      0@      [@      �?      f@      @              @      $@     @W@      M@      @      2@                                              �?              @                                      @      @                       @                                      7@              G@      �?                              "@               @      @       @                                      6@             �@@      �?                              @               @      @                                              �?              *@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJf�AhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @f'X���?�	           ��@       	                    �?�譈t��?N           �@                          �;@�&�?�           �@                            @�ѷDc��?�           t�@������������������������       ���<�?           ��@������������������������       ��3�{ӣ�?�            �p@                           �?���C4�?:             W@������������������������       �     ��?
             0@������������������������       ��Q��X�?0             S@
                           @�DAZ�o�?Q           H�@                            @�����?j            �@������������������������       ���s�9�?p           0�@������������������������       ��a@���?�            �y@                           �?xl3����?�           ��@������������������������       ��V�DJl�?�            �u@������������������������       �΄#����?           py@                            @��B%M�?Z           ��@                          @@@mm���?�           ؅@                          �<@沞����?�           `�@������������������������       �+���ݽ�?�           �@������������������������       �EQEQ�?             E@������������������������       ���A���?             .@                           @��e���?�            0p@                          �5@�[�@�'�?�            @n@������������������������       �@ApAg�?=            �Y@������������������������       ��zN��N�?R            `a@������������������������       �،A��_�?             1@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      7@      G@      ;@     �Z@     ��@      C@     ��@      2@      @     �S@     �K@     ��@     ��@      2@     @n@      d@      *@      D@      9@     �V@     �@      6@     ��@      0@      �?      O@      F@      �@     �v@      ,@     �h@     @Q@       @      1@      4@      9@     `g@      &@     �s@       @              >@      7@     �p@     �d@       @     @R@      P@       @      1@      4@      8@     �e@      &@      q@      @              :@      2@      o@      d@      �?     �Q@     �K@      �?      0@      4@      6@     �`@      "@     @h@      @              5@      2@     �d@     @`@      �?      N@      "@      �?      �?               @     �D@       @      T@                      @              U@      >@              &@      @                              �?      ,@             �C@      �?              @      @      0@      @      �?       @                                              @              @                               @      @      �?                      @                              �?      $@              B@      �?              @      @      $@      @      �?       @     �V@      &@      7@      @     @P@      t@      &@     �@       @      �?      @@      5@     �s@     �h@      (@     �_@      M@      "@      1@       @      E@     �e@      @      p@      @              &@      (@     `i@     @Z@      "@     �T@      :@      @      "@       @      <@      [@      @     �`@                      &@      @     �[@      Q@      @     @P@      @@      @       @              ,@     �P@      @      _@      @                      @      W@     �B@      @      2@     �@@       @      @      @      7@     @b@      @     �o@      @      �?      5@      "@      \@     �V@      @     �E@      0@      �?      @              (@     @T@      �?     @W@       @      �?      $@      @      L@      B@              <@      1@      �?       @      @      &@     @P@      @      d@       @              &@      @      L@     �K@      @      .@      B@      $@      @       @      0@     �g@      0@     �m@       @      @      0@      &@      g@     �f@      @     �E@      :@      @      @       @      ,@      a@      0@      c@       @      @      *@      "@     �`@     �a@      @      C@      8@      @      @       @      ,@     �`@      0@     �b@       @      @      *@       @     �`@     ``@      @      C@      8@      @      @       @      ,@     �_@      0@     �a@       @      @      *@       @     @\@     �_@      @      C@                                               @              "@                                      5@      @                       @                                       @              �?                              �?              "@                      $@      @                       @     �J@             @U@                      @       @      I@     �E@              @      $@      @                       @     �F@             �S@                      @       @     �H@     �D@              @      @      @                       @      *@             �@@                      @      �?      ,@      :@              @      @      �?                              @@              G@                              �?     �A@      .@               @                                               @              @                                      �?       @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJg�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @9+]�{��?�	           ��@       	                   �?@@5n���?�           �@                          �0@�?_So
�?�           b�@                           @0[�-x�?c            �b@������������������������       ��3�a-v�?2            �T@������������������������       ��0!j#;�?1            �P@                           !@��?T           8�@������������������������       �n.���?J           �@������������������������       ����[���?
             2@
                           @��@�4Q�?)            �O@                           �?JC�@��?            �E@������������������������       ��㙢�c�?             7@������������������������       ��G�z��?             4@������������������������       ���Q���?             4@                          �;@,D��C{�?�           d�@                           �?']�֭�?]           �@                          �0@M,1����?           �z@������������������������       ���a_j�?
             3@������������������������       ����Epe�?           �y@                          �9@2�W���?Q           ��@������������������������       ��XA�U��?,           �}@������������������������       �hE#߼�?%             N@                           @
i��f��?d            �b@                           �?�+�wɃ�?$             J@������������������������       �EQEQ�?             5@������������������������       ��-��?             ?@                          �<@Je��{x�?@            �X@������������������������       ��Q����?             4@������������������������       �vb'vb'�?3            �S@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @h@      <@      G@      ?@     �]@     h�@      A@     Ԑ@      2@       @     �T@     @U@     �@     �@      4@     �m@     `c@      6@      <@      ;@     �V@      �@      9@     ��@      *@      @      P@     �Q@     �}@     �w@      2@     �g@      c@      6@      <@      ;@     �V@     ��@      8@     ��@      &@      @      P@     �Q@     p}@     0w@      2@     @g@      "@               @      �?      @     �D@              2@      �?      �?      @      @      ;@      >@              "@      @               @               @      ?@              @      �?              �?       @      2@      0@               @      @                      �?       @      $@              ,@              �?       @      �?      "@      ,@              @      b@      6@      :@      :@     �U@     �~@      8@     �@      $@      @     �N@     �P@     �{@     Pu@      2@      f@      b@      6@      :@      :@     �U@     0~@      5@     �@      $@      @     �N@     �P@     �{@     @u@      2@      f@                                              &@      @      �?                                      �?      �?              �?       @                                      "@      �?      A@       @                      �?      @      @               @       @                                      @      �?      <@       @                              @                       @                                              @              3@                                                                       @                                      �?      �?      "@       @                              @                       @                                              @              @                              �?       @      @                     �C@      @      2@      @      ;@     �e@      "@     �w@      @      @      3@      ,@     �l@     �`@       @     �H@      A@      @      2@      @      6@      a@      "@     �s@      @      �?      3@      *@     @k@     �^@             �F@      4@      @      &@      �?      .@     �P@      @     �]@       @      �?      ,@      @     �T@      P@              8@       @                              �?      �?                                       @       @       @      @              @      2@      @      &@      �?      ,@     @P@      @     �]@       @      �?      (@      �?     @T@     �N@              2@      ,@      @      @      @      @     �Q@      @     @h@      �?              @      $@     �`@      M@              5@      ,@      @      @      @      @     @P@      @     `f@      �?              @      $@     @[@      H@              3@                                      �?      @              .@                                      :@      $@               @      @                              @      B@             �Q@       @       @              �?      *@      $@       @      @                                      @      @              <@               @              �?      @      @               @                                      �?      �?              (@                              �?      �?      @               @                                      @      @              0@               @                      @      @                      @                              �?      ?@              E@       @                              "@      @       @       @                                              "@              @                                       @      �?               @      @                              �?      6@              B@       @                              @      @       @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�	�fhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx                            �;@.��N���?�	           ��@       	                   �0@�^�_��?�           �@                           �?��?"md�?�            �o@                           �?��)V��?;            @V@������������������������       �JG��S��?#             K@������������������������       ��l8b��?            �A@                            @�`��[�?Z            `d@������������������������       �����n��?H            @`@������������������������       �^1�[��?            �@@
                           �?(tU���?            �@                            @lZ�3�;�?�           ��@������������������������       �A�}�an�?�           ��@������������������������       ���x�|�?�            @x@                            @�-�@��?�           ��@������������������������       ���=��?8           ��@������������������������       ���&`��?J           �~@                           @�KyU#\�?           �{@                           �?Ѧr�X��?           @{@                           @j]���~�?)            �Q@������������������������       �x9/���?!             L@������������������������       ��$I�$I�?             ,@                           @��|**4�?�            �v@������������������������       ��������?�            �t@������������������������       �H�%s��?            �A@������������������������       �                     "@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      6@     �C@      8@     @]@     �@     �B@     ��@      0@      "@     �Q@     �L@     ��@     P@      .@     �r@     �h@      2@     �B@      8@      [@     ��@     �A@     0�@      .@      @     @P@     �I@     P�@     `}@      *@     pq@      *@               @       @      1@      K@       @     �D@                      @      $@     �G@      A@              8@      �?              �?      �?      (@      6@      �?      @                      @      @      0@      0@               @                      �?      �?      (@      "@      �?      @                      @       @      $@      $@              �?      �?                                      *@              @                       @      @      @      @              �?      (@              �?      �?      @      @@      �?      A@                      �?      @      ?@      2@              6@      $@              �?      �?       @      <@      �?      7@                      �?      @      <@      *@              2@       @                              @      @              &@                              �?      @      @              @     �f@      2@     �A@      6@     �V@     �@     �@@     �@      .@      @     �M@     �D@     ؂@     @{@      *@     �o@     @W@      "@      6@      0@     �G@     �n@      1@     pu@      &@      @      >@      5@     `o@     `h@      @      a@     �R@      @      0@      .@      >@     `g@      &@     @m@      $@      @      :@      3@     �e@     �a@      @     �[@      2@      @      @      �?      1@     �M@      @     @[@      �?              @       @     �S@      K@              :@     �V@      "@      *@      @      F@     �p@      0@     0�@      @       @      =@      4@      v@      n@       @     �]@      R@      @       @      @      C@     `i@      ,@     @v@       @       @      <@      ,@     �l@      h@      @     �X@      2@       @      @      �?      @     @P@       @     @h@       @              �?      @     @^@      H@      �?      3@      9@      @       @              "@     @R@       @     @g@      �?      @      @      @     �Q@      ?@       @      7@      9@      @       @              "@     @R@       @      f@      �?      @      @      @     �Q@      ?@       @      7@      @                                      3@              4@                       @       @      (@      @              @      @                                      &@              2@                       @       @       @      @              @                                               @               @                                      @                              2@      @       @              "@      K@       @     �c@      �?      @      @      @     �M@      <@       @      2@      2@      @       @              "@      J@       @     �`@      �?      @      @      @      J@      ;@       @      2@                                               @              8@                              �?      @      �?                                                                              "@                                                                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�ǿAhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?f)���l�?�	           ��@       	                   �1@�5����?           X�@                          �0@��R���?�             r@                            �?:}R���?>            @Y@������������������������       �     $�?$             P@������������������������       �u�t��?            �B@                            @��7�B��?w            �g@������������������������       ��$��(�?[            `b@������������������������       �U�	�S�?             E@
                           @w��|��?i           Е@                           @������?�           ��@������������������������       �f�}����?1           @�@������������������������       �.�F���?i            �d@                            @\=ӇS��?�            pt@������������������������       �WШ��?�             n@������������������������       �s�k����?4            �U@                            @&��y��?x           f�@                           @��qMu�?�           ��@                          �7@o���|��?           �@������������������������       �,d����?            �@������������������������       �������?�            �w@                            �?���(h��?�            �v@������������������������       ��������?F             ^@������������������������       ���m�L��?�            �n@                          �5@��8��?�           �@                           @�\���?�            �r@������������������������       ��]t�l�?�            0q@������������������������       �p�u=q��?             7@                           @�en���?�            �u@������������������������       �ᦛ?�?�            �l@������������������������       ��QDr	�?>            �\@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �f@      C@      ?@      ;@     �U@     ��@      B@     l�@      .@      *@     @T@     �L@     ��@     ��@      0@     �p@     �T@      4@      4@      2@     �J@     Pq@      5@     px@      *@       @      A@      <@     �u@     �l@      @     �`@      3@      �?      @      @      *@      C@      @      C@      @       @      @       @     �N@     �H@              B@      @                      @      @      &@      @      &@              �?      @       @      ;@      7@              @      @                      @      @      "@       @      @                              �?      5@      (@              @      @                               @       @      �?      @              �?      @      �?      @      &@               @      *@      �?      @              @      ;@      @      ;@      @      �?      @      @      A@      :@              ?@      (@      �?      @              @      2@      @      ,@      @      �?      @      @      :@      6@              9@      �?              �?                      "@              *@                                       @      @              @      P@      3@      .@      .@      D@     �m@      .@     v@      "@      @      ;@      4@     �q@     �f@      @     �X@     �J@      1@      .@      .@      B@     �e@      @      q@      @      �?      9@      2@     �l@     @_@      �?      S@     �G@      0@      ,@      *@      <@      b@      @     �l@      @      �?      4@      *@     �i@      W@      �?     @Q@      @      �?      �?       @       @      >@      �?     �D@                      @      @      9@     �@@              @      &@       @                      @     @P@      $@     @T@      @      @       @       @     �L@     �L@      @      6@      "@       @                       @     �I@      $@      I@      @               @       @     �B@      G@      @      5@       @                               @      ,@              ?@              @                      4@      &@              �?      Y@      2@      &@      "@      A@     �u@      .@     ��@       @      @     �G@      =@     �{@     �r@      "@     �`@      U@      1@       @       @      9@     0p@      ,@     P|@      �?      @      F@      8@     �r@     �k@      "@     �\@     �R@      *@      @      @      *@     �k@      *@     `t@              @     �A@      2@     `m@     �f@      @      Q@     @P@      @      @      @       @     @c@      @      i@              @      2@      *@     �c@     @a@      @      I@      "@      @      �?      �?      @     �P@      @     @_@              �?      1@      @      S@      F@       @      2@      $@      @      @      �?      (@     �C@      �?     �_@      �?              "@      @     @P@      C@       @      G@       @      @              �?              @             �N@      �?              @              7@      *@      �?      @       @              @              (@      @@      �?     �P@                      @      @      E@      9@      �?      E@      0@      �?      @      �?      "@      V@      �?     �p@      �?      �?      @      @     �a@     �S@              5@       @              @      �?      @      G@      �?     �X@                       @      @     �Q@      G@              .@       @              @      �?      @      F@      �?     @T@                       @      @      Q@      G@              ,@                                               @              2@                                       @                      �?       @      �?                      @      E@             �e@      �?      �?      �?       @     @R@     �@@              @      @      �?                      @      5@              `@              �?      �?              H@      ,@              @      �?                                      5@             �E@      �?                       @      9@      3@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJJ��JhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?s>#�s�?�	           ��@       	                    @5��?a           ��@                          �1@MZ��;�?t           H�@                           @rw����?�             o@������������������������       �x9/���?�             l@������������������������       ��������?             8@                           @��j���?�           h�@������������������������       �R����?b           ��@������������������������       ��j}s�)�?s            �h@
                            �?2��-��?�            �v@                           �?@�(ݾ2�?�             j@������������������������       ��5?,R�?             B@������������������������       ���u�-�?o            �e@                           @���e�?e            `c@������������������������       �{�1��8�?G            �Z@������������������������       ��q�q\�?             H@                          �;@�D){���?_           ��@                           @�M&��?�           ��@                            @�X�����?           ��@������������������������       ��j^'=�?u           `�@������������������������       ��A�^�T�?�            �l@                           !@��
8WI�?�           Ȑ@������������������������       �?�Bu�H�?�           ��@������������������������       �9��8���?             (@                           @�'��?�            �l@                           @��8���?�             h@������������������������       �0�od N�?i             c@������������������������       ���/5�?            �C@                           �?���?            �C@������������������������       �     ��?             0@������������������������       ���<b���?             7@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      =@      F@      9@      X@     ��@      B@     ��@      7@      (@     �S@     �I@     ��@     �@      4@     �n@     �\@      2@     �A@      &@      N@     �s@      3@     �|@      *@      @      A@      ;@     �s@     �k@      &@     �_@     �W@      *@      @@      &@     �K@     `o@      @      w@      (@      @      ?@      8@     0p@      c@       @     �Y@      .@      �?      @      �?      &@     �D@      @      D@      �?       @      @      @      G@      D@      @      ;@      .@      �?      @      �?      &@      D@      @      ?@      �?       @       @      @     �F@     �@@      @      7@                                              �?              "@                      �?      �?      �?      @              @      T@      (@      9@      $@      F@     @j@       @     �t@      &@      @      <@      4@     �j@     @\@      @      S@     �N@      "@      3@       @     �@@      e@       @     �q@      &@      @      ;@      0@     @g@     �V@      @     �O@      3@      @      @       @      &@     �D@             �G@                      �?      @      ;@      7@              *@      4@      @      @              @     �P@      *@     �W@      �?      �?      @      @      L@     �P@      @      7@      .@      @       @              @     �F@      $@     �F@                       @      �?      =@      ?@      @      0@      �?      @                      �?      @              2@                                      @                       @      ,@      �?       @              @      E@      $@      ;@                       @      �?      6@      ?@      @      ,@      @              �?              �?      5@      @     �H@      �?      �?      �?       @      ;@      B@              @      @                              �?      0@      @      B@              �?      �?       @      0@      8@              @      �?              �?                      @              *@      �?                              &@      (@              @     @Z@      &@      "@      ,@      B@     ps@      1@     �@      $@      @      F@      8@     |@     �q@      "@      ^@     @Y@      $@      "@      *@     �A@     �p@      ,@     �@      @      @     �C@      7@     �x@     0q@       @      \@     �I@      @      @      @      .@     �Y@      @     �p@       @              $@      $@      h@     �X@       @     �H@     �F@      @      @      @      ,@     @T@      @      e@       @               @      @      a@      R@       @     �B@      @              �?      @      �?      5@              Y@                       @      @      L@      :@              (@      I@      @       @      @      4@      e@      &@     Ps@      @      @      =@      *@     �i@      f@      @     �O@      I@      @       @      @      4@     `d@      &@     @s@      @      @      =@      *@     �i@     �e@      @     �O@                                              @              �?                                       @      @                      @      �?              �?      �?      D@      @      X@      @      @      @      �?     �I@      &@      �?       @      @      �?              �?      �?     �B@      @      R@      @      @      @      �?     �D@      &@      �?       @      @      �?              �?      �?      8@      @      P@      @      @      @      �?      <@      @      �?       @                                              *@               @                                      *@      @                                                              @              8@                       @              $@                                                                      @              @                       @              @                                                                                      2@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�I^shG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?���k�z�?�	           ��@       	                    @�N�H)�?L           D�@                            @�[E,�?�           ��@                          �=@�YI}��?           ��@������������������������       �`mu���?�           �@������������������������       �g�WH��?             ;@                           �?<�Ӎ���?�             w@������������������������       �xJ'�L�?�            �n@������������������������       ��<��?V             _@
                           @`*�Kr��?r           �@                           �?���98�?�            �p@������������������������       �<۪zJ�?7            @U@������������������������       ����hz�?{            �f@                            �?$��+��?�            pq@������������������������       ���')>Y�?g            `b@������������������������       ���wC���?Y            �`@                            @̠�0���?e           �@                           @L���p�?�           ��@                            �?�z���|�?D           D�@������������������������       �qQ��Y��?�           (�@������������������������       ���;5��?�            �r@                           @/��mԚ�?�            `k@������������������������       ��p)���?E             [@������������������������       �'�[���?G            �[@                          �2@B�)���?�           `�@                          �0@L���Y&�?l            �e@������������������������       ��8��8��?             8@������������������������       �Q��<J�?_            �b@                          @@@��b�/��?)            ~@������������������������       ��a!����?           �|@������������������������       �6�80\��?             3@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `e@      @@     �E@      ?@     @\@     ��@      ;@     4�@      .@      @     �P@     �Q@     ��@     x�@      5@     �p@     @W@      .@      =@      *@     �N@     `r@      1@     �y@      "@      @      ;@     �D@     �t@      m@      *@      c@     �M@      $@      8@      $@     �J@     �i@       @     0q@      @      @      3@      :@     `n@     `a@      @     �[@     �H@      @      ,@      "@     �E@     @c@      @     �e@      @      @      2@      8@     �a@     @V@      @     �U@     �G@      @      ,@      "@      D@      c@      @      d@      @      @      2@      8@     @a@      U@      @     �U@       @                              @      �?              ,@                                       @      @                      $@      @      $@      �?      $@     �J@      @      Y@                      �?       @     �Y@      I@              7@      @      @      @              @      =@      @     �Q@                      �?       @      S@      9@              .@      @              @      �?      @      8@              =@                                      ;@      9@               @      A@      @      @      @       @     �U@      "@      a@       @               @      .@     �V@     �W@      @     �E@      ;@      @      @      �?      @      F@      @     �N@       @              @      @     �A@      H@              7@      @                      �?       @      *@      @      9@      �?              @              3@      @              @      6@      @      @              �?      ?@      @      B@      �?                      @      0@      E@              0@      @       @       @       @      @     �E@       @     �R@                      @      "@     �K@      G@      @      4@      @      �?      �?       @      �?      ;@       @      <@                      @      @      7@      ;@       @      0@       @      �?      �?              @      0@             �G@                               @      @@      3@      @      @     �S@      1@      ,@      2@      J@     �u@      $@     ��@      @      @     �C@      =@     @|@     `r@       @     @\@      O@      .@      "@      ,@      F@     �n@       @     �z@       @      @     �A@      6@     �r@      l@       @     �X@     �N@      *@       @      (@      @@     �j@       @     �u@       @      @      >@      3@     �o@     @j@      @     �R@      E@      &@      @      $@      2@     �d@      @     �r@      �?              6@       @      j@     �c@      �?      H@      3@       @      @       @      ,@     �H@       @      K@      �?      @       @      &@      G@      K@      @      :@      �?       @      �?       @      (@      @@             �R@                      @      @      G@      ,@      @      8@                      �?       @      &@      .@              C@                              �?      :@       @              @      �?       @                      �?      1@              B@                      @       @      4@      @      @      2@      0@       @      @      @       @     �X@       @     �p@      @              @      @     �b@     �Q@              .@      @              �?      @       @      (@              Q@                      �?      �?      K@      5@              @                                               @              *@                                      @      @              �?      @              �?      @       @      $@             �K@                      �?      �?      I@      1@              @      (@       @      @      �?      @     �U@       @     �h@      @              @      @     @X@     �H@              $@      &@       @      @      �?      �?     �U@       @     �g@      @              @      @      W@     �H@              $@      �?                              @                       @                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ?ZhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @bZo�-��?�	           ��@       	                     �?y�O��?�           ��@                           @ns�#��?{           (�@                           @U�1���?�           (�@������������������������       �H� �U��?*           p|@������������������������       �j� ��?a            �c@                           �?�8��8J�?�             x@������������������������       �ŀz	k�?Z            �a@������������������������       ���|i��?�             n@
                          �1@�z��n�?{           \�@                           @�������?�            pt@������������������������       �e/H�n��?w            �f@������������������������       ��a�2�4�?]             b@                           @bk4�"D�?�           @�@������������������������       �Õ jzQ�?           ��@������������������������       ��?N�ю�?�            �m@                           �?���3�?�           4�@                           @���q�?G           8�@                           @6���Y�?5           �~@������������������������       �k���&^�?	           `z@������������������������       �*p긹��?,            @Q@������������������������       ��m۶m��?             <@                          �2@�:�D��?|           0�@                           �?2���o�?l            �d@������������������������       �Sl �?'            �K@������������������������       ��6Z���?E            �[@                           �?�|��_�?           z@������������������������       �N�p3*<�?-            �P@������������������������       �(p7O��?�            �u@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �l@      <@     �C@      6@     �Y@     h�@      @@     �@      1@      @     @S@     �K@     X�@      �@      A@     pp@      f@      4@      <@      4@     �S@     �{@      9@     8�@      *@      @     �P@     �E@     P@     �z@      ?@     �k@      J@       @      @      @      7@      e@      *@     Ps@      @              .@       @     `h@     �a@      "@     �D@     �B@      �?      @      @      2@      \@      @     `i@      �?              @      @     @\@     �R@      @      <@      <@      �?      @      @      0@      W@       @     �a@      �?               @      @      W@     �H@       @      1@      "@                               @      4@       @      O@                      �?       @      5@      9@      @      &@      .@      @      �?       @      @      L@      "@     �Z@      @              (@       @     �T@     �P@      @      *@       @      �?      �?              @      2@      �?      A@      @              @              A@      <@       @      @      @      @               @       @      C@       @      R@                      "@       @      H@     �C@       @      @     @_@      (@      8@      *@      L@     Pq@      (@      y@      "@      @      J@     �A@      s@     �q@      6@     �f@      5@       @      @               @      J@      �?      G@      �?       @      1@      $@     �K@      N@      @      C@      *@       @      @              @      A@      �?      3@      �?              (@      @     �@@      8@      @      ;@       @              @              @      2@              ;@               @      @      @      6@      B@      @      &@      Z@      $@      1@      *@      H@      l@      &@     @v@       @       @     �A@      9@     `o@     @l@      .@     �a@     @U@      $@      0@      $@     �@@      h@      "@     0r@      @       @      >@      8@     �h@     �i@      .@     �^@      3@              �?      @      .@     �@@       @     @P@      �?              @      �?     �J@      3@              3@     �I@       @      &@       @      8@      f@      @     �w@      @       @      $@      (@     �n@     @^@      @      E@      D@      @      @       @      2@     �W@      @     �a@      �?       @      @      @     @Z@      O@              7@      C@      @      @       @      ,@     @V@      @     @a@      �?       @      @      @     @Y@      L@              5@     �@@      @      @       @      *@     �R@      @     �\@      �?              @      @     �V@     �H@              5@      @      @      �?              �?      ,@      �?      7@               @               @      $@      @                       @                              @      @              @                                      @      @               @      &@       @      @              @     �T@      @     �m@      @              @      @     �a@     �M@      @      3@      @               @              �?      5@             �J@                      �?             �N@      0@              @                                               @              2@                                      9@      "@              �?      @               @              �?      3@             �A@                      �?              B@      @              @      @       @      @              @     �N@      @     @g@      @               @      @      T@     �E@      @      *@       @              �?                      &@      �?      5@                                      *@      ,@              @      @       @       @              @      I@       @     �d@      @               @      @     �P@      =@      @      "@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��4hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @+������?�	           ��@       	                    �?L�*`�?�           <�@                            �?h&�׍�?           ̓@                           �?d9��Z�?W           �@������������������������       �� ���?R            �_@������������������������       �:���H�?           (�@                           @�	"P7��?�             s@������������������������       ��|�l%�?�             q@������������������������       �     ��?             @@
                            �?R�]Yhq�?�           ��@                          �@@Z������?�           �@������������������������       ��45�h��?�           ��@������������������������       �333333�?             $@                           @�M���?�            @v@������������������������       ���E>D�?k            @d@������������������������       ���`����?t            @h@                          �2@/X7�?�           ��@                          �1@�K�;(h�?�            @p@                           @����+�?W            �a@������������������������       �#JS��%�?0            @S@������������������������       �     d�?'             P@                           @N ?sI��?Q            �]@������������������������       �?��K>7�?-            �P@������������������������       �1(?cwr�?$            �J@                           �?�3�����?�           8�@                           @5�?7�?�            �u@������������������������       �     ��?�             p@������������������������       �����<�?4            �V@                          �3@Ξ�X[��?           �|@������������������������       ��
�'��?'            @P@������������������������       ��X	���?�            �x@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      D@      F@      <@      [@     ��@      C@     ܐ@      ,@      .@     @S@      M@     ��@     ��@      7@     �l@      d@      @@      A@      :@     @U@     ~@     �@@     �@      $@      $@     @Q@     �C@     x�@     �y@      5@     �h@     @V@      ,@      :@      (@     �I@     �m@      .@     �p@      @      @      B@      4@     @j@     �e@      "@     �X@     �Q@      "@      7@      "@      D@     �h@       @     `i@      @              =@      (@      d@     @_@      @      O@      @       @      �?       @      @      .@             �B@                      *@      @      6@      "@              "@      P@      @      6@      @      A@      g@       @     �d@      @              0@      "@     `a@      ]@      @     �J@      2@      @      @      @      &@     �B@      @      O@      �?      @      @       @     �H@     �G@      @     �B@      2@      @       @      @      &@      A@      @     �E@      �?      @      @       @     �H@      C@      @     �B@                      �?                      @              3@                                              "@                     �Q@      2@       @      ,@      A@     �n@      2@     �{@      @      @     �@@      3@     �s@     @n@      (@     �X@     �H@      2@      @      (@      1@      g@      (@     �w@       @              6@      &@     �o@     �f@      @      Q@     �H@      2@      @      (@      1@     `f@      (@     �w@       @              6@      $@     �o@     `f@      @     �P@                                              @                                              �?      �?      �?              �?      6@              @       @      1@      N@      @     �M@      �?      @      &@       @      O@      O@      @      ?@      $@              @      �?      @      1@              :@      �?      @       @      �?      C@      >@      @      4@      (@              �?      �?      (@     �E@      @     �@@                      "@      @      8@      @@      @      &@     �F@       @      $@       @      7@      j@      @     @w@      @      @       @      3@     �h@      `@       @      >@      &@              �?       @      @     �D@             �R@                      �?      "@     @R@      >@              *@       @                              @      ;@              D@                      �?      "@      =@      .@               @       @                                      3@              :@                      �?              3@      @              @      @                              @       @              ,@                              "@      $@      "@              @      @              �?       @              ,@             �A@                                      F@      .@              @      @                                      @              .@                                      A@      @               @                      �?       @              @              4@                                      $@      $@              @      A@       @      "@              3@     �d@      @     �r@      @      @      @      $@     @_@     �X@       @      1@      5@      @      @              (@     �R@       @     �Y@      @      @      @      �?      G@     �J@       @      $@      5@      @      @              "@     �M@       @     �O@      @      @      �?      �?      A@     �E@       @      @              �?       @              @      0@             �C@                      @              (@      $@              @      *@      @       @              @      W@      @     `h@      �?       @      �?      "@     �S@     �F@              @       @                              �?      "@      @     �@@                                      @      @                      @      @       @              @     �T@             @d@      �?       @      �?      "@      R@     �D@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJk�� hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @���?�	           ��@       	                     �?�9����?�           ��@                            �?�˶��?@           ��@                           �?x?}���?~           ��@������������������������       ��cR3?�?j            �d@������������������������       ���)o��?           ��@                           �?ru�<��?�           ��@������������������������       ����;\I�?�            �u@������������������������       �ސ4q���?�           H�@
                           @ҞoZ{��?�            �@                           �?��|YN�?�            �j@������������������������       �s��F�?J            @Z@������������������������       ��u�Ë��?A             [@                          �4@�+u���?           �z@������������������������       ��(�A��?�            �o@������������������������       ���޶�,�?u            `f@                           �?�J���?�           ��@                          �8@�����Z�?F           0�@                           �?��8���?�             x@������������������������       ��@8ݓ��?/            @R@������������������������       �<b&:�d�?�            ps@                           �?�XO��?Z            �`@������������������������       ����^B{�?             2@������������������������       ���_�#3�?J             ]@                           �?٥@�q�?�           �@                           �?!�#���?�            �x@������������������������       �f1�����?<            �V@������������������������       ���[���?�            �r@                           @RQY�?�            @k@������������������������       �~�U92��?9            @V@������������������������       ��L��}
�?W             `@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      ?@     �B@      7@     �T@     ��@      @@     L�@      5@      @     �W@      P@     0�@     �@      2@     �p@     �d@      8@      8@      2@     �Q@     p|@      9@     P�@      0@      �?     �S@      M@     �@      x@      0@     �k@      a@      *@      2@      0@      J@     pw@      6@     ��@      (@      �?     �G@      =@     y@     �p@      $@     �a@     �N@      @      �?      (@      0@     �d@       @     Pt@      @              .@      ,@     @i@     ``@      @     �G@      @                       @      @      4@      �?      N@                      @             �@@      0@              .@     �K@      @      �?      $@      (@     `b@      @     �p@      @               @      ,@      e@     �\@      @      @@     �R@      @      1@      @      B@      j@      ,@     q@      @      �?      @@      .@     �h@     @a@      @     �W@      4@      @      @      @      *@      D@      �?      T@      �?              ,@      @     �P@      L@       @     �B@     �K@       @      *@              7@      e@      *@      h@      @      �?      2@      $@     �`@     �T@      @     �L@      <@      &@      @       @      2@      T@      @      ]@      @              @@      =@     �[@     @]@      @     �T@      @      @       @      �?      @      5@      �?      D@      @              0@      @     �H@      @@       @      =@              @              �?      �?      3@      �?      2@      @              @      �?      6@      *@       @      2@      @       @       @              @       @              6@                      *@      @      ;@      3@              &@      8@      @      @      �?      ,@     �M@       @      S@      �?              0@      9@     �N@     @U@      @     �J@      $@      @      @      �?      @      C@      �?      B@                      &@      1@      5@     �M@      @     �D@      ,@      �?      �?              "@      5@      �?      D@      �?              @       @      D@      :@              (@      E@      @      *@      @      *@     �f@      @     �x@      @      @      .@      @     pp@     @_@       @     �G@      >@      @       @      @      $@     @W@      @     �`@       @      @      $@      @     @_@     �M@      �?      9@      ,@      @      @      @      $@     �R@      @     �T@              @      $@      @      X@     �H@              6@      @                              @      $@              3@                      @      �?      ,@      $@              @      "@      @      @      @      @     @P@      @     �O@              @      @      @     �T@     �C@              .@      0@      �?       @                      2@             �I@       @                      �?      =@      $@      �?      @       @              �?                      @              @                                      @       @                      ,@      �?      �?                      *@             �G@       @                      �?      9@       @      �?      @      (@      @      @      �?      @     �V@      �?     @p@      @              @      �?     @a@     �P@      �?      6@      @              @      �?       @      P@      �?     `d@      @              @      �?      R@     �I@      �?      4@       @              @              �?      &@      �?      B@                                      .@      .@              @      @                      �?      �?     �J@             �_@      @              @      �?     �L@      B@      �?      *@      @      @       @              �?      :@             @X@                      �?             �P@      .@               @       @               @              �?      "@              A@                                     �C@       @                      @      @                              1@             �O@                      �?              ;@      *@               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�x4lhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @����?�	           ��@       	                     �?����?�           �@                           @�asM��?�           Ԑ@                           �?�7�h���?           @�@������������������������       ���v/FO�?�            �s@������������������������       ����]��?E           ��@                           @�$����?�            �m@������������������������       �B{	�%��?             "@������������������������       �{[����?�            �l@
                          �1@�#�;d�?[           `�@                          �0@n��@��?�            v@������������������������       ��jt����?E            �]@������������������������       �rT=�^�?�            `m@                            �?<�j6	/�?�           ܕ@������������������������       ��+���?1           Ȋ@������������������������       � &'A���?W           ��@                           @�*��D�?�           �@                           �?�c�;��?A           �@                           �?���U��?�            t@������������������������       ��,F�z�?t             f@������������������������       ��n�K�?W             b@                          �6@<T��~��?v            @h@������������������������       �tٻ��?D            @Z@������������������������       �_��0e�?2            @V@                          �5@�ϬjQ�?v           ȁ@                           �?��P��?�            `o@������������������������       �$M=ֱ��?T            �\@������������������������       ���Ooo6�?Z             a@                           @�����?�            �s@������������������������       ������?�             n@������������������������       �H�~�?5            @S@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      ;@      E@      ,@     �Z@     �@      >@     8�@      3@      &@     @T@     �Q@     p�@     x�@      5@     �o@      c@      6@      ?@      *@     @U@     �~@      6@     ��@      ,@      "@     �Q@      N@     �@      y@      2@     @j@      H@      $@      @      @      8@      i@      $@     pt@      @              .@      0@     �j@     �a@      @     �H@     �@@      @      @      @      2@     �c@      $@     �n@      @              *@      $@     �e@      _@       @      @@      &@              �?      �?      (@     �K@      @      V@      �?              @       @      N@      H@       @      0@      6@      @      @      @      @     �Y@      @     �c@      @              @       @     �\@      S@              0@      .@      @              �?      @      E@             �T@      �?               @      @     �C@      0@      @      1@                                              �?              @                      �?                                              .@      @              �?      @     �D@              S@      �?              �?      @     �C@      0@      @      1@     @Z@      (@      8@       @     �N@     r@      (@     �x@      "@      "@     �K@      F@     pr@     `p@      &@      d@      5@      @      @      �?      *@     �R@      @      H@      @      @      *@      (@     �I@     �N@       @      B@      @      �?       @      �?      @      3@              $@       @      @      @      @      (@      =@      �?      0@      1@       @      @              @      L@      @      C@      �?      �?       @      @     �C@      @@      �?      4@      U@      "@      2@      @      H@     �j@       @     �u@      @      @      E@      @@     �n@      i@      "@     @_@     �I@       @      (@      @      7@     �b@      @     `l@                      :@      1@     �c@     @[@      @     @R@     �@@      @      @      @      9@     �P@       @      ^@      @      @      0@      .@     �U@      W@      @      J@     �A@      @      &@      �?      6@     �f@       @     �w@      @       @      &@      $@      n@     @_@      @     �F@      (@              @      �?      "@     �P@      �?     �f@              �?       @      @     @a@     �N@              8@      @                              @     �J@      �?     �Z@                      @       @     �T@      G@              1@      @                              @     �C@      �?     �H@                      @       @     �E@      6@              @                                              ,@             �L@                                     �C@      8@              $@      @              @      �?      @      ,@             @S@              �?      @      �?      L@      .@              @      @              @      �?       @      $@              @@                      @             �@@      &@              @      �?              @              @      @             �F@              �?              �?      7@      @               @      7@      @      @              *@     @\@      @     �h@      @      �?      @      @     �Y@      P@      @      5@      $@      �?       @               @      B@      @      V@       @      �?      @      @     �G@      ?@              (@      @      �?                      @      (@      @      C@              �?               @      7@      .@              "@      @               @              @      8@       @      I@       @              @      @      8@      0@              @      *@      @       @              @     @S@       @     @[@      @                       @      L@     �@@      @      "@      (@      @       @              @     �L@       @     @V@       @                       @      A@      7@      @      @      �?                              �?      4@              4@      �?                              6@      $@               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJt+hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �:@'��g��?�	           ��@       	                     @�@���?M           (�@                           �?iw��4!�?�           Ģ@                           @�4�ͯ��?�           h�@������������������������       �ٔ�٨�?6           0�@������������������������       �D˩�m��?b            �b@                           @z�G�n��?Z            �@������������������������       ��?�4���?           ��@������������������������       ��@f�y2�?J           `@
                           �?l��q���?[           ��@                           @��a��?           pz@������������������������       ��t�Yl��?�            �x@������������������������       �V}��b�?             9@                          �9@��9�C��?S           X�@������������������������       �
�o��p�?7            ~@������������������������       �z3�Vf`�?            �D@                           @&����?n           ��@                           �?���L��?A           �~@                          �<@{y��?�            �h@������������������������       ���#�X��?8            �W@������������������������       �
٭�\��?K            @Z@                            �?�e���?�            Pr@������������������������       ���Fe;�?0            �S@������������������������       ��^��cQ�?�            �j@                           �?��dc�_�?-            @R@������������������������       �z3����?
             5@                          �;@.�T�6�?#             J@������������������������       �      �?              @������������������������       ��E]t��?             F@�t�b��     h�h4h7K ��h9��R�(KKKK��h��B�       �j@      E@      C@      9@      [@     ��@      D@     X�@      :@      @     �U@      K@     ��@     �}@      1@     Pq@     �g@      >@     �A@      8@     �W@     0�@     �A@     �@      3@      @     �S@      I@     Ȃ@     `{@      .@     �o@      b@      0@      :@      4@     @R@     0z@      <@     ��@      1@      �?     @Q@     �F@     �y@     pt@      ,@     �h@     �S@      $@      2@       @     �D@     �h@      &@      k@      0@      �?      ?@      :@     @e@      a@      @      U@      P@      $@      2@      @      <@     �c@      &@     `g@      0@      �?      ?@      8@      d@     @\@      @     @Q@      .@                      �?      *@     �C@              =@                               @      $@      8@              .@     @P@      @       @      (@      @@     �k@      1@     �w@      �?              C@      3@      n@     �g@      "@     �\@      E@      @      @       @      0@     �a@      @      j@      �?              6@      (@      g@     �_@      @      Q@      7@      @      �?      @      0@     @T@      &@      e@                      0@      @      L@     �O@      @     �G@      G@      ,@      "@      @      6@     `d@      @      s@       @       @      $@      @     �g@     �[@      �?      L@      ;@      @      @      �?      .@     �V@      @     @Y@       @       @      @      �?     @S@      K@              =@      9@      @      @      �?      (@     �U@      @     �X@       @       @      @      �?     @Q@      H@              <@       @                              @      @               @                                       @      @              �?      3@      @       @      @      @     @R@      @     `i@                      @      @     @\@     �L@      �?      ;@      3@      @       @      @      @     �Q@      @      h@                      @      @      X@      J@      �?      8@               @                      �?       @              &@                                      1@      @              @      7@      (@      @      �?      *@     @[@      @     �j@      @       @      @      @     @Y@     �D@       @      6@      7@      (@      @      �?      (@      Y@      @      e@      @       @      @      @     @V@      C@       @      3@      (@      &@      @      �?      @      @@      @     �O@       @              @      �?      ;@      9@              $@      @      "@      �?      �?              4@      @      9@      �?              �?              1@      "@              @       @       @       @              @      (@              C@      �?              @      �?      $@      0@              @      &@      �?                       @      Q@       @     @Z@      @       @       @      @      O@      *@       @      "@      �?                               @      *@       @      9@       @                              :@      @              @      $@      �?                      @     �K@              T@      @       @       @      @      B@      "@       @      @                                      �?      "@             �F@                                      (@      @              @                                      �?       @              @                                      @                                                                      �?              C@                                      @      @              @                                              �?              @                                               @               @                                                             �A@                                      @      �?              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJH�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�T���i�?�	           ��@       	                   �<@��aH�0�?E           h�@                            @�@z�y3�?�           (�@                           �?wM�<0��?�           �@������������������������       ���ǟd��?           {@������������������������       �"-�COE�?�           ��@                          �6@R�f��%�?           �|@������������������������       �?"J'��?�            �s@������������������������       �P�G�� �?X            `a@
                           @�5?,R��?S             b@                           @�j�~%W�?A            �\@������������������������       �Z�g{��?2             W@������������������������       ��nkK�?             7@                            �?�n��>�?             =@������������������������       �;�;��?	             *@������������������������       �      �?	             0@                          �;@�Ss���?_           ޠ@                            @L��z��?�           ��@                           @0�ѩeB�?a           <�@������������������������       �xRa�85�?\           x�@������������������������       ��K8#�?            z@                           @�����?V           �@������������������������       ��&k'(�?�            �m@������������������������       �%U����?�            s@                            �?6
e��?�            0p@                          �?@vʾ��?4            �U@������������������������       �<�g���?&            @P@������������������������       ��Ra����?             6@                           @�YeD��?t            �e@������������������������       �c��-8�?Q            �_@������������������������       ��=��h��?#             G@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@     �B@      C@      9@     �W@     ��@      :@     ��@      4@      @     �P@     �P@     ��@     �~@      4@     �n@     �[@      9@      8@      *@     �L@     @t@      .@     �y@      (@      @     �B@     �D@     �s@      m@       @     �_@     �V@      3@      7@      *@      K@     ps@      .@     @v@      $@      @     �A@      C@     `r@     �k@      @     �^@      R@      $@      4@      &@     �H@     `l@      "@     �l@      "@      @      =@      @@     @h@     �d@      @     �V@      >@       @      @      @      8@      U@      �?      S@      @       @      ,@      "@      M@     @R@       @      C@      E@       @      *@      @      9@     �a@       @      c@      @      �?      .@      7@      a@     �V@      @     �J@      2@      "@      @       @      @      U@      @      `@      �?      �?      @      @      Y@     �L@              ?@      (@      @       @       @      @      E@      @     @W@              �?      @      @     @S@     �@@              =@      @       @      �?                      E@      @     �A@      �?                              7@      8@               @      4@      @      �?              @      *@              J@       @               @      @      7@      (@      @      @      0@      @      �?              @      *@             �B@       @               @      @      5@      @      @      @      ,@      @      �?              �?      *@             �@@       @               @      @       @       @      @      @       @                               @                      @                                      *@       @                      @                                                      .@                                       @       @                                                                              @                                       @      @                      @                                                      $@                                               @                     �Y@      (@      ,@      (@     �B@     �u@      &@     p�@       @      @      >@      :@     �{@     `p@      (@     �]@     @W@      $@      ,@      (@      A@     �q@      "@     (�@      @      �?      =@      6@     py@     �n@      &@     �Z@     �Q@      $@      "@      $@      ?@     �j@      "@     �x@      @      �?      :@      .@      r@     �f@      "@     �U@      M@      @      @      "@      .@     @d@      @     p@      @      �?      0@      "@     @j@     �`@      @     �G@      *@      @      @      �?      0@     �J@      @     �`@                      $@      @      T@     �F@      @      D@      6@              @       @      @      R@             �k@       @              @      @     @]@     @P@       @      4@       @               @      �?      �?      2@             �\@                       @      @      K@      6@              $@      ,@              @      �?       @      K@             �Z@       @              �?      @     �O@     �E@       @      $@      "@       @                      @     �M@       @     @Z@       @       @      �?      @      D@      1@      �?      (@      @                               @      (@              G@      �?                       @      $@      @              @      @                               @      "@              D@      �?                              @      @               @                                              @              @                               @      @      @               @      @       @                      �?     �G@       @     �M@      �?       @      �?       @      >@      $@      �?       @      @       @                      �?      8@       @      G@      �?       @      �?       @      8@      @      �?       @                                              7@              *@                                      @      @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhM�9hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @n��Zt�?�	           ��@       	                   �0@�Fj���?�           ��@                           �?�P�'6�?k             e@                           @���m�.�?;            �W@������������������������       �^��I5v�?5            �T@������������������������       �"pc�
�?             &@                           @59���|�?0            �R@������������������������       �A�S���?$            �L@������������������������       � )O��?             2@
                           @�<��z��?u           @�@                           �?�!ݵݵ�?�           8�@������������������������       ��JH�.�?           x�@������������������������       �1��z���?�            �u@                           �?�-�C��?�           H�@������������������������       ��;���t�?�           ؃@������������������������       �$o���<�?�           ��@                           @��E��?�            �@                           �?0+e�?*           p�@                           �?v����?�            �u@������������������������       � �?���?�            0q@������������������������       ���Β��?/            @R@                          �2@���ï�?E            @������������������������       ��Cc}h,�?G             \@������������������������       �Fق!�>�?�             x@                           @��̵�?�             s@                           �?��<L��?u            @h@������������������������       ��.+K�j�?#            �H@������������������������       �����}��?R             b@                          �5@��>4և�?H             \@������������������������       ���#���?*            �O@������������������������       �?`[�?            �H@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �l@      A@      J@      7@     �U@     ��@     �B@     �@      8@       @     �S@      H@     Ѕ@     H�@      4@     �m@      g@      <@     �C@      0@     �P@     p{@      >@     X�@      4@      @     �P@     �G@     �|@     �y@      1@     �g@      (@               @              @     �C@      @      7@              �?      @       @      ;@     �A@              .@      @               @              @      4@      @      *@              �?              �?      (@      5@              $@      @               @              @      ,@      @      $@              �?              �?      (@      3@              $@                                              @              @                                               @                      @                                      3@              $@                      @      �?      .@      ,@              @       @                                      3@               @                      @      �?      (@      @              @      @                                                       @                                      @       @              �?     �e@      <@     �B@      0@     �N@      y@      ;@     ��@      4@      @     �N@     �F@     �z@     `w@      1@     �e@      T@      *@      =@      "@      B@     �f@      @     @u@       @      �?      7@      5@     `j@     �_@      "@     @R@     �M@      @      .@      @      >@     �`@       @      k@       @      �?      1@      2@      b@      X@      "@      K@      5@      @      ,@      @      @      I@       @     �^@                      @      @     �P@      >@              3@      W@      .@       @      @      9@      k@      7@      x@      (@      @      C@      8@     �k@      o@       @     @Y@     �I@      @      @      @      (@     �X@      0@     �a@      @       @      0@      (@     �X@      [@      @     �J@     �D@       @      @      @      *@     �]@      @     �n@      @       @      6@      (@     @^@     �a@      �?      H@     �G@      @      *@      @      5@     �g@      @     py@      @       @      (@      �?      n@      b@      @     �G@      C@      @      $@      @      *@      c@      @     �q@      @       @      @      �?     @f@     �Z@      @      C@      5@      @      @              @     �Q@      �?     �W@       @      �?      �?             �P@     �K@      �?      3@      2@              @              @      J@             �S@       @      �?      �?              I@     �F@      �?      0@      @      @                      �?      2@      �?      0@                                      1@      $@              @      1@              @      @      @     �T@      @      g@       @      �?      @      �?     �[@     �I@       @      3@       @              @       @       @      0@              =@                              �?      B@      .@              @      .@               @      @      @     �P@      @     �c@       @      �?      @             �R@      B@       @      *@      "@       @      @       @       @     �C@      �?     �_@                      @              O@      C@              "@      �?                              @      4@             �W@                      @              E@      9@              @      �?                                      @              .@                       @              0@      @              @                                      @      .@             �S@                      �?              :@      2@              �?       @       @      @       @      @      3@      �?     �@@                      @              4@      *@              @      @                       @      �?      @      �?      8@                      @              *@       @              �?      @       @      @               @      *@              "@                                      @      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��\_hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �<@ܐ+�N��?�	           ��@       	                     @��}���?	           t�@                            �?Rbվ�?�           ��@                           �?gv&��?b           ��@������������������������       ������?�            �w@������������������������       ��h^�K�?h           ��@                           �?Si�ma�?4           `�@������������������������       ���´t�?~           ��@������������������������       ��R|D�?�           �@
                           �?�����0�?�           ��@                          �;@�
���?l           ��@������������������������       ����6S�?]            �@������������������������       ��&%�ݒ�?             5@                           @.h��"�?           �{@������������������������       ��^M橍�?�             t@������������������������       ����f!�?M            �^@                           �?,'Zw��?�            �p@                           �? _����?F            �X@                           @��?,�?#            �H@������������������������       ����#E��?            �D@������������������������       �      �?              @                           @�u�)�?#            �H@������������������������       ��g�eX�?            �A@������������������������       �/����?             ,@                            �?��$2
�?w            �e@                          @@@�?�(ݾ�?E             Z@������������������������       �l�����?;             V@������������������������       �     ��?
             0@                           @�2y���?2            @Q@������������������������       �� B�~�?*             M@������������������������       ���!pc�?             &@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@     �@@      ?@      :@     �W@     ��@      ?@     ��@      5@      $@     @S@      K@      �@     ��@      8@     �n@      h@     �@@      =@      :@     @V@     p�@      <@     ��@      1@      "@     @Q@      K@     Ї@     �@      5@     �l@     @c@      ;@      6@      5@     @R@      |@      6@     h�@      1@       @     �K@      F@     �@     �x@      3@     �g@     �K@      (@      @      "@      3@     `f@      "@     �p@      @               @      $@     `h@     �_@       @     �@@      :@      @      @      @      (@     �R@      @     @T@       @              @       @     @T@     �K@       @      0@      =@       @      �?      @      @      Z@      @     �g@      @              �?       @     �\@      R@      @      1@     �X@      .@      2@      (@      K@     �p@      *@     �u@      (@       @     �G@      A@      t@     �p@      &@     �c@      B@      "@      $@      @      8@     �[@      �?     �Z@      @      �?      1@      (@     �^@      U@      @     �F@     �O@      @       @      @      >@     �c@      (@     �n@      @      @      >@      6@     �h@      g@       @     @\@      C@      @      @      @      0@     �e@      @     �t@              �?      ,@      $@     �n@     �\@       @     �C@      :@       @      @      @       @      W@      @     �h@              �?      @       @     �^@     �P@       @      4@      :@       @      @      @       @     �U@      @     �f@              �?      @       @     �^@     �P@       @      4@                                              @              .@                                      �?                              (@      @       @      �?       @     �T@      @     �`@                       @       @      _@      H@              3@      @      @       @              @     �J@       @     �Y@                      @      �?     �X@      @@              ,@      @                      �?      @      =@      �?      >@                      @      �?      :@      0@              @      (@               @              @      B@      @      \@      @      �?       @              E@      :@      @      1@       @               @              @       @              D@       @               @              @      0@      �?       @      @               @               @       @              ,@       @               @              @       @      �?      @      @               @               @       @              "@       @               @               @       @      �?      @                                                              @                                       @                      �?       @                               @                      :@                                      @      ,@               @       @                               @                      7@                                       @      @               @                                                              @                                      �?      $@                      @                              �?      <@      @      R@       @      �?      @             �A@      $@       @      "@      @                                      4@      �?      B@       @               @              9@       @              @      @                                      ,@      �?     �A@      �?               @              7@      @              @                                              @              �?      �?                               @      @              �?      �?                              �?       @       @      B@              �?      @              $@       @       @       @      �?                              �?      @       @      ;@              �?      @              "@       @       @       @                                              �?              "@                                      �?                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�:�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@���"%��?�	           ��@       	                     @*l���?�           D�@                           �?�]Z���?7           ��@                            �?&"mCy�?�           �@������������������������       �����(�?           ��@������������������������       �c�>�� �?�            pr@                           @��4��?b           8�@������������������������       ��3e���?�           h�@������������������������       �:KVE��?�           �@
                           �?���J�f�?{           ؎@                           @�v'8\�?            �|@������������������������       ����x6w�?�            �t@������������������������       �*h��5�?\             `@                          �9@K�Z�R`�?[           ��@������������������������       �L�ȱCW�?6           �}@������������������������       ����{�?%            �K@                           �?9��ǔ{�?           pz@                          @A@�>$*a�?k             d@                           �?�b�U5�?d            `b@������������������������       �Bf�����?8            @U@������������������������       ���A�9�?,             O@������������������������       �:/����?             ,@                           @r�l�w��?�            `p@                           @��y����?�            �k@������������������������       ���R��?|             h@������������������������       ���(\���?             >@                          �=@L�usr��?            �C@������������������������       ��ӭ�a��?             2@������������������������       �և���X�?             5@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@      <@     �F@      :@     �Z@     h�@      @@     $�@      .@      @      U@      J@     @�@     (�@      <@     p@      f@      8@      C@      9@     �W@      �@      @@     ��@      $@      @     �S@      I@     0�@     (�@      5@     @n@     �a@      (@      >@      5@     @T@     @{@      8@     ��@      "@       @     �P@      E@     `|@     �w@      4@     �g@      Q@      @      2@      *@     �H@     �i@      *@     �i@      @      �?      :@      :@     �l@     �d@      &@     �X@      M@              (@      *@     �@@     �d@      "@     �d@       @              2@      *@     `f@     @\@      @     �N@      $@      @      @              0@      D@      @     �D@      @      �?       @      *@      J@     �J@      @     �B@      R@      @      (@       @      @@     �l@      &@     Px@      @      �?      D@      0@     �k@     �j@      "@      W@     �@@      @      @      @      7@      Y@      @      i@      �?              $@      @     �\@      T@      �?     �C@     �C@      @      @      @      "@      `@       @     �g@       @      �?      >@      &@      [@     �`@       @     �J@     �B@      (@       @      @      *@     �a@       @     �t@      �?      �?      *@       @      l@      a@      �?      J@      7@      @      @       @      $@     @Q@      @     �_@      �?      �?      (@      @     �Y@     @P@              ;@      ,@      @      @       @      "@     �J@      @     �S@                      $@       @      U@      E@              7@      "@      �?                      �?      0@      @      H@      �?      �?       @       @      2@      7@              @      ,@      @      @       @      @     �Q@       @      i@                      �?      @     �^@      R@      �?      9@      ,@      @      @       @       @     �P@       @      g@                      �?      @     @Y@     �P@      �?      7@              @                      �?      @              1@                                      5@      @               @      0@      @      @      �?      (@     @S@             �e@      @      �?      @       @     �P@      @@      @      .@      $@      @      @              @      3@             �K@      @              @      �?      9@      .@      @      "@      "@      @      @              @      3@              J@      @              @      �?      6@       @      @      "@      @      @      @              @      ,@              ;@      @              @      �?       @       @      @      @      @              �?              �?      @              9@                                      ,@      @              @      �?                                                      @                                      @      @                      @                      �?      @      M@             �]@       @      �?       @      �?     �D@      1@      @      @      @                      �?      @     �J@             @V@       @      �?      �?      �?     �B@      1@      @      @      @                              @      D@              T@      �?      �?      �?      �?      ?@      1@      @      @                              �?              *@              "@      �?                              @                                                                      @              =@                      �?              @                                                                                      .@                      �?               @                                                                      @              ,@                                       @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?^[�Uȥ�?�	           ��@       	                    �?!��3�?Q           \�@                           �? ��IS�?n           ��@                            �?!�ҝ9�?�            �n@������������������������       �"sLj�'�?3            �T@������������������������       ��YJz��?h            �d@                          �:@�����4�?�             v@������������������������       ���� ���?�            `q@������������������������       ��˹�m��?.             S@
                            �?���b�?�           ��@                           @�� n��?�           (�@������������������������       ��,����?�            �x@������������������������       ��	C֣��?�            �o@                           @�n8R�F�?I           �@������������������������       � �R=���?F            @Z@������������������������       �� �s�E�?           y@                            @�b��?L           �@                          �;@��ϸ��?�           �@                          �0@��g���?R           p�@������������������������       ��P�!�c�?3            �V@������������������������       �EM���?           �@                           @6�����?m            �c@������������������������       �� ~�[g�?V             _@������������������������       ��� =[�?             A@                          �2@4�	va�?�           ��@                           �? #���?c            @f@������������������������       �-b�m?K�?"            �L@������������������������       �
��	�g�?A            @^@                          @@@F,����?*           `|@������������������������       �x ��"��?           �z@������������������������       ��p�F�:�?             7@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        k@     �B@      B@      :@     �Y@     ؅@      ?@     ��@      4@      .@     @U@     �L@     ��@     �@      1@     �p@     �\@      6@      ;@      ,@     �N@     �t@      (@     �y@      0@      @      =@      >@     �q@     �l@      "@     @b@      H@      @      2@      @      <@     �Y@             @c@      "@       @      *@      "@     �U@     �P@       @      J@      (@      @       @      �?      2@     �B@             �Q@      @              $@      @      :@      <@              9@      @               @      �?      @      $@              =@                      @      @      @      "@              $@      @      @      @              .@      ;@             �D@      @              @       @      3@      3@              .@      B@      @      $@       @      $@     �P@              U@      @       @      @      @      N@      C@       @      ;@      7@      �?      @       @      "@     �K@              O@      @       @      �?      @     �M@      ;@              4@      *@      @      @              �?      &@              6@                       @              �?      &@       @      @     �P@      .@      "@      &@     �@@      m@      (@     0p@      @      @      0@      5@      i@     �d@      @     �W@      E@      @      @      @      3@     �b@      @     `b@      @      �?      @      $@     �Z@     @U@      @      I@      6@      @       @      @      @     �X@      @     @T@      @              @      @     �Q@      K@      �?      <@      4@      @      �?       @      ,@      I@      �?     �P@      �?      �?              @      B@      ?@       @      6@      8@      "@      @      @      ,@      U@      @      \@       @      @      "@      &@     �W@     �S@      @      F@       @      �?                      @      8@      @      8@                      �?       @      $@      6@              @      0@       @      @      @      $@      N@      @      V@       @      @       @      "@      U@     �L@      @      C@     �Y@      .@      "@      (@      E@     �v@      3@     ��@      @      "@      L@      ;@     P{@     `q@       @     �^@     @U@      *@      "@      &@     �@@      p@      2@     {@      @      @     �I@      5@     �p@      j@       @      Z@     @T@      (@      "@      &@     �@@     �k@      ,@     �v@       @      @      H@      4@     �n@      i@      @     �X@      @                      �?              7@              (@                       @       @      1@      2@              $@      S@      (@      "@      $@     �@@      i@      ,@     �u@       @      @      G@      2@     �l@     �f@      @     @V@      @      �?                             �@@      @     @R@      �?              @      �?      8@      @       @      @      @      �?                              =@      @     �G@      �?               @              6@      @       @      @                                              @              :@                      �?      �?       @                              1@       @              �?      "@      [@      �?      l@      �?      @      @      @     �d@     �Q@              3@      "@                              @      ;@              G@                      @      @     �M@      5@              @      �?                                      �?              :@                                      2@      "@               @       @                              @      :@              4@                      @      @     �D@      (@              @       @       @              �?      @     @T@      �?     @f@      �?      @              @     �Z@     �H@              ,@      @       @              �?      @      T@      �?      e@      �?                      @      Y@     �H@              ,@      �?                               @      �?              "@              @                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ:�ThG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx         
                     @蒾6ˎ�?�	           ��@       	                    !@I$!3n��?�           �@                           �?��/���?�           Υ@                           @�uf\�p�?           ��@������������������������       �з��`{�?�           p�@������������������������       �06eg�w�?/            �Q@                           @(�ebu�?�           �@������������������������       ��hG/C��?�           ��@������������������������       ���7����?           �y@������������������������       �B{	�%��?             2@                          �;@s��\;0�?�           @�@                           �?�]��K�?g           ȍ@                           @�7�i�k�?           �y@������������������������       �`�;�ߐ�?�            `q@������������������������       ��&5D�?Y             a@                           @p�H��?\           ؀@������������������������       �XV<�?�            �m@������������������������       ���nʠ��?�            �r@                           �?(-A#��?e            �b@                           �?��S�r
�?             <@������������������������       �0�����?             5@������������������������       �����>4�?             @                           @.u�m���?R            �^@������������������������       ��>4և��?             <@������������������������       ��[`��>�?A            �W@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@      D@      >@      7@     �W@     ��@      8@     Ԑ@      ;@      $@     �U@     �Q@     ��@     (�@      6@      n@      c@      @@      9@      4@     �R@     �~@      1@     ��@      6@      @      R@     @P@     ��@      x@      4@     �h@     �b@      @@      9@      4@      R@     P~@      (@     ��@      6@      @      R@     @P@     ��@      x@      4@     �h@     �P@      &@      0@      @      G@     @m@       @     pp@      5@      @      ?@      A@     �l@     �c@      &@     �[@      P@      &@      .@      @     �F@     �l@       @      n@      2@      @      ?@      A@     �j@     �b@      &@     �X@       @              �?              �?      @              6@      @                              1@      @              *@     @U@      5@      "@      *@      :@     `o@      @     �z@      �?      �?     �D@      ?@     0s@     `l@      "@     �U@     @S@      &@       @      &@      3@      i@      @     Pr@              �?      :@      7@     �l@     @c@       @      P@       @      $@      �?       @      @      I@      �?     �`@      �?              .@       @     @S@     @R@      �?      6@      �?                               @      @      @      �?                                               @                     �H@       @      @      @      5@      i@      @     x@      @      @      .@      @     �k@     ``@       @      F@      F@       @       @      @      1@     �d@      @     0t@       @              .@      @     �h@      _@      �?      D@      8@       @       @              .@     �T@      @     �[@      �?              &@      �?     �S@     �M@              2@      6@      @       @              "@     �P@      �?      O@      �?              @      �?     �H@     �D@              .@       @      @                      @      0@      @      H@                      @              >@      2@              @      4@                      @       @      U@      @     �j@      �?              @      @     �]@     @P@      �?      6@      &@                      @              6@             �Z@                       @      �?     �L@      4@              0@      "@                               @      O@      @     �Z@      �?               @       @     �N@     �F@      �?      @      @              @              @      A@              O@      @      @              �?      8@      @      �?      @                                              �?              1@                              �?      @      �?              �?                                              �?              .@                              �?      @                                                                                       @                                      @      �?              �?      @              @              @     �@@             �F@      @      @                      1@      @      �?      @      �?              @              @      @               @      �?      @                      @      �?                      @                              �?      >@             �B@       @                              (@      @      �?      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?���G��?�	           ��@       	                     @p��%CD�?/           ��@                           @�`�!x�?           X�@                           @�
t�d�?�           ��@������������������������       ���"��?x           ��@������������������������       ������C�?�            �l@                          �4@�׬]l�?           �y@������������������������       ���"$�c�?k            �e@������������������������       ��0��#�?�            �m@
                           �?��	����?,           0}@                          �9@SPt֭�?i            �d@������������������������       �h�"�`��?Y            �a@������������������������       ��q�q�?             8@                           @#�n��Q�?�            �r@������������������������       ������?�            �i@������������������������       ��IBD�A�?=            �W@                           �?������?z           @�@                           @��SP��?�            �u@                          �4@�X�s�V�?a            �c@������������������������       ��-YS��?-            @R@������������������������       ���l���?4             U@                          �;@�s)m<��?{            �g@������������������������       ��Q��{�?j             d@������������������������       �f?����?             ?@                          �;@���!X��?�           �@                           @Җ�����?           ��@������������������������       �c��� ��?'           ��@������������������������       �b�I�1��?�           �@                           @`Cl��?�            @l@������������������������       �UUUUUU�?{             h@������������������������       �8�
t�F�?             A@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      :@      G@      <@     @[@     �@      <@     ��@      3@      &@     �R@      N@     ��@     ��@      5@     �p@     �Z@      4@      =@      *@      Q@     pr@      ,@     �x@      ,@      @      ?@      =@      s@     �l@      @     �a@     �R@      (@      8@      *@     �L@     @k@      $@     pp@       @      @      8@      9@     �k@     `e@      @     @Z@      J@      @      0@      *@      H@      a@      @     �g@      @      @      0@      *@     �c@     �X@      @     �P@     �C@      @      ,@      *@     �D@     @Y@      @      `@      @      @      *@      &@      Y@     @R@       @     �H@      *@      �?       @              @     �A@      �?      N@               @      @       @     �L@      :@      �?      2@      7@      @       @              "@     �T@      @     �R@      @      �?       @      (@      P@      R@      @      C@       @      @       @              �?     �D@      @      >@              �?      @      @      1@      @@      @      &@      .@                               @     �D@      @     �F@      @              �?      @     �G@      D@              ;@      ?@       @      @              &@     @S@      @     �`@      @              @      @     �T@      M@      �?     �B@      &@      @      �?              @      @@      @     �D@                      @       @      B@      ,@              ,@      $@      @      �?              @      =@      @     �@@                      @              :@      ,@              ,@      �?                                      @               @                               @      $@                              4@      @      @               @     �F@      �?     �W@      @              �?       @     �G@      F@      �?      7@      4@       @      @              @      >@      �?     �K@      @              �?       @     �@@     �A@      �?      ,@              @                      @      .@             �C@                                      ,@      "@              "@     �X@      @      1@      .@     �D@     `u@      ,@     ��@      @      @      F@      ?@     0z@      s@      ,@     �_@      4@              @      @      "@      H@      @      W@                      @       @     �P@     �M@       @      @@      "@               @      @       @      ;@              @@                       @       @     �E@      *@              6@      @                                      @              (@                      �?              >@      @              .@      @               @      @       @      6@              4@                      �?       @      *@      @              @      &@              @      �?      @      5@      @      N@                      @              7@      G@       @      $@      &@              @      �?      @      0@      @     �E@                      @              4@      D@       @      $@                                              @              1@                                      @      @                     �S@      @      (@      &@      @@     `r@      &@     Ѓ@      @      @      C@      =@     v@     �n@      (@     �W@     �R@      @      (@      $@      @@      o@      $@     ؀@       @      @     �A@      :@     @s@      m@      @     @V@     �F@       @      @      @      *@     �_@      @     `q@      �?              1@      (@      h@     @]@      @     �B@      =@      @      @      @      3@     @^@      @     Pp@      �?      @      2@      ,@      ]@      ]@      @      J@      @                      �?              G@      �?     �W@      @       @      @      @     �F@      (@      @      @      @                      �?             �D@      �?      R@      @       @       @      @      E@      $@      @      @                                              @              7@                      �?              @       @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�AmhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@3�Q���?�	           ��@       	                     @�s�M��?�           L�@                            �?N��� �?<           ģ@                           �?��6��?�           ��@������������������������       �T���l��?	           0�@������������������������       �$�6S#�?�           �@                           �?�M<T��?�           ��@������������������������       ��k\���?�            @m@������������������������       �n�5�?           �|@
                          �2@x�b.d�?l            �@                           �?7�\�~��?�            �q@������������������������       �l�����?Z            �`@������������������������       �ʮ��?Z            �b@                           �?x���1�?�           H�@������������������������       �r07W�A�?�            �p@������������������������       �^�*��?           �y@                            �?~ln)k~�?           0z@                            �?�5���?�             l@                           �?�Z�k%�?P            �[@������������������������       �����K�?             2@������������������������       ��@#U�?E            @W@                           �?p+>[��?I            �\@������������������������       �Y�����?             F@������������������������       ��݃�R��?.            �Q@                           �?Yy�o���?}            @h@                          �?@�kWw��?:            �V@������������������������       �^�VCr�?/            �Q@������������������������       �r`�����?             3@                            @�t���]�?C             Z@������������������������       ��η���?             ?@������������������������       �*�l�Ø�?/            @R@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        l@      :@      8@      4@     @Z@     `�@     �B@     <�@      0@      *@      U@      R@     @�@     �~@      5@     `o@     �h@      6@      6@      4@     �X@     H�@      A@     �@      $@      *@      S@      Q@      �@     0}@      2@     @l@      d@      1@      0@      3@     �U@     �|@      9@     ��@      "@      (@      O@     �K@     �|@     `u@      2@     �g@      \@      (@      "@      *@     �H@     v@      1@     �~@      @      @      ?@      >@     @v@     �k@       @      _@     �J@      @      @      @      ?@      f@      @     �f@      @      @      (@      .@     �b@     @V@      @      N@     �M@      @      @      @      2@      f@      &@     0s@                      3@      .@     �i@     �`@      @      P@     �H@      @      @      @     �B@      [@       @     @Z@      @      @      ?@      9@     �Z@     �]@      $@     �P@      2@      @      @      @      &@      =@       @      9@      @              @      .@      G@     �H@       @      2@      ?@       @      @      @      :@     �S@      @      T@      �?      @      :@      $@     �N@     �Q@       @      H@      C@      @      @      �?      *@     �c@      "@     u@      �?      �?      ,@      *@      j@     @_@              B@      @      �?              �?      @     �C@       @     �W@                      @      @      T@      @@              .@       @                      �?      @      7@             �H@                      @      @      ;@      ,@              "@      @      �?                              0@       @     �F@                       @      �?     �J@      2@              @      ?@      @      @              $@     @]@      @     `n@      �?      �?      "@      "@      `@     @W@              5@      0@      @      �?              @     �H@      @      Q@              �?       @      �?     �K@     �I@              @      .@      �?      @              @      Q@       @     �e@      �?              �?       @     �R@      E@              ,@      9@      @       @              @     �P@      @     �e@      @               @      @      R@      6@      @      9@      @      @      �?              @     �F@      �?     @U@       @               @      �?     �D@      ,@              *@      @                               @      .@      �?     �I@       @              @              6@      @              @                                               @              @                      @              @                       @      @                               @      *@      �?      G@       @              �?              0@      @               @      @      @      �?              �?      >@              A@                      @      �?      3@      @              "@       @                                      @              ,@                      @      �?       @      @              @       @      @      �?              �?      7@              4@                      �?              &@      @              @      2@              �?              @      6@       @     �U@      @                      @      ?@       @      @      (@      *@              �?              @      @             �D@       @                       @      "@      @              @      @              �?              @      @              B@                               @      "@      @               @       @                                                      @       @                                      �?              @      @                                      .@       @      G@       @                      �?      6@      �?      @      @      @                                      @       @       @                              �?      @              @      @      �?                                      &@              C@       @                              2@      �?               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJW�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @��d؉��?�	           ��@       	                    @�������?�           ĥ@                           @��Ռ �?%           *�@                            �?(��O �?�           `�@������������������������       �ݴ׊Od�?�           ��@������������������������       ����r|�?Q           8�@                          �5@	�}Mh�?G           �@������������������������       ��1��>b�?�            �s@������������������������       ����c�?v            �g@
                          �;@h.���?�           h�@                            �?`� �?�           ��@������������������������       �7�w[��?3           �}@������������������������       ���FA6�?`             c@                           �?
�-6�?;            @V@������������������������       �騷}*_�?             ;@������������������������       ��AI-���?(             O@                          �;@;0b�@�?�           ��@                           �?<%�3~q�?o           ��@                           �?Y�X*�q�?           �z@������������������������       �l(�����?e             c@������������������������       �FP��.�?�            q@                          �2@�(��m�?Z           X�@������������������������       �|��
�?d             d@������������������������       �E4� )��?�            �x@                          �=@��`]���?]            `b@                           @*�o\��?+             O@������������������������       ��^�q��?            �@@������������������������       ��CE5��?             =@                           �??c�����?2            @U@������������������������       �:/����?             <@������������������������       ���a0��?!            �L@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      <@     �G@      7@     �X@     ��@      :@     �@      4@      "@      T@     @P@     �@     ��@      1@      p@     �f@      0@     �B@      3@     �S@      |@      5@     0�@      *@      @      R@      L@     �@     px@      0@     �j@      c@      &@      A@      1@     �P@     Pu@      (@     ��@      @       @      K@      E@     w@     0p@      $@     @c@      ]@      &@      7@      *@      H@      q@      "@     �w@      @             �D@      C@     �q@     `i@       @     �\@      J@      @      @      @      ,@      ]@      @      f@      �?              (@      .@     @_@     �O@       @     �@@      P@       @      4@      @      A@     �c@      @     @i@       @              =@      7@     `c@     �a@      @     �T@      B@              &@      @      2@     �P@      @     @d@      @       @      *@      @     @V@      L@       @     �C@      5@               @      @      *@      J@       @     @Z@       @       @      *@      @      @@     �D@              5@      .@              @      �?      @      .@      �?     �L@      �?                      �?     �L@      .@       @      2@      =@      @      @       @      *@     @[@      "@     @e@      @      �?      2@      ,@     �a@     �`@      @     �M@      <@      @      @       @      *@     @Y@      "@      `@      @      �?      2@      (@      ]@     �^@      @     �K@      8@      @      @       @      (@     �T@       @      Z@       @      �?      $@      @     �X@     �T@       @      A@      @       @                      �?      3@      �?      9@      @               @      @      2@      D@      @      5@      �?                                       @             �D@                               @      8@      "@              @      �?                                      @               @                                      @      @              @                                              @             �@@                               @      2@      @                     �C@      (@      $@      @      3@     �i@      @      x@      @      @       @      "@     �l@     �a@      �?     �E@      >@      (@      $@      @      1@     `f@      @     �s@       @      @       @      @      j@     @a@      �?      D@      &@       @      @      �?      0@     �T@      @     @\@      �?      @      @      @      S@     �Q@              6@      @      @       @               @     �@@       @      @@                      @              A@      6@              &@      @      @      @      �?      ,@     �H@      @     @T@      �?      @      �?      @      E@     �H@              &@      3@      @      @      @      �?     @X@             @i@      �?              @      @     �`@     �P@      �?      2@      @               @      @              ;@              F@                      �?             �G@      :@               @      0@      @      �?              �?     �Q@             �c@      �?               @      @     @U@     �D@      �?      $@      "@                               @      <@             @Q@      @       @               @      6@      @              @       @                                      0@              A@                                      @      @               @      �?                                      @              4@                                       @      @              �?      �?                                      &@              ,@                                      �?      �?              �?      @                               @      (@             �A@      @       @               @      3@                      �?      @                                       @              @       @                       @      $@                      �?       @                               @      $@              =@      @       @                      "@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�P_hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @A3��r��?�	           ��@                            �?�c$�	�?�           �@                           !@���t��?N           ��@                           �?k&_��?D           ��@������������������������       ������?[           ��@������������������������       ��ܯ���?�           8�@������������������������       �>
ףp=�?
             4@                          �;@0�!8���?�           ��@	       
                   �4@J�J��?�           �@������������������������       �����m��?�            pu@������������������������       ���(x]��?�            �p@                           �?���.�?&            �L@������������������������       �窷uJ��?             3@������������������������       �D�n�3�?             C@                           �?$s0��?�           P�@                          �;@��:�a�?�            �t@                          �8@Q�=.�?�            `r@������������������������       �-���?�            �o@������������������������       �1��D�\�?            �C@                           �?Z;����?             A@������������������������       �R���Q�?             4@������������������������       ��X�C�?             ,@                           @4p6�֜�?�           `�@                           @O�D^���?�           �@������������������������       �W)#���?�           ��@������������������������       �
ц�s�?	             *@                          �3@^Ƒڋ��?B            @Z@������������������������       ���d�T��?            �D@������������������������       �     ��?'             P@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@      >@     �C@      0@     @_@     h�@      A@     @�@      0@      "@     �R@     �K@     ��@     �@      ,@     �p@      f@      9@      ?@      *@     �X@      @      ;@     ��@      &@      @     �O@      G@     �~@     `w@      &@     @m@      a@      1@      3@      *@     �O@     �y@      4@     �@      @      �?     �G@      ;@     �x@     �o@      @      c@     �`@      1@      3@      *@     �N@     y@      1@     ��@      @      �?     �G@      ;@     �x@     �o@      @      c@      R@      @      0@      @     �E@     �g@       @     `l@      @      �?      7@      (@     `d@     �W@      @     @T@     �O@      $@      @      @      2@     @j@      "@     �u@       @              8@      .@     �l@     �c@      �?     �Q@       @                               @      $@      @      �?                                               @                     �C@       @      (@              B@     �U@      @     �^@      @      @      0@      3@      Y@      ^@      @     �T@      B@       @      (@              B@     �T@      @      X@      @      @      .@      3@     @V@      ]@      @      T@      4@      @      @              1@      I@      �?     �H@              @      &@      0@      B@      P@      @      N@      0@      @      @              3@     �@@      @     �G@      @      @      @      @     �J@      J@              4@      @                                      @       @      ;@                      �?              &@      @      @       @                                               @       @      @                                              @      @       @      @                                       @              4@                      �?              &@      �?                     �B@      @       @      @      :@     `g@      @     �y@      @       @      (@      "@      m@     @`@      @     �@@      @               @      �?      @      K@      �?      [@                      @      @     �S@     �G@              3@      @               @      �?       @      I@      �?     @V@                      @      �?      S@     �E@              1@      @               @      �?       @     �D@      �?     �U@                      @      �?      O@     �A@              .@      @                                      "@              @                                      ,@       @               @                                      �?      @              3@                               @       @      @               @                                              @              &@                               @       @      �?                                                      �?                       @                                              @               @      >@      @      @       @      7@     �`@      @     �r@      @       @      @      @     `c@     �T@      @      ,@      =@      @      @       @      5@     �\@      @     �o@      @       @      @      @     @`@      T@      @      *@      =@      @      @       @      5@      [@      @     @o@      @       @      @      @     �_@      T@      @      *@                                              @              @                                      @                              �?       @      �?               @      3@       @      G@       @              �?              9@      @              �?                                               @       @      9@                      �?              @      �?              �?      �?       @      �?               @      &@              5@       @                              6@       @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ �hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?���w�?�	           ��@       	                   �:@�\`�]�?C           �@                            @����0�?�           ��@                            �?	�n�7��?�           ��@������������������������       ���8���?�             x@������������������������       ���)���?�           h�@                           @������?            y@������������������������       �|�E��?�            p@������������������������       ��|�H�?W            �a@
                           @j�[�v�?�            pp@                            �?h`z\��?�            �l@������������������������       �b���i��?,            �P@������������������������       �y�v�J�?f            �d@������������������������       �     P�?             @@                           @�B�����?b           
�@                          �4@��Z�Ai�?I           ��@                           @�\��/��?           `{@������������������������       ���x�6L�?�             u@������������������������       ��~�:p��?<             Y@                           @�.�?� �?*            ~@������������������������       ��D���?           �y@������������������������       �Lh/����?)             R@                          �<@<��5��?           ��@                           !@�,�¦_�?�           ��@������������������������       ������c�?�           h�@������������������������       ��g���e�?             &@                            �?�T�[j�?T            @a@������������������������       �l�����?             F@������������������������       �x���T��?:            �W@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      7@      K@      2@     �]@     ��@     �@@     ��@      7@      "@      Q@     �N@     �@     �@      1@     �p@     �X@      (@     �C@      $@      R@     �r@      3@      |@      *@      @      @@      7@      r@     �l@       @     �`@      U@      $@     �@@      $@     �P@     pq@      1@     0v@      "@      @      :@      7@     �l@      i@      @      \@      P@      @      :@      "@     �L@     �i@      *@     �l@       @      @      3@      6@     �c@     �b@      @     @W@      2@       @      @      @      *@     �Q@      @      [@      �?              "@      "@     �N@     �L@      @      2@      G@      @      4@      @      F@      a@      @     �^@      @      @      $@      *@     �W@     �V@      @     �R@      4@      @      @      �?      "@     @R@      @      _@      �?      @      @      �?     �R@     �J@              3@      *@      @      @      �?      @     �H@             �Q@                      @             �M@     �@@              (@      @              @              @      8@      @      K@      �?      @              �?      0@      4@              @      .@       @      @              @      4@       @     @W@      @              @             �M@      =@      �?      4@      .@       @      @              @      0@       @      S@      @              @             �I@      ;@      �?      3@                                      @      $@       @      @@                      �?               @      @              @      .@       @      @              @      @              F@      @              @             �E@      8@      �?      (@                                              @              1@                                       @       @              �?     �V@      &@      .@       @      G@     �t@      ,@     0�@      $@      @      B@      C@      ~@     @q@      "@      a@     �G@      @       @       @      5@     @[@       @     `r@      @       @       @      *@     �n@     �X@      @     �K@      8@              @       @      @     �P@             @]@                      @      @     ``@     �E@      @      >@      7@              �?      �?      @      M@             @S@                      @       @     �[@     �A@              7@      �?              @      �?      @      "@              D@                              @      4@       @      @      @      7@      @      @              ,@      E@       @      f@      @       @      @      @     @\@     �K@       @      9@      7@      @      @               @      A@       @      c@               @      @      @      V@     �K@       @      7@                                      @       @              9@      @                       @      9@                       @      F@      @      @      @      9@     �k@      (@      x@      @      �?      <@      9@     �m@     @f@      @     @T@      F@      @      @      @      9@      h@      &@      t@      @      �?      9@      6@     @j@     �e@      @     �R@      F@      @      @      @      9@      g@      &@     �s@      @      �?      9@      6@      j@     �e@      @     �R@                                              @              @                                      �?                                                                      =@      �?      P@                      @      @      :@      @              @                                              @              8@                              @      @      @                                                              8@      �?      D@                      @              3@      �?              @�t�bub��     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?8�s���?�	           ��@       	                     @VE�0�?]           `�@                            �?+R��	��?           ��@                           �?k�!w��?           z@������������������������       �Ҙ_&��?n            @e@������������������������       ��u�x�8�?�            �n@                           �?6�{>��?           p�@������������������������       �-�����?g            �d@������������������������       ��������?�           @�@
                           @`�0y���?>           �~@                           �?qgsz? �?           Py@������������������������       ���?N�0�?�            @o@������������������������       ��ql���?\            `c@                          �4@�u]�u]�?8             U@������������������������       �4�%�p�?             �I@������������������������       �ܛ)��	�?            �@@                            @��p���?c           �@                          �0@���t�H�?�           ��@                           @�\/�@g�?4            �T@������������������������       ��v:���?             A@������������������������       �r�q��?             H@                          �1@��^p�,�?�           p�@������������������������       �H$�QR�?k            `f@������������������������       �x����2�?P           ��@                           @X�����?t           �@                          �2@��"ñ��?           �z@������������������������       ��\Fs��?K            �\@������������������������       �͓!g���?�            �s@                           �?��N&�g�?a            �b@������������������������       ���_�L�?             9@������������������������       ��!wI2�?T            �_@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      <@      H@      =@     �X@     8�@      D@     ��@      2@      @     @T@     �Q@     Ȇ@     ��@      ,@     `o@      Y@      .@     �A@      .@     �N@     t@      4@     py@      (@      @      <@     �A@      s@      o@      @     �a@      S@      "@      =@      *@      I@     �k@      ,@     @p@      $@      @      5@      @@     �i@      h@      @     @^@      2@      �?       @       @      1@     @U@      @     @Z@      �?              @       @      Q@     �O@      �?      C@      @      �?       @      �?      @      4@      �?     �F@                      @      @      <@      >@              8@      *@                      �?      $@     @P@      @      N@      �?              �?      @      D@     �@@      �?      ,@      M@       @      ;@      &@     �@@      a@      $@     `c@      "@      @      1@      8@      a@      `@      @     �T@       @       @      ,@      @      "@      E@              1@      @              @      �?      3@      1@              7@      I@      @      *@      @      8@     �W@      $@     @a@      @      @      &@      7@     �]@      \@      @      N@      8@      @      @       @      &@     �X@      @     `b@       @              @      @     @Y@      L@              3@      7@      @      @              $@     @U@      @     @[@       @              @      @     �U@     �H@              1@      2@      @      @              @     �I@       @      Q@       @              @              I@      A@              @      @       @                      @      A@       @     �D@                      �?      @     �B@      .@              $@      �?      �?               @      �?      ,@       @      C@                       @              ,@      @               @      �?                       @      �?      *@       @      8@                       @              @      @                              �?                              �?              ,@                                      &@      @               @     @X@      *@      *@      ,@      C@     `t@      4@     h�@      @             �J@      B@     pz@     �q@       @     �[@     �S@      (@       @      *@     �@@     �l@      1@     @~@      @             �H@      >@      s@     @k@      @     �X@      @                      �?              9@              (@                      @       @      *@      $@              "@       @                                      1@              �?                       @       @       @       @                      @                      �?               @              &@                       @              @       @              "@      R@      (@       @      (@     �@@     `i@      1@     �}@      @             �F@      <@     0r@      j@      @     @V@      0@               @                      8@      @     �P@                      @      @      0@     �@@              $@      L@      (@      @      (@     �@@     `f@      *@     `y@      @              D@      9@     0q@     �e@      @     �S@      3@      �?      @      �?      @     �X@      @      m@       @              @      @     �]@      Q@       @      *@      1@              @      �?      @      L@      @     �g@       @               @      @     �T@      I@              (@      @              �?              �?       @             �J@                              �?      A@      "@               @      (@              @      �?      @      H@      @      a@       @               @      @      H@     �D@              $@       @      �?                              E@              F@                       @       @     �B@      2@       @      �?                                              "@               @                                               @                       @      �?                             �@@              B@                       @       @     �B@      $@       @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJL�6hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �6@�}_"��?�	           ��@       	                     @��
���?Z           ��@                           �?��6q�5�?�           $�@                           @�0����?<           ��@������������������������       �Ubږ���?�           p�@������������������������       ��ES0�3�?�            �h@                          �0@�F��ɩ�?w           ��@������������������������       �DSbq���?,             Q@������������������������       �Q_��?K           ��@
                           �?B{�}�?�           ��@                           �?�r��dn�?�            �r@������������������������       �^��$8�?P            �^@������������������������       ��ȓ�)��?~            �f@                           �?W�7�L\�?�             u@������������������������       �x�߿��?�             i@������������������������       ���d�!�?V            �`@                           �?�Ɨ7���?x           �@                            �?��`+
��?�            �t@                          �9@��M��?<            @W@������������������������       ��-�����?!             G@������������������������       ��{T�H�?            �G@                           @��:m��?�             n@������������������������       ������;�?i            �a@������������������������       ���z����??            @X@                            @(�wd�?�           А@                           �?���0`�?�           І@������������������������       �pN�,m�?K            �]@������������������������       ��2-H
��?v           �@                          �@@[ٵ�|N�?�            �u@������������������������       ��$nҢ��?�            �t@������������������������       �޾�z�<�?             *@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@      C@     �C@      <@     �Y@     ��@      G@     (�@      &@      (@      T@     �L@     �@      @      ,@     �q@     @d@      6@      ;@      5@     �R@     �y@      @@     �@      @      "@      K@     �D@     @|@     Ps@      $@     �h@     �_@      0@      9@      ,@      N@      t@      7@      }@      @      @      H@     �B@     �r@     �n@      $@     �d@      O@      *@      5@      @      B@     `c@      ,@     `g@       @      @      :@      0@     ``@     �]@      @     �U@     �H@       @      .@      @     �A@      [@      "@     �b@              @      9@      $@      Z@     @U@      @      S@      *@      @      @              �?     �G@      @     �B@       @       @      �?      @      ;@     �@@      �?      &@     @P@      @      @      "@      8@     �d@      "@     Pq@      �?      �?      6@      5@     �d@      `@      @      T@      @                       @              1@              "@                              @      .@      "@              "@      O@      @      @      @      8@     �b@      "@     �p@      �?      �?      6@      1@     �b@      ^@      @     �Q@     �A@      @       @      @      .@     �V@      "@     @j@       @      @      @      @     �c@      O@              @@      .@      @      �?      �?      *@     �I@      @      U@              @      @       @     �P@     �@@              4@      @      �?                      @      :@      @      4@                      @             �B@      @              &@       @      @      �?      �?      @      9@      �?      P@              @      �?       @      =@      :@              "@      4@       @      �?      @       @     �C@      @     �_@       @              �?       @     �V@      =@              (@      "@              �?      @              7@      @     �R@       @              �?       @     �F@      7@              $@      &@       @                       @      0@             �I@                                     �F@      @               @     �J@      0@      (@      @      <@     �j@      ,@     �z@      @      @      :@      0@     �s@     `g@      @     �T@      6@      @      �?      @      @     �F@      �?     �Q@      �?              &@      @      T@      L@      �?      9@      @                       @       @      &@              4@                       @      @      @@      @               @      @                              �?      $@              $@                      �?      @      "@      @              �?      �?                       @      �?      �?              $@                      �?              7@      �?              @      0@      @      �?      @       @      A@      �?     �I@      �?              "@      @      H@      I@      �?      1@      $@      @              @              ,@              E@                      @       @      :@      =@      �?      @      @              �?               @      4@      �?      "@      �?               @      �?      6@      5@              &@      ?@      *@      &@       @      8@      e@      *@     v@      @      @      .@      "@     �m@     ``@      @     �L@      0@      $@      @       @      0@      ]@      &@     `k@       @              .@      @     @c@      Z@       @      I@      @       @              �?      @      "@      �?      F@                      �?      @      3@      .@              0@      &@       @      @      �?      *@     �Z@      $@     �e@       @              ,@      @     �`@     @V@       @      A@      .@      @      @               @     �J@       @     �`@      @      @               @     �T@      ;@      �?      @      *@      @      @               @     �J@       @      _@      @      @               @     �T@      ;@      �?      @       @                                                      $@                                      �?                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ.COdhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@�F�' I�?�	           ��@       	                    �?�I��h�?�           ��@                            @�&�����?2           �|@                          �2@%e�*���?�            �s@������������������������       �9��8���??             X@������������������������       �B�P���?�             k@                          �6@9���d<�?b            �b@������������������������       �_1"g.��?E            �Y@������������������������       �#�tV�?            �G@
                            @6UorSP�?R           "�@                           @�L���?W           �@������������������������       ����A�?W           ��@������������������������       ���^5��?            �@                           �?��4�^��?�           �@������������������������       ��]���)�?�            �u@������������������������       �;�J�>�?            �|@                           @d��ϼ�?(           �~@                           @h�k:<q�?           �z@                           @hCG���?�            �u@������������������������       �7@�%��?�            pq@������������������������       ����F�?.            @Q@                            �?G[����?,            @S@������������������������       ��Q����?             D@������������������������       ��fj��?            �B@                          �<@      �?'             P@                            �?�?�(ݾ�?             :@������������������������       �*L�9��?             &@������������������������       �z�G�z�?	             .@                           �?�S����?             C@������������������������       �N��)x9�?
             ,@������������������������       ��q�q�?             8@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@     �C@     �G@      6@     @T@     ��@      :@     8�@      2@      &@     �P@      L@      �@     P�@      ,@     �n@     �e@      ?@      D@      4@      R@     h�@      7@     (�@      (@      $@      K@     �K@     Ȅ@     @~@      &@     �k@      ?@      �?       @      �?      (@     �H@       @     @_@      @              "@      @     �T@     �T@      �?      I@      5@      �?      @      �?      $@      8@       @     �S@      @               @      @      O@      F@      �?     �G@      ,@              @              �?       @      �?      >@      @              @       @      *@       @      �?      "@      @      �?      �?      �?      "@      0@      �?     �H@      @              @      �?     �H@      B@              C@      $@              @               @      9@              G@                      �?              5@      C@              @      $@              @               @      5@              ?@                      �?              *@      3@              @                      �?                      @              .@                                       @      3@                     �a@      >@      @@      3@      N@     ��@      5@     @�@      @      $@     �F@      J@     0�@      y@      $@     `e@     @\@      1@      8@      *@     �J@     �y@      3@     @�@      @      "@      D@      H@     px@     �s@      $@     �a@     �O@      @      &@      &@      :@     `g@      @     Pp@      �?              $@      (@     @i@     @Y@      @      J@      I@      &@      *@       @      ;@     @l@      .@     0r@      @      "@      >@      B@     �g@     `j@      @     �V@      <@      *@       @      @      @     �_@       @      r@       @      �?      @      @     �g@     �V@              =@      ,@       @       @      �?      @      N@       @     @W@              �?      @      �?     @T@      G@              4@      ,@      @              @      �?     �P@             `h@       @              �?      @     �[@      F@              "@      <@       @      @       @      "@     �R@      @      i@      @      �?      (@      �?     �Q@      C@      @      8@      <@       @      @       @      "@     �P@      @      d@      @      �?      "@      �?     �N@     �B@      @      7@      9@       @      @       @      "@     �H@      @     �`@      @      �?      "@      �?      J@      3@      @      5@      8@       @      @       @      @     �E@      @      Z@      @      �?      �?      �?      D@      2@      �?      ,@      �?                              @      @              =@                       @              (@      �?       @      @      @                                      1@              <@                                      "@      2@               @                                              @              4@                                      @      &@              �?      @                                      *@               @                                      @      @              �?                                              "@              D@                      @              $@      �?              �?                                              @              0@                      @               @      �?              �?                                                              @                      @               @      �?              �?                                              @              (@                                                                                                              @              8@                                       @                                                                      @              @                                      @                                                                      �?              4@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?���`���?�	           ��@                          �0@�UY64�?-           ܚ@                            @�|a2U�?=             Y@                            �?EQEQ�?5             U@������������������������       ��렵0�?%            �N@������������������������       �`������?             7@������������������������       �     ��?             0@                           �?���,�?�           L�@	       
                     @����[�?S           �@������������������������       ��l��?�            �r@������������������������       �ѧ�I� �?�             o@                           @��L���?�           Ȑ@������������������������       ����Z2D�?           �z@������������������������       ����aSG�?�           @�@                            @BhI����?[           $�@                            �?b5�$9r�?�           ��@                           @GAr���?�           p�@������������������������       ���1>�?�           p�@������������������������       �Ic�2�?'           �~@                           @rE�6���?�            `x@������������������������       �NwR����?\            �b@������������������������       ��`6�:C�?�            @n@                           �?�^��Կ�?�           ��@                           �?z���}��?�            �y@������������������������       ��x���?=            �W@������������������������       ��H5~�?�            �s@                           @rw2'�$�?�            �j@������������������������       �/��N�^�?7            @V@������������������������       �0��Q�(�?V            @_@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �f@     �C@     �D@      8@     @X@     8�@      A@     �@      1@      @      R@      N@     (�@     ��@      3@     q@     @V@      7@      9@      .@      P@      u@      8@     �y@      (@      @      =@      ?@     �p@      l@      $@     �b@      @      @      �?      �?      "@       @      @      0@      �?      �?       @      @      ,@      0@      �?      .@       @      @      �?      �?       @       @      @      ,@      �?      �?              @      ,@      &@      �?      &@      �?              �?      �?       @      @      @       @      �?                      @      "@      "@              "@      �?      @                               @              @              �?                      @       @      �?       @      �?                              �?              �?       @                       @                      @              @     �U@      4@      8@      ,@     �K@     �t@      3@     �x@      &@      @      ;@      ;@     p@      j@      "@     �`@      ;@      "@      *@       @      1@     @X@      @     `b@       @              &@      @      R@      Q@      @      L@      ,@      @      $@       @      "@     �F@      @      R@      @              @       @      ;@      C@       @     �G@      *@      @      @               @      J@      �?     �R@      �?              @       @     �F@      >@       @      "@     �M@      &@      &@      @      C@      m@      .@     �n@      @      @      0@      7@      g@     �a@      @     �S@      7@      @      @      �?      &@     @]@      $@      V@      �?              @       @      U@     �I@       @      9@      B@      @       @      @      ;@      ]@      @     �c@       @      @      (@      5@     @Y@     @V@      @      K@     @W@      0@      0@      "@     �@@     Pw@      $@     x�@      @      �?     �E@      =@     `{@     Ps@      "@     �^@     @T@      (@      &@      @      >@     �q@       @     �z@      @      �?      D@      9@     �r@     �l@       @     @Z@      I@      &@      @      @      2@     @l@      @     @v@       @              7@      0@     `m@     �d@       @     �O@     �B@      @      @       @      *@     `a@      @     `f@      �?              *@       @      b@     �W@       @      D@      *@      @               @      @     �U@       @      f@      �?              $@       @     �V@     �Q@              7@      ?@      �?       @      �?      (@      K@       @     �R@      �?      �?      1@      "@     @P@     �P@      @      E@       @      �?      @              @      *@      �?      9@      �?      �?       @      @     �C@      0@      @      .@      7@              @      �?      @     �D@      �?     �H@                      "@      @      :@      I@      �?      ;@      (@      @      @      @      @     @W@       @     p@       @              @      @     @a@     �S@      �?      2@      $@       @      @      @      �?      Q@       @     `e@                      �?      @      S@      I@      �?      2@      @              @                      (@      �?      B@                                      .@      ,@              @      @       @              @      �?      L@      �?     �`@                      �?      @     �N@      B@      �?      &@       @       @       @               @      9@             �U@       @               @      �?      O@      <@                                       @               @      @              D@                              �?     �A@      @                       @       @                              6@              G@       @               @              ;@      6@                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ+��9hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�_�O[l�?�	           ��@       	                   �;@�$ߠ���?           ��@                            �? ��#��?I           ��@                           �?�x~v�?�           X�@������������������������       �\��U�?           ��@������������������������       ��Pi�6��?�           Џ@                           �?�A ���?�           0�@������������������������       ���c���?�            `t@������������������������       �>
ףp��?�             t@
                            �?�|�M��?�            �q@                           @���"&��?O            �\@������������������������       ���"�3c�?C            �W@������������������������       ��G�z�?             4@                           @��+�Y/�?n            �e@������������������������       �F��;5�?a            �b@������������������������       ��0�~�4�?             6@                           @��a��?�           <�@                           @�fH��E�??           �~@                          �7@����?!           �{@������������������������       ��i����?�            �s@������������������������       ��ܡ*���?R            �_@                           �?����|��?             F@������������������������       ���%����?            �@@������������������������       ��zv��?             &@                          �5@� �+Lm�?�           0�@                          �2@�qr�s�?�             s@������������������������       �$ou8���?Z            @a@������������������������       �Z��5;j�?h             e@                           @��
KF�?�            @s@������������������������       ��$_�V�?�            pp@������������������������       �\�D9�"�?            �F@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@     �B@     �C@      :@     �Y@     ؃@      :@     �@      4@       @      T@     �R@     P�@     �~@      :@     �o@     �c@      >@      =@      6@     �T@     �}@      5@     ��@      (@      @     �O@     �O@     P@     @v@      5@     �j@      b@      ;@      <@      2@      S@      {@      4@     (�@      &@      @      L@     �M@     �|@     �t@      .@     �h@      [@      .@      5@      *@      G@     �u@      0@     ��@      @       @     �@@      A@     �v@      k@       @     �^@     �H@      @      3@      $@     �@@     @g@      "@     �i@      @       @      2@      0@     `b@      V@      @     �N@     �M@      "@       @      @      *@     �c@      @     @t@       @              .@      2@      k@      `@       @     �N@     �B@      (@      @      @      >@     @V@      @     �\@      @      @      7@      9@      X@     �\@      @     �R@      &@      @      @      @      1@     �G@      @     �P@      @      �?      @      1@     �H@      H@      @     �C@      :@      @      @       @      *@      E@              H@      �?       @      1@       @     �G@     �P@      @     �A@      *@      @      �?      @      @     �E@      �?     @\@      �?              @      @      E@      :@      @      0@      @                              @      *@      �?     �K@                       @       @      2@      (@              @      @                              @      &@      �?     �C@                       @       @      1@      &@              @                                               @              0@                                      �?      �?                      $@      @      �?      @       @      >@              M@      �?              @       @      8@      ,@      @      (@      $@      @      �?      @       @      <@             �C@      �?              @       @      7@      ,@      @      (@                                               @              3@                                      �?                             �A@      @      $@      @      4@     �c@      @     �x@       @      @      1@      &@     �n@     �`@      @     �D@      (@              "@      @      @      K@       @     �g@       @              &@      @      _@      M@              3@      (@               @      �?      @     �G@       @     �f@       @               @      @     �\@      H@              0@       @               @      �?              B@       @      ^@                      @             �V@      B@              *@      @                              @      &@              N@       @              @      @      9@      (@              @                      �?      @              @               @                      @              "@      $@              @                      �?      @              @              @                      @              @       @               @                                               @              @                                      @       @              �?      7@      @      �?              1@      Z@      @     `j@      @      @      @       @     @^@     @S@      @      6@      &@      @                      (@      @@       @     �[@              @      @      @      M@     �D@              4@      @                              @      ,@              D@                      @      @     �B@      .@              "@      @      @                      @      2@       @     �Q@              @               @      5@      :@              &@      (@      @      �?              @      R@      �?      Y@      @                      �?     �O@      B@      @       @      (@      @      �?              @      L@      �?     �U@      @                      �?     �L@      :@      @       @                                              0@              *@                                      @      $@                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJC�gNhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�)����?�	           ��@       	                     �?�UŴ��?�           ��@                          �:@���]��?$           N�@                          �9@��%�`��?t           P�@������������������������       �WwN?B��?@           �@������������������������       � �Z���?4            �T@                           �?NX
�a��?�            0q@������������������������       �333333�?E             Y@������������������������       �0*��D�?k            �e@
                           @�im���?�           p�@                          �1@���2�?6           �~@������������������������       ����rm�?9            �U@������������������������       ���z�;��?�            @y@                          �2@�hB����?�            `h@������������������������       ��~_� �?'            �N@������������������������       �r/�����?\            �`@                           �?���;��?�           Б@                           @���{^�?@           0�@                           @*EDڅ�?�            `u@������������������������       �a�hg���?�            �n@������������������������       �ޟ���|�?5            �W@                           @��7V�?t             f@������������������������       ��H�y!�?Q            �_@������������������������       ��(\����?#             I@                          �2@O��B�d�?�           p�@                           @��.��q�?h            `c@������������������������       ���{8���?;            �T@������������������������       ��2�tk~�?-             R@                           �?������?%           0}@������������������������       �����C�?'            �J@������������������������       �p+9����?�            �y@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        g@      F@     �H@      @@     �X@     X�@     �A@     �@      5@      @     �Q@     �R@     ��@     �@      6@     @q@     �a@     �A@     �@@      9@      T@      {@      <@     ��@      .@      @      P@      O@     �@     �w@      4@     �k@      Y@      8@      6@      3@      I@     �u@      3@     @�@       @      �?     �E@     �B@     �y@     �p@      (@     �a@     �V@      0@      4@      1@     �D@     �s@      .@     �~@       @      �?      D@     �@@     �u@     �n@      (@     �^@     �V@      0@      4@      ,@      D@      r@      ,@     0~@      @      �?     �B@     �@@     �t@     `l@      (@      ^@      �?                      @      �?      8@      �?      &@       @              @              1@      2@               @      "@       @       @       @      "@      A@      @     �V@                      @      @     �P@      :@              2@      @      @       @      �?      @      ,@      @      =@                      @              (@      (@               @      @       @              �?      @      4@             �N@                              @      K@      ,@              $@     �E@      &@      &@      @      >@      V@      "@     @a@      @      @      5@      9@     �W@     @[@       @     @T@      =@      &@      @      @      3@      M@      @     @Z@      @      @      5@      0@      Q@     �Q@      @     �M@      "@      @              @      @      .@      �?      @                      @      @      0@      @      @      $@      4@       @      @      �?      ,@     �E@      @     �X@      @      @      1@      *@      J@     �O@      @     �H@      ,@              @       @      &@      >@       @     �@@              �?              "@      :@     �C@      �?      6@      @               @                      *@       @      @                              @      @      7@              @      &@              @       @      &@      1@              <@              �?              @      5@      0@      �?      1@      E@      "@      0@      @      2@      g@      @     �z@      @              @      *@     �k@     �_@       @     �K@      @@      @      $@       @      &@     �V@      @     �b@      @              @      @      W@     @R@              ?@      1@       @       @       @      @     �Q@      @     @U@      �?              @      @      R@     �E@              6@      .@       @       @       @      @     �D@      @      Q@      �?              @       @      H@     �A@              0@       @                              @      =@              1@                      @      @      8@       @              @      .@      @       @              @      5@       @     �P@       @                      �?      4@      >@              "@      .@       @       @               @      $@      �?      H@       @                      �?      ,@      7@              @              �?                      @      &@      �?      2@                                      @      @              @      $@      @      @      @      @     �W@       @     q@      @              �?      @     @`@      K@       @      8@       @              @       @       @      0@              M@                              �?     �I@       @              $@      �?                       @              @              >@                                     �A@      @              @      �?              @               @      $@              <@                              �?      0@      @              @       @      @      �?      @      @     �S@       @     �j@      @              �?      @     �S@      G@       @      ,@       @                                      $@      �?      4@                                      @      &@               @      @      @      �?      @      @      Q@      �?     `h@      @              �?      @      R@     �A@       @      (@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�6�_hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @��~����?�	           ��@       	                   �?@����?�            �@                          �2@�e�d��?�           t�@                            �?~�S�P��?�           h�@������������������������       �˶��02�?h           ��@������������������������       ���7N�?�            �i@                           �?R�����?�           ��@������������������������       �6�l��2�?           Љ@������������������������       ��V ���?�           ̑@
                           �?�橻�-�?&            �Q@                          �@@2G�����?             :@������������������������       �      �?	             0@������������������������       ���Q��?             $@                           @�ˠT��?             F@������������������������       ��>�>�?             >@������������������������       �T�r
^N�?             ,@                           �?dr)����?�           $�@                           @��,�%�?&           ~@                          �2@�+� �_�?�            �t@������������������������       ��0%t]�?5            �V@������������������������       �p���s�?�            @n@                           @�4Vk�Y�?`            �b@������������������������       �������?%            �J@������������������������       ���Ͱ��?;            �W@                          �2@h<a��?�           @�@                           @�5ǡG��?h            �b@������������������������       ���<���?Z            @`@������������������������       �Tg�x�P�?             5@                           @�O]�?$           }@������������������������       ���_q��?	            z@������������������������       �G��+'��?            �G@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@      >@      D@      >@     @Y@     p�@      ;@     4�@      5@      @     �T@     �P@     p�@     Ȁ@      .@     `m@     @g@      3@      ;@      ;@     @S@     �}@      5@     ��@      1@      @     �S@      M@     �@     �y@      ,@     @h@     @g@      3@      ;@      ;@     @S@     @}@      4@     ��@      .@      @     �S@     �L@     @      y@      ,@     @h@     �Q@       @      (@      @      7@     �`@      "@     �d@      @      �?      A@      6@     �[@      _@      "@     �K@     �J@              "@      @      0@     @Z@      @     �`@      @              ,@      ,@      V@      V@      @     �@@      1@       @      @       @      @      >@      @      >@              �?      4@       @      7@      B@      @      6@      ]@      1@      .@      6@      K@     �t@      &@     �~@      &@      @     �F@     �A@      x@     `q@      @     `a@      K@      "@      (@      @      A@      d@      @     �g@      @      �?      3@      2@     �a@     �[@      @      L@      O@       @      @      .@      4@     �e@       @      s@      @      @      :@      1@     �n@     �d@       @     �T@                                              &@      �?      A@       @                      �?      &@      $@                                                               @              3@                                      �?      @                                                              �?              .@                                                                                                              �?              @                                      �?      @                                                              "@      �?      .@       @                      �?      $@      @                                                              @      �?      @       @                               @      @                                                               @              "@                              �?       @                              =@      &@      *@      @      8@     �e@      @     �y@      @      �?      @      "@     @n@     @_@      �?     �D@      8@      @      $@              4@     �V@      @      b@      �?              @      @     �U@      P@      �?      6@      .@       @      $@              2@      Q@      @     �V@                      @       @     �N@      F@              0@      @              @               @      2@              <@                       @       @      7@      @              @      (@       @      @              0@      I@      @     �O@                      �?              C@     �D@              &@      "@      @                       @      7@      �?     �J@      �?              �?       @      :@      4@      �?      @       @      @                      �?      @              2@      �?                              (@      @      �?      @      @                              �?      2@      �?     �A@                      �?       @      ,@      ,@               @      @      @      @      @      @      U@       @     �p@      @      �?              @     `c@     �N@              3@                      �?       @      �?      &@             �L@                               @     �N@      &@              @                      �?       @      �?      "@              E@                               @      M@      $@              @                                               @              .@                                      @      �?                      @      @       @      �?      @     @R@       @      j@      @      �?              @     �W@      I@              ,@      @      @       @      �?      @      P@       @     �h@      �?      �?              @     �T@     �F@              $@      �?       @                              "@              (@       @                              (@      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��VhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @R�k��?�	           ��@       	                     �?��N@���?�            �@                          �0@it*ɑ�?5           Ġ@                           @(�gA~8�?J            �]@������������������������       ��Q#1�?            �G@������������������������       �)O���?,             R@                          �:@�����{�?�           ��@������������������������       ��9�je��?           d�@������������������������       �e�bLV$�?�             u@
                          �4@ �'~���?�           p�@                          �3@�nN7���?�            pt@������������������������       �z�(��?�            �o@������������������������       ���� :�?.            �R@                           @��w���?�            pv@������������������������       ��Io���?�            �s@������������������������       ��6�G���?             G@                          �=@��� ��?�           �@                           �?d' ND�?|           H�@                          �0@u�'����?%           �}@������������������������       �N贁N�?             .@������������������������       ��.��\a�?           �|@                           �?�����?W           ��@������������������������       ����ӡ��?�            Pu@������������������������       ��b�'�?{            �g@                           �?��Q��?2             T@������������������������       �      �?              @                           @B{	�%��?+             R@������������������������       �}�'}�'�?#             N@������������������������       ���8��8�?             (@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@     �A@     �H@      >@     �Y@     ��@      A@     ��@      2@      @     �S@      P@     Ї@     @}@      1@     �p@     �d@      7@     �B@      :@      U@     ��@      >@      �@      0@      @     �M@     �K@     0�@     �u@      0@     �j@     �]@      4@      :@      1@     �K@     �y@      :@     H�@      "@              C@     �@@     �y@     �l@      $@      c@      @               @      �?      @      5@      �?      1@       @                      @      <@      3@              (@      �?              �?                      @      �?      @                               @      3@      &@              @      @              �?      �?      @      1@              (@       @                      @      "@       @              "@      \@      4@      8@      0@      I@     �x@      9@     ��@      @              C@      <@     �w@     �j@      $@     �a@     @Y@      (@      6@      $@      E@     �t@      3@     p}@      @              :@      7@      s@      h@      $@      ^@      &@       @       @      @       @     �O@      @     @X@      �?              (@      @     �S@      4@              4@      H@      @      &@      "@      =@     @\@      @     �]@      @      @      5@      6@     �Z@     �]@      @     �O@      5@              @      @      .@     �N@      @      K@              �?      (@      .@     �A@      O@      @      B@      1@               @      @      *@     �H@      @     �G@              �?       @      "@      ?@     �D@       @      :@      @              �?               @      (@              @                      @      @      @      5@      @      $@      ;@      @       @      @      ,@      J@      �?     @P@      @      @      "@      @      R@     �L@              ;@      :@      @      @      @      ,@      D@      �?      I@      @      @       @      @     @Q@      H@              :@      �?              �?                      (@              .@      @              �?              @      "@              �?     �C@      (@      (@      @      3@     @d@      @     �w@       @       @      3@      "@     �n@     �]@      �?     �I@      B@      (@      (@      @      .@     �b@      @     �u@      �?       @      3@      @     �k@     �]@      �?     �I@      4@      $@       @              (@      T@      @     @`@      �?       @      2@      �?     @W@      O@              @@                                      �?      �?       @      �?                       @      �?      �?       @              @      4@      $@       @              &@     �S@      �?      `@      �?       @      0@              W@      N@              <@      0@       @      @      @      @     �Q@      �?      k@                      �?      @      `@      L@      �?      3@      &@      �?      @      @       @      D@      �?     @b@                      �?      @     @Q@      D@      �?      2@      @      �?      �?              �?      ?@             �Q@                               @     �M@      0@              �?      @                              @      &@              B@      �?                       @      7@                               @                              �?      �?              @                                                                      �?                              @      $@              @@      �?                       @      7@                              �?                              @      @              >@      �?                       @      0@                                                                      @               @                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�AeqhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �2@6��g��?�	           ��@       	                    @���0�?�           ��@                           �?����$�?�           p�@                           �?	iv^��?�            �r@������������������������       �dE�?[             b@������������������������       �k���?g            �c@                            @1�Y
�?+           �}@������������������������       �=�^�&_�?�            �w@������������������������       �9-�.]�??            @Y@
                            @�����?�            �q@                           @�)��?�?�            �n@������������������������       �9�5�3�?u            @h@������������������������       �:J�����?"             J@                           �?�������?             A@������������������������       �VUUUUU�?             .@������������������������       �d�����?             3@                           �?h�G4~-�?           F�@                            �?�O����?�           ��@                           �?�T�f�?�           �@������������������������       �'6�i���?�             k@������������������������       �p�ݯ�?           �|@                          �9@+ʔ���?G           (�@������������������������       �����	�?�            y@������������������������       �?��C��?O             ]@                            @<�Z�?           ��@                           @�Ųe��?�           H�@������������������������       ��4��!�?           ��@������������������������       �֔]�?�            `w@                           �?���bDg�?'           �~@������������������������       ��N��'�?/            �R@������������������������       �ƵHPS�?�             z@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `i@      ?@      C@      6@     �Z@     ��@     �A@     ��@      @      @     �R@      L@     ��@     ��@      1@     `q@     �R@      @      1@      @     �@@      f@       @     �l@              �?      :@      9@     `i@     �e@       @      S@     �I@      @      *@      @      7@     �a@      @     `c@                      2@      3@     �d@      _@      @     �J@      2@              "@      �?      *@     �G@      @     �T@                      @      @     �F@      K@       @      5@      &@              @              (@      *@       @      D@                      @      @      9@      5@       @       @      @              @      �?      �?      A@      �?      E@                                      4@     �@@              *@     �@@      @      @      @      $@     @W@      @     @R@                      ,@      .@     �]@     �Q@      @      @@      ;@      @      @      @      @     @S@      @     �N@                      (@      *@      R@     �N@      @      ?@      @      @                      @      0@              (@                       @       @     �G@      "@              �?      7@              @              $@      B@       @     �R@              �?       @      @     �C@      I@      @      7@      6@              @              $@      ?@      �?      N@              �?       @      @      <@     �H@      @      7@      2@              @               @      =@      �?     �H@                      @      @      :@      ?@      @      2@      @              �?               @       @              &@              �?      @      @       @      2@              @      �?                                      @      �?      .@                                      &@      �?                      �?                                      �?              @                                      @      �?                                                              @      �?      "@                                      @                              `@      8@      5@      2@     @R@     p~@      ;@     ��@      @      @      H@      ?@     ��@     0v@      "@     @i@      Q@      *@      1@      &@      H@     �j@      "@     pr@      @       @      5@      0@     �i@     �a@      @     @^@      E@      @      "@      @      ;@     `a@      @     �c@       @              *@      "@      \@     �P@       @      S@      "@      @      @      @      *@      B@             �E@                      $@      �?     �A@      5@             �A@     �@@      @       @      @      ,@     �Y@      @     @\@       @              @       @     @S@      G@       @     �D@      :@      @       @      @      5@     �R@      @     `a@      �?       @       @      @     �W@      S@       @     �F@      1@      @      @      @      5@      J@      @     �X@      �?       @       @      @     @T@      N@       @     �B@      "@      @      @                      6@      �?      D@                              �?      *@      0@               @     �N@      &@      @      @      9@      q@      2@     ��@      @      �?      ;@      .@     0v@     �j@      @     @T@      I@      @       @      @      6@     �g@      *@     �u@       @      �?      6@      *@     `p@     �c@      @     @R@     �D@      @       @       @      2@     `a@      $@     �k@       @              .@      @     �f@     �Y@      @      H@      "@      @              @      @      I@      @     �_@              �?      @      @      T@      L@              9@      &@      @       @       @      @     @U@      @     �j@       @              @       @     @W@     �J@      �?       @      @                                      $@      @      =@                                      "@      2@              �?      @      @       @       @      @     �R@      �?      g@       @              @       @      U@     �A@      �?      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��ehG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @zb�Z4��?�	           ��@       	                    @    ���?�            �@                            �?I��"�%�?           �@                          �=@x�_�?�           Ј@������������������������       �sI��P4�?�           h�@������������������������       ��h�!�?            �F@                          �1@�@�Ԫ�?&           |�@������������������������       �<�'܀w�?�            �n@������������������������       �B$yCɒ�?�           X�@
                          �:@@���=�?�           8�@                           @$�g���?�           ��@������������������������       ��h\�x�?           Pz@������������������������       ���"Ac��?�             k@                           @h���%�?O             a@������������������������       �H�7�&��?             .@������������������������       ��D���?G            �^@                           �?᜗  k�?�           $�@                           @����Gq�?�            �t@                           �?5�Qa&�?�            pr@������������������������       �1w�5�?y             g@������������������������       ��g���?@            �[@������������������������       ��������?            �A@                           �?U��0�4�?�           ��@                          �=@r.!ƎQ�?�            `s@������������������������       ��q�m'�?�             r@������������������������       �      �?             4@                           �?8�n��?*           �|@������������������������       ���.�t�?7            �U@������������������������       ���\9��?�             w@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �l@      7@      B@      6@     �Z@     `�@      ;@     �@      4@      @     �U@     �Q@     ��@     �@      *@     Pp@     �e@      5@      7@      1@      V@     �~@      5@     ؆@      .@      @     �R@     �M@     �~@     �w@      (@     `k@     �`@      &@      4@      &@     @R@     �v@      .@     �~@      *@      @      M@      F@     �v@     �o@      $@     �e@     �C@      @      @      @      1@     �b@      @     �n@      @              0@      1@     @b@     �W@      @      G@     �C@      @      @      @      .@     @b@      @     �k@      @              0@      1@     �`@     @W@      @     �F@                                       @      @              8@                                      (@      �?              �?     �W@      @      1@       @      L@     `j@      &@      o@      $@      @      E@      ;@     `k@     �c@      @     �_@      4@       @      @      �?      "@     �L@      �?      :@       @      �?      @      @      D@     �D@      �?      9@     �R@      @      &@      @     �G@     @c@      $@     �k@       @      @     �A@      6@     `f@     �]@      @     �Y@     �C@      $@      @      @      .@     �_@      @     �m@       @      �?      0@      .@     �_@     @_@       @      G@     �B@      $@      @      @      .@     �[@      @     �d@       @      �?      *@      &@     �Z@     �\@       @      B@      8@       @       @      @      @      T@       @     �Y@       @               @      @     @U@     �R@      �?      2@      *@       @      �?              &@      ?@       @     @P@              �?      @      @      5@      D@      �?      2@       @                                      .@       @     �Q@                      @      @      4@      &@              $@                                                              (@                      �?       @                                       @                                      .@       @      M@                       @       @      4@      &@              $@     �L@       @      *@      @      3@     �h@      @     �v@      @              *@      &@     `m@     @`@      �?      E@      1@               @              @     �I@      @     �W@                      @       @     �W@      >@              8@      *@               @               @      E@      @     �T@                      @      �?      W@      =@              5@       @               @               @      =@      �?      N@                       @      �?      G@      6@              (@      @                                      *@      @      7@                      @              G@      @              "@      @                               @      "@              &@                      �?      �?      @      �?              @      D@       @      &@      @      .@      b@       @     �p@      @              @      "@     �a@      Y@      �?      2@      2@              "@       @      $@     �L@       @     @V@      @              @       @     �E@      M@              &@      (@              "@       @      "@      L@       @     �T@       @              @       @     �D@      M@              &@      @                              �?      �?              @      @                               @                              6@       @       @      @      @      V@             `f@                       @      @     @X@      E@      �?      @      $@               @              @       @              B@                                      ,@      $@              @      (@       @              @      �?      T@             �a@                       @      @     �T@      @@      �?      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�ghG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?.����?�	           ��@       	                     @z��/�?F           H�@                          �?@�Pp4i�?"           �@                           @�QV��w�?           p�@������������������������       ���u��t�?�           �@������������������������       �g	J�R��?;            �U@                            �?�H���?             ?@������������������������       �      �?
             0@������������������������       ��X�%��?
             .@
                           @t>��!_�?$           p}@                           @�@=��?�            0w@������������������������       �hy��?�            @m@������������������������       �\��)�?W             a@                           @��#����?=             Y@������������������������       �� {�/��?*             Q@������������������������       �     �?             @@                            @�[�R
�?T           �@                            �?VЈDd��?�           ��@                          �0@�]�����?�           8�@������������������������       ��ߋm��?*            �P@������������������������       ���D����?�           0�@                           �?��a���?�             w@������������������������       ��Y�R_�?.            �Q@������������������������       �rvT����?�            �r@                           @�_��<�?{           ȁ@                          �2@8�b����?&           �{@������������������������       ��D �D �?M            �]@������������������������       �xt�>v��?�            `t@                          �4@M�*`W��?U             _@������������������������       ���x�(��?!             G@������������������������       �^�"R��?4            �S@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        j@      ?@      E@      7@     �[@     H�@      ;@     ̐@      8@      $@     �T@      P@     x�@     �@      5@      p@     @Z@      4@      <@       @      P@     �t@      $@     �y@      0@      @     �E@      A@     Ps@     @l@      @     �`@     �P@      .@      7@       @      I@     @o@      $@     0q@      (@      @     �C@      >@     @k@     �c@      @      [@      P@      .@      7@       @      I@     �n@      $@     0p@      (@      @     �C@      >@      k@     @c@      @      [@      O@      .@      3@       @     �F@     @m@      $@     �m@      $@      @     �C@      =@     �i@      a@      @      X@       @              @              @      $@              6@       @                      �?      (@      1@              (@      @                                      @              0@                                      �?      @                                                               @              (@                                               @                      @                                      @              @                                      �?      @                      C@      @      @              ,@     �S@             �`@      @      �?      @      @     �V@     �P@       @      8@      >@      @      @              (@     �P@             �V@       @              @       @     �S@      K@       @      5@      9@      �?      @              @     �A@             �K@       @              @              J@     �B@              0@      @      @                       @      @@              B@                               @      :@      1@       @      @       @              �?               @      (@              E@       @      �?      �?       @      *@      *@              @       @              �?                      &@              <@       @      �?               @      @      "@              @                                       @      �?              ,@                      �?              $@      @                     �Y@      &@      ,@      .@      G@      v@      1@     ؄@       @      @     �C@      >@     �{@     �q@      ,@     �_@     �T@       @      $@      &@      D@     @p@      *@     �{@      @      �?      A@      ;@     �s@     �l@      ,@     �Z@     �K@      @      @      &@      7@     @j@      $@     �w@      @              0@      0@     `o@     �d@      @     �R@      @                                      0@               @                       @       @      &@      "@              *@      I@      @      @      &@      7@     @h@      $@     0w@      @              ,@      ,@      n@     �c@      @     �N@      ;@       @      @              1@      I@      @      P@       @      �?      2@      &@     �O@      O@      "@     �@@       @               @              @      .@              $@       @      �?      �?              0@      @       @      @      9@       @      @              ,@     �A@      @      K@                      1@      &@     �G@     �L@      �?      ;@      5@      @      @      @      @      W@      @      l@      @       @      @      @      `@     �I@              3@      2@      �?      @      @      @     �N@      @     �g@      @       @       @      @     �W@     �B@              1@      @                      @       @      @             �E@                              �?     �E@      &@              @      (@      �?      @      �?      @      K@      @     @b@      @       @       @       @      J@      :@              ,@      @       @                      �?      ?@             �A@                      @             �@@      ,@               @       @      �?                      �?      @              0@                      @              (@      @              �?      �?      �?                              ;@              3@                                      5@       @              �?�t�bub�     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�`�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx         
                    �?�GWK��?�	           ��@       	                    @�n�*� �?f           ��@                           @X!t��?]           X�@                          �=@��&8,>�?]           �@������������������������       ��8m.�C�?:           �@������������������������       �d}h���?#             L@                           @�派o�?            �y@������������������������       �0�n�"��?�             o@������������������������       �*�hi&�?j            �d@������������������������       �0�����?	             2@                           @�(��n�?K            @                          �7@8�0��?�           Ԙ@                          �0@�|{z��?�           ��@������������������������       ���Z���?4            �T@������������������������       �c�H���?�           X�@                          �?@!�Z�0��?'           �|@������������������������       �Rm/6��?           Pz@������������������������       �\���(\�?             D@                           @D��dS�?X           `�@                           @�=��?           �z@������������������������       ��4�-���?�            @v@������������������������       �������?-             R@                           @     ��?K             `@������������������������       �)\���h�?1             T@������������������������       ��8��8��?             H@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      C@     �A@      8@     �Z@     ��@      ?@     `�@      4@      @      V@     �J@     ��@     �}@      4@     0r@     @]@      3@      <@      .@      O@     �s@      3@     �{@      ,@      @      C@      @@     �r@     @l@      @      `@     @\@      3@      <@      .@      O@     �s@      0@     �{@      ,@      @      C@      @@     �r@      l@      @     �^@     �V@      .@      7@      ,@      L@     �m@      $@     0t@      "@      @      B@      2@     �l@      d@      @      Z@     @T@      .@      7@      ,@     �H@     �m@      $@     �r@       @      @      B@      0@      l@     �c@      @      Z@      $@                              @      @              9@      �?                       @      @       @                      6@      @      @      �?      @     �S@      @     �]@      @      �?       @      ,@     �P@     �O@       @      3@      4@      @      @      �?      @      J@      @     �L@      @                       @     �E@      A@      �?      $@       @      �?                      �?      :@      �?     �N@      �?      �?       @      @      8@      =@      �?      "@      @                                       @      @      �?                                      �?       @              @     @Z@      3@      @      "@     �F@      v@      (@     ��@      @       @      I@      5@     pz@     �n@      .@     `d@     @V@      &@      @       @      @@     �n@      $@     0�@      @      �?     �@@      3@     `t@      c@      $@     �^@      R@      @      @      @      (@      h@       @      w@      �?      �?      :@      *@     �i@     �]@      @     �U@      @                                      :@              2@                      @      @      ,@      @              @     �P@      @      @      @      (@     �d@       @      v@      �?      �?      7@      $@      h@     @\@      @     �S@      1@       @      �?      �?      4@      K@       @     �b@      @              @      @     �]@     �A@      @     �B@      0@       @      �?      �?      3@      J@       @     �_@      �?              @      @     �[@     �A@       @     �@@      �?                              �?       @              5@       @                               @              �?      @      0@       @      �?      �?      *@     �Z@       @      c@       @      �?      1@       @     @X@     @W@      @      D@      0@      @      �?      �?       @     �T@       @     �_@       @      �?      0@             @S@     @Q@      @      0@      @      @      �?      �?      @     �R@             �Z@       @      �?      &@             �P@     �N@      @      &@      "@                              @       @       @      5@                      @              &@       @              @              @                      @      8@              9@                      �?       @      4@      8@              8@              @                      @      5@               @                      �?       @      *@      2@              "@                                              @              1@                                      @      @              .@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�+.hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @�.FH�a�?�	           ��@       	                     @�SZR�e�?f           �@                           �?W����?*           $�@                          �>@�U.�J��?�           x�@������������������������       �<|M����?�           ��@������������������������       �     ��?	             0@                          �<@� %�?�           Є@������������������������       �9�,H��?�           ��@������������������������       ��Ł�r��?             C@
                           �?4�@}K��?<           @                           �?���·g�?�            @o@������������������������       �����P�?w            @h@������������������������       ��m۶m��?#             L@                           @@�+����?�            �n@������������������������       ���;���?�            @l@������������������������       ���kv�?             5@                          �0@��m�
M�?P           ��@                           @�V�½��?C            �X@                            �?��+j��?.            �P@������������������������       ��G�z�?             D@������������������������       �θ	j�?             :@                           �?~fL���?            �@@������������������������       ��d�����?             3@������������������������       ��m۶m��?             ,@                           �?�@��5�?           ��@                          �1@8p����?           ��@������������������������       ���Q�d��?B            �\@������������������������       ����;Q��?�           ��@                           !@
LQZǤ�?�           �@������������������������       �M]aw��?�           ��@������������������������       �paRC4%�?             1@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      >@     �A@      =@      Z@     �@      >@     d�@      5@      $@     �S@      M@     ��@     @      *@      m@     �W@      ,@      :@      0@      M@      s@      @     �@      &@      @      ?@      ?@     �w@     �e@      @     @^@      U@      &@      1@      ,@      I@     `l@      @     pt@      @       @      ;@      <@     �p@      `@      @      V@      B@      @      &@      $@      B@     �[@       @      a@      @       @      2@      ,@     �[@     �P@      @      L@     �A@      @      &@      $@      B@     @[@       @     �_@      @       @      2@      ,@     �[@     �P@      @     �J@      �?                                       @              $@                                                              @      H@      @      @      @      ,@      ]@      @     �g@       @              "@      ,@     �c@     �O@       @      @@      F@      @      @      @      ,@      Z@      @     �g@                      "@      "@      c@     �N@      �?      <@      @      �?                              (@               @       @                      @      @       @      �?      @      $@      @      "@       @       @     �S@             @g@      @       @      @      @     @[@     �F@             �@@      @      @      @              @      G@              U@      @               @      �?     �I@      ;@              0@      @      @       @              @      D@             �O@                       @      �?     �D@      2@              .@                      @                      @              5@      @                              $@      "@              �?      @               @       @      @     �@@             �Y@               @       @       @      M@      2@              1@      @               @       @             �@@             �V@                       @       @     �K@      2@              1@                                      @                      &@               @                      @                             �W@      0@      "@      *@      G@     y@      8@     ��@      $@      @     �G@      ;@     px@     0t@       @      \@      @               @      �?       @      3@      �?      &@                       @       @      2@      :@              &@      @               @      �?      �?      ,@               @                      �?       @      *@      *@               @       @               @                       @               @                              �?      &@      @              @      �?                      �?      �?      @              @                      �?      �?       @      @              �?      �?                              �?      @      �?      @                      �?              @      *@              @      �?                              �?       @      �?      @                                      @      @                                                              @                                      �?              �?      @              @     �V@      0@      @      (@      F@     �w@      7@     h�@      $@      @     �F@      9@     Pw@     �r@       @     @Y@     �K@      &@      @      @      ;@     @b@      $@     �i@       @      @      1@      *@     �b@     �]@      @      H@      @      @       @              @      4@       @     �A@              @      @       @      *@      "@              @     �H@       @       @      @      5@     �_@       @      e@       @      �?      *@      @      a@     @[@      @      F@     �A@      @      @      "@      1@     �m@      *@     x@       @       @      <@      (@     �k@     `f@      @     �J@     �A@      @      @      "@      1@     �l@      *@     �w@       @       @      <@      (@     �k@      f@      @     �I@                                               @              @                                      �?       @               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��`hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �<@���Rj�?�	           ��@       	                   �0@�zaM��?�           (�@                           @�(E��?�            �j@                           �??(� ���?_            `c@������������������������       ��.��6i�?1            �S@������������������������       �vq`����?.             S@                           @;�^
�$�?"            �M@������������������������       ��ۘ9��?            �G@������������������������       �UUUUUU�?             (@
                           @3�o�f�?f           |�@                          �1@B��yK�?�           p�@������������������������       ��ܩ���?�             g@������������������������       �8���.�?3           ��@                            @K	�5]�?�           ��@������������������������       �w=}e��?V           ��@������������������������       ��A���?\           ��@                           @B�a����?�            Ps@                            @+��9���?�            �i@                          �=@v�9w�q�?M            �^@������������������������       ��h�*$��?             C@������������������������       ��=d���?2            @U@                           �?6�]��?3            @T@������������������������       �ffffff�?             D@������������������������       �>YV����?            �D@                           @ܥ�Xk��?=            @Z@                            �?	�J0��?,            �R@������������������������       �I��&���?             =@������������������������       �$G�h��?             G@������������������������       �<+	���?             >@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      @@     �A@      4@     �[@     ��@      ;@     @�@      0@       @     @R@     �R@     X�@     �|@      2@     `q@     `i@      =@     �A@      4@     �Z@     ��@      8@     �@      $@       @      P@     @Q@     �@     �{@      1@     `p@      &@      �?      @      @      &@      D@       @     �@@      �?              @      *@      <@     �C@      �?      9@      @      �?      �?      @      "@      =@       @      9@      �?              @      (@      6@      4@              6@      �?      �?      �?      @       @      0@      �?       @      �?                      @      ,@      0@              @      @                              �?      *@      �?      1@                      @      @       @      @              3@      @               @               @      &@               @                              �?      @      3@      �?      @      @               @                      &@               @                              �?      @      1@      �?              @                               @                                                               @       @              @      h@      <@      @@      1@     �W@     ��@      6@     (�@      "@       @     �N@      L@     8�@     py@      0@     �m@     �W@       @      8@      "@     �I@     �m@      "@     �y@       @      �?      7@      9@     pt@     �_@      @     @T@      3@              @              @      D@             �D@                              @      C@      4@      @      &@      S@       @      1@      "@      H@     �h@      "@      w@       @      �?      7@      6@     r@     �Z@      @     �Q@     @X@      4@       @       @      F@     pt@      *@     `�@      @      @      C@      ?@      t@     �q@      $@     �c@     @R@      &@      @      @     �A@     �k@      &@     �w@      @      @     �@@      :@     @k@     @j@      $@      a@      8@      "@      �?       @      "@     @Z@       @     @j@       @       @      @      @     �Y@     �Q@              4@      3@      @                      @     �I@      @     @a@      @              "@      @      D@      ,@      �?      0@      1@      @                      @     �C@      @     @T@      @              @      @      6@      @      �?      ,@      $@      @                       @      =@      @      B@      @              @      @      &@       @              *@      @      @                              @              &@                      @      �?      @      �?              @      @                               @      8@      @      9@      @              �?      @       @      �?              $@      @                               @      $@             �F@       @                              &@       @      �?      �?      @                              �?      @              0@       @                              @       @      �?                                              �?      @              =@                                      @                      �?       @                                      (@             �L@      �?               @      �?      2@      $@               @      �?                                       @              G@                       @      �?      @      "@               @                                                              3@                              �?      @      @                      �?                                       @              ;@                       @              @      @               @      �?                                      @              &@      �?                              (@      �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�XOhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?Ya�����?�	           ��@       	                   �;@�("]�0�?A           ��@                            @�N��F(�?�           p�@                            �?^t/�+��?�           8�@������������������������       ����:�?           h�@������������������������       ��u���2�?�            r@                           @� ����?           �|@������������������������       �rĜ��m�?           `{@������������������������       ���8��8�?             8@
                          �?@��P�4��?\            �a@                            �?���*�{�?H             [@������������������������       �Q?��2��?%             M@������������������������       ���MbX�?#             I@                           @�RMw�?            �A@������������������������       �9��8���?             8@������������������������       �b���i��?             &@                           @�����?E           ��@                           @ �Ub��?#           �@                          �0@�1r����?.           <�@������������������������       �����k�?             C@������������������������       ��������?           ��@                          �=@[�.H���?�            `w@������������������������       �X/ �>��?�            �u@������������������������       �J��LQ�?             7@                            �?�<Tp��?"           �}@                          �7@_c�>��?<            �X@������������������������       �K�m_8��?3            �T@������������������������       ��r����?	             .@                           @��#.y�?�            pw@������������������������       ��A8K%q�?`            �f@������������������������       ���}��?�            `h@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@      @@      ?@      9@      Y@     h�@      8@     �@      7@      (@      S@     �U@     8�@      ~@      3@     pr@     @X@      7@      7@      (@      N@      s@      $@      {@      *@      @      B@      E@     �r@     �m@      (@     �c@      V@      1@      3@      (@     �J@     @r@      $@     @x@      &@      @      ?@      E@     �q@      l@       @     �a@      P@      ,@      1@      (@      D@     �i@      @     �m@      &@      @      9@      B@     �g@     �d@       @     �^@     �H@      @      $@      $@      9@      f@      @     `i@      @      �?      3@      3@      c@     �Y@      @      V@      .@      "@      @       @      .@      ?@       @     �A@      @      @      @      1@      C@      P@      @     �A@      8@      @       @              *@     @U@      @     �b@              �?      @      @      W@      M@              3@      8@      @       @              &@      S@      @     �b@              �?      @      @     �V@      I@              2@                                       @      "@               @                                       @       @              �?      "@      @      @              @      (@              G@       @              @              4@      (@      @      0@       @      @      @              @      @              =@                      @              1@      @      @      .@      @      @      @               @      @              $@                      @              "@      �?              *@      @                              @      @              3@                                       @      @      @       @      �?                                      @              1@       @                              @      @              �?                                               @              ,@       @                              @       @              �?      �?                                      @              @                                              @                     �W@      "@       @      *@      D@     �u@      ,@     ��@      $@      @      D@      F@     �}@     `n@      @      a@     �T@      @      @      $@      ;@     0q@      $@     P@      @      @      9@      =@     �w@     `j@      @     @X@     �K@      @      @       @      9@     �h@       @     �x@      @      @      5@      ;@     @s@     �b@      @     �S@       @                                      @              @                              �?      .@       @              @     �J@      @      @       @      9@     @h@       @     px@      @      @      5@      :@     Pr@     �a@      @     �R@      <@      �?               @       @     @S@       @     �Z@       @              @       @      Q@     �N@      �?      2@      <@      �?               @       @     �R@       @     @Y@                       @       @     �M@     �N@      �?      .@                                               @              @       @               @              "@                      @      (@      @      @      @      *@     �R@      @     `c@      @              .@      .@      X@      @@       @      D@              @               @              (@             �I@      �?               @              (@      "@       @      @              @               @              (@              C@      �?               @              $@      "@       @      @                                                              *@                                       @                              (@       @      @      �?      *@      O@      @      Z@      @              *@      .@      U@      7@              B@      @              @      �?      @      8@      �?      H@       @              @      @     �L@      @              3@       @       @                      @      C@      @      L@      �?              $@       @      ;@      2@              1@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�N0JhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @.΋�w�?�	           ��@       	                    �?"�=1l��?�           .�@                           @���^��?"           �@                           @���e��?R           �@������������������������       �r-�T��?�            �@������������������������       �����?U             `@                          �8@��a��?�             t@������������������������       �c>��J�?�            �n@������������������������       �L ���u�?0            @S@
                          �0@��	fV�?�           P�@                            �?JR��?9            �U@������������������������       ��E��Y��?+             O@������������������������       ��z6�>�?             9@                            �?1�k;�?�           ��@������������������������       �L,<H]�?�           �@������������������������       �H��5��?�            �w@                           �?����?�           Ȑ@                           @�ȫRK�?1           �|@                           @����g�?�            `r@������������������������       ��!����?�            �o@������������������������       ��������?             D@                          �1@t*�$ �?e            �d@������������������������       �N�zv�?             6@������������������������       ���l���?W            �a@                          �2@ ;͐P�?�           8�@                           @�����?m             e@������������������������       �����K�?K             ]@������������������������       ��E��
��?"             J@                           @���Vo��?           �{@������������������������       �~+��4�?�            �x@������������������������       ������j�?             H@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      :@      E@      =@      [@     ��@      C@     ��@      4@      @     �P@     �L@     p�@     x�@      0@     @l@      e@      7@      ?@      9@     �W@     �}@      ?@     h�@      .@      @     �K@      H@     p@     �{@      *@     �g@      V@      &@      8@      1@      J@     @l@      4@     �p@      $@      @      6@      ;@     `j@     �h@      @      X@      Q@      "@      3@      1@     �F@     `f@      "@     �h@       @      @      5@      6@     `c@      `@      @      S@      P@      @      3@      .@     �D@     �b@       @     `f@      @      @      &@      ,@     �a@     �[@      @      O@      @       @               @      @      >@      �?      2@       @              $@       @      .@      3@              ,@      4@       @      @              @     �G@      &@      R@       @       @      �?      @      L@     @Q@      @      4@      4@       @      @              @      E@       @      I@       @       @      �?      @     �F@     �E@      @      &@                                      �?      @      @      6@                                      &@      :@              "@     @T@      (@      @       @      E@     `o@      &@      |@      @             �@@      5@     @r@     �n@      @     @W@      @                                      7@              &@                      @      @      .@      0@              @      @                                      ,@              &@                      @      �?      *@      "@              @                                              "@                                              @       @      @              �?      S@      (@      @       @      E@     �l@      &@     P{@      @              >@      ,@     Pq@     �l@      @     �U@     �E@      $@      @      @      5@     �e@      "@     �w@      @              *@      "@      k@      c@      @     �H@     �@@       @       @       @      5@      L@       @     �N@      �?              1@      @      N@     �S@       @     �B@     �I@      @      &@      @      ,@     �f@      @     py@      @       @      &@      "@     �j@     �\@      @     �B@     �@@      @      "@       @      @     �V@      @     @`@      @      �?      "@      @     @V@      J@      �?      4@      1@      �?      @       @      @      P@      @     @P@       @              @       @     �Q@     �@@              .@      *@      �?      @              @      L@      @      N@       @               @       @      Q@      9@              $@      @               @       @               @              @                      @              @       @              @      0@       @       @                      ;@       @     @P@      �?      �?      @       @      2@      3@      �?      @       @                                      @       @      @                      @      �?       @       @              @      ,@       @       @                      8@              O@      �?      �?              �?      0@      1@      �?       @      2@               @       @      @     @V@       @     Pq@       @      �?       @      @     �_@     �O@       @      1@       @              �?      �?      @      2@              O@                                     �J@      1@              @      @                      �?              *@             �B@                                      F@      (@              @      @              �?              @      @              9@                                      "@      @              �?      $@              �?      �?      @     �Q@       @     �j@       @      �?       @      @     @R@      G@       @      (@      @              �?      �?      @     �K@       @     �h@      �?      �?       @      @     @Q@      F@       @      $@      @                                      0@              2@      �?                       @      @       @               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��KhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?3	��z�?�	           ��@       	                    �?hd񑂯�?           (�@                           �?ro�����?:           �}@                          �6@�%Nn[#�?v            @f@������������������������       �CMu���?R            �^@������������������������       ��m۶m��?$             L@                           �?�B����?�            �r@������������������������       ��� �U�?_            �a@������������������������       ��gb�8�?e            �c@
                            �?`*�m���?�           X�@                          �:@�z�����?s            �i@������������������������       ��Cb��?k            �g@������������������������       �     ��?             0@                           �?��q��?c           ��@������������������������       � �{��t�?�            �t@������������������������       �#�XoC�?�            �j@                          �<@D�	��R�?�           ��@                            @S6-���?�           &�@                            �?`��K���?J           p�@������������������������       �Cy[K�?�           �@������������������������       ����$eE�?�           |�@                           @���<���?�           ��@������������������������       �; ~|��?�           0�@������������������������       ��������?             1@                           @��޵o9�?�            �m@                          �A@���:Z��?x            �g@������������������������       ��i�r�?q            �f@������������������������       ��<ݚ�?             "@                            �?^��y�p�?            �F@������������������������       ��z6�>�?             9@������������������������       ��G�z��?             4@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@     �B@      F@      5@     �[@      �@      @@     P�@      3@      @     �Q@     �H@     ��@     p~@      ;@      q@     �R@      @      0@       @      =@     �h@      @     �r@      @      �?      4@      3@     pq@     �c@      @     �X@      4@      @       @      @      @     �R@      @     �`@      �?              0@      $@      W@     �L@       @     �I@      @              �?              @      7@              F@      �?               @      @     �D@      7@             �@@      @              �?              �?      2@              =@      �?               @       @      8@      &@              >@                                       @      @              .@                               @      1@      (@              @      1@      @      @      @      �?      J@      @     �V@                      ,@      @     �I@      A@       @      2@      @              @      �?             �A@      @      D@                      @      �?      3@      (@      �?      "@      $@      @               @      �?      1@              I@                      @      @      @@      6@      �?      "@     �K@      @       @      @      9@     �^@      @     �d@      @      �?      @      "@     `g@     �Y@      @     �G@      ,@               @      @      @     �H@      �?     �D@                              �?      K@      >@      �?      @      ,@               @      @      @      H@      �?     �B@                              �?     �E@      >@      �?      @                                              �?              @                                      &@                             �D@      @      @      �?      5@     �R@       @     @_@      @      �?      @       @     �`@      R@      @     �E@      ?@      @      @      �?      0@     �G@       @      O@      @      �?      @      @     �Q@      G@      @      =@      $@              �?              @      ;@             �O@      �?              �?      @      O@      :@              ,@     �]@      ?@      <@      *@     @T@     �}@      :@     @�@      ,@      @      I@      >@     �~@     �t@      4@     �e@     �[@      <@      9@      *@     @S@     �{@      8@     Ѕ@      $@      @     �G@      =@     �{@     �s@      3@      d@     �V@      0@      3@      $@      M@     �t@      3@     p{@      @      @     �E@      5@     `s@     �m@      1@      a@      6@      &@      &@      @       @      `@      @      g@      @              (@      @      `@     @S@      @      :@      Q@      @       @      @      I@     @i@      ,@     �o@      @      @      ?@      0@     �f@      d@      $@     �[@      5@      (@      @      @      3@     �[@      @     0p@      @      �?      @       @      a@      T@       @      9@      5@      (@      @      @      3@     �Y@      @      p@      @      �?      @       @     �`@     @S@       @      8@                                              @              �?                                      @      @              �?      @      @      @              @     �@@       @     �[@      @              @      �?     �D@      &@      �?      *@      @      @      @              @      8@       @     �W@      @              @      �?      8@       @      �?      *@      @      @      @              @      4@       @     @W@      @              @      �?      7@      @      �?      *@                                              @               @                                      �?       @                                                      �?      "@              .@                                      1@      @                                                              @               @                                      @      @                                                      �?       @              @                                      $@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJt�xhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@���Q^��?�	           ��@       	                   �8@�Yh޺�?�           P�@                           �?]�����?f           z�@                           @����w]�?V           D�@������������������������       ���J�R�?�           0�@������������������������       ����MK�?�            Pt@                            @�1�?t%�?           ��@������������������������       ����]%��?           Ԓ@������������������������       �x���o�?           p{@
                            @��,u;�?+           �~@                            �?�0v���?�            u@������������������������       �V9q@���?�             p@������������������������       ��IW�U7�?.            �S@                           �?�Lw-+�?a            @c@������������������������       ����o^M�?&             N@������������������������       ��ͯ3��?;            �W@                            @��:���?           z@                           �?��5����?�            pr@                           �?	�DG��?E            �Z@������������������������       �u#�����?             C@������������������������       �t�F��?,             Q@                          �=@�/�%�?x            �g@������������������������       �������?1             R@������������������������       �������?G            @]@                           @�N�����?T            �^@                           �?�u���?G            �Y@������������������������       ���ˠ�?             &@������������������������       ���Y[}Q�?@            �V@������������������������       ��������?             4@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@     �A@     �I@      =@     �X@     0�@     �E@     X�@      1@      "@     �O@     @R@     Ȇ@     �@      6@     pp@      i@      =@      H@      =@      V@     ��@      D@     ��@      ,@       @      L@      P@     ��@      ~@      1@     �n@     �f@      9@      G@      2@      T@      @      B@     ȉ@      (@       @     �K@      M@     �@     �x@      1@      j@     @V@      ,@     �B@      @     �G@      m@      .@      s@       @      @      3@      ;@     @n@      h@      *@     �Z@     @P@      "@      <@      @      G@     �d@       @     �m@      @      @      1@      .@     �g@     @b@      @     �V@      8@      @      "@              �?      Q@      @     �Q@       @      @       @      (@     �I@     �G@      "@      .@      W@      &@      "@      *@     �@@     pp@      5@     8�@      @      �?      B@      ?@      s@      i@      @     �Y@      S@      &@      @      "@      =@     �h@      2@     �t@      @      �?      A@      :@     @j@     �c@      @     �W@      0@              @      @      @     @P@      @     �g@      �?               @      @     �W@     �F@              @      3@      @       @      &@       @     @Q@      @     @_@       @              �?      @     @]@     �U@             �B@      2@      @              &@       @     �F@      @     @R@       @              �?      @     �R@     �M@              @@      ,@                      "@      @      @@      @     �O@       @              �?      �?      L@      I@              3@      @      @               @      �?      *@              $@                              @      3@      "@              *@      �?               @                      8@              J@                              �?      E@      ;@              @      �?               @                      *@              5@                                      *@      "@              �?                                              &@              ?@                              �?      =@      2@              @      ,@      @      @              &@     @T@      @      d@      @      �?      @      "@     �P@      >@      @      2@      $@      @       @              @     �N@      @     �X@      @              @      @      F@      :@      @      .@      "@      @       @              @       @             �C@                      @              ,@      *@              @      @                              �?      @              4@                                      @       @               @      @      @       @              @       @              3@                      @              $@      &@              @      �?       @                      �?     �J@      @      N@      @              @      @      >@      *@      @       @              �?                      �?      .@              <@                      �?      @      @      @      @      @      �?      �?                              C@      @      @@      @               @      �?      8@      @       @      @      @              �?              @      4@             �N@              �?               @      6@      @              @      @                              @      1@              L@              �?               @      .@       @               @      �?                                      @              @                                              �?                      @                              @      *@             �I@              �?               @      .@      �?               @                      �?              �?      @              @                                      @       @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�#�UhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �2@)���|�?�	           ��@       	                    @sZ�m��?�           �@                            @y�����?�           `�@                          �0@���?^           ��@������������������������       ��a�Sp�?L            �_@������������������������       �ڎ����?           �{@                           �?q4�Q���?�            �n@������������������������       �bRJxw��?C            �Y@������������������������       �|/)e�!�?\            �a@
                           �?8�\ی��?�            Pq@                           @��ͻ��?Z             c@������������������������       �b�L^E��?-            @R@������������������������       ����Q8�?-             T@                           @��z4���?M             _@������������������������       �J#��PJ�?=            �X@������������������������       �,�wɃ�?             :@                           �?t�.?�?�           �@                          �;@XVf���?           D�@                          �5@ep/���?�           ��@������������������������       �ﰻl+�?7           �~@������������������������       �X*�a!5�?b           �@                           @����?i            �d@������������������������       ��Z����?_            @b@������������������������       ��G�z�?
             4@                            @4u%����?�           ܘ@                            �?D=�Q�?�           p�@������������������������       ����i��?           ��@������������������������       ��[I��?�            @r@                           �?��r�)��?*           �}@������������������������       ��~�t�?W            `a@������������������������       �G���H��?�             u@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      <@     �C@      5@     @^@     ��@      <@     ��@      2@       @      S@      Q@     ��@      �@      "@      p@      S@      @      (@      @      4@     �f@       @     �p@      @      �?     �B@      7@     �j@     �c@      @      S@      M@      @      @      @      ,@      b@      @     �f@      �?              8@      1@     @f@      [@      @      M@     �G@      @      @       @      "@     @[@      @      _@      �?              3@      *@      Y@     �U@      @      D@      .@       @      @              @      3@       @      .@                      @      @      ?@      4@              @      @@      @      �?       @      @     �V@       @     @[@      �?              *@      @     @Q@     �P@      @      B@      &@       @      @      @      @     �A@             �M@                      @      @     �S@      6@              2@      @       @       @              @      7@              .@                      @      @      ;@      (@               @       @              �?      @      �?      (@              F@                      �?      �?     �I@      $@              $@      2@              @      �?      @     �B@      @     @T@      @      �?      *@      @      A@      I@              2@      (@              @      �?      @      ;@      @      >@      @      �?       @      @      6@      <@              "@      &@              �?      �?      @      *@              @      @                      @      &@      .@              @      �?              @              �?      ,@      @      9@              �?       @       @      &@      *@              @      @              �?                      $@      �?     �I@                      &@      �?      (@      6@              "@      @              �?                      @      �?     �G@                      $@      �?      "@      $@              @                                              @              @                      �?              @      (@               @     @`@      5@      ;@      .@     @Y@     �@      4@     ��@      ,@      @     �C@     �F@     �~@     `v@      @     �f@      Q@      &@      ,@      @      N@     @o@      $@     @s@      "@      @      2@      3@      k@      d@             @S@     �H@      $@      (@      @      L@     �l@      $@     @o@       @      @      $@      2@      i@     `a@              O@      ?@      @      @      �?     �H@     �V@      @     �]@      @      @      @      "@     @S@     �M@              :@      2@      @       @      @      @     �a@      @     ``@      @      �?      @      "@      _@      T@              B@      3@      �?       @              @      3@              M@      �?               @      �?      0@      6@              .@      3@      �?       @              @      2@              G@      �?               @      �?      &@      6@              *@                                              �?              (@                                      @                       @      O@      $@      *@       @     �D@     @p@      $@     @�@      @      @      5@      :@     q@     �h@      @     @Z@      G@      @      &@      @      A@     �g@      "@     pu@      @       @      5@      4@      g@     �b@      @     @V@      9@      @      �?      @      4@     �b@      @     �q@       @              &@      1@     �b@     �Y@      @      H@      5@              $@      �?      ,@      D@      @     �O@       @       @      $@      @      A@      G@      �?     �D@      0@      @       @      �?      @      R@      �?      j@      �?      �?              @     @V@     �H@              0@      @                      �?      �?      0@             �Q@              �?              �?      1@      0@              (@      *@      @       @              @      L@      �?     @a@      �?                      @      R@     �@@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�"~hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?a&��j�?�	           ��@       	                     @�&{�G�?I           D�@                            �?zQ��C�?#           L�@                           @&P�f��?           `z@������������������������       �M��l��?�            `h@������������������������       ���Ch��?�            `l@                           @��
yTy�?           h�@������������������������       ��g^F���?�           �@������������������������       �_j����?/             S@
                          �;@U=�g�?�?&           �{@                          �5@I��d�?�            �x@������������������������       ���-!���?�             m@������������������������       ������?f            `d@                           �?�:��X��?*            �I@������������������������       ��ˠT�?	             &@������������������������       �
ףp=
�?!             D@                          �6@Rxj���?S           �@                           @�=� �3�?P           p�@                            @�l���?l           ��@������������������������       ��~�7*�?           �{@������������������������       ������e�?g            �d@                           @��r�1~�?�           ��@������������������������       �q�r���?�            �m@������������������������       ���gƴ��?O           ��@                           @V���"��?           ��@                           �?kFm��?�           0�@������������������������       �2{�69�?Q            �_@������������������������       �4TR�t��?�           @�@������������������������       ����J�?             6@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      4@      ?@      .@      \@     ��@      <@     �@      1@      $@      T@      M@      �@     8�@      9@     �l@     �Z@      ,@      5@      @      R@     �t@      0@     Pz@      (@      @     �A@      A@      t@      k@      $@      `@     �T@      @      0@      @      K@     �n@      ,@     r@      (@      @      8@      <@     �l@     �e@      $@     @Y@      0@      @              �?      4@     @V@      @     �Z@      �?              "@      *@     �R@     �M@      @      6@      $@                      �?      @      K@      �?      J@                      @      @      >@      1@       @      &@      @      @                      *@     �A@      @      K@      �?              @      @      F@      E@      @      &@     �P@      @      0@      @      A@     �c@      $@     �f@      &@      @      .@      .@     �c@     �\@      @     �S@     @P@      @      0@      @     �@@     �b@       @     @c@      &@      @      .@      *@     �b@     �Y@      @     �P@      �?                              �?       @       @      =@                               @      "@      (@              (@      9@      @      @              2@     �T@       @     �`@                      &@      @     @V@      E@              ;@      3@      @      @              0@     @S@       @     @[@                      &@      @     @T@     �C@              9@      &@      @      �?              0@      C@      �?     �Q@                      @      @      D@      2@              4@       @       @      @                     �C@      �?     �C@                      @             �D@      5@              @      @              �?               @      @              7@                              �?       @      @               @                                              �?              @                              �?      @      �?              �?      @              �?               @      @              3@                                      @       @              �?      W@      @      $@      $@      D@     �v@      (@     ��@      @      @     �F@      8@      ~@     �r@      .@     @Y@     �R@       @       @       @      9@      l@      @     pw@      @       @      =@      0@     0s@     �i@      "@     @S@      A@               @       @      $@     @X@             �e@       @               @       @     �d@     @Q@       @      =@      ;@              @              "@     �T@             @]@       @               @       @     �Z@      H@       @      :@      @              �?       @      �?      .@              L@                                      M@      5@              @     �D@       @              @      .@      `@      @     @i@      �?       @      5@       @     �a@      a@      @      H@       @                      �?       @      F@      �?      T@               @      @      @      B@      C@      @      .@     �@@       @              @      *@      U@      @     �^@      �?              2@      @     �Z@     �X@       @     �@@      1@      @       @       @      .@     �`@      @     �q@       @       @      0@       @     �e@     �X@      @      8@      1@      @       @       @      .@     �_@      @     �q@       @       @      0@       @     �d@     �W@      @      8@      �?                              �?      .@      @      B@                      @       @      A@      9@              @      0@      @       @       @      ,@      \@      @      o@       @       @      *@      @     @`@     @Q@      @      2@                                               @              �?                                      "@      @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ%�cDhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �2@ :N�K��?�	           ��@       	                    @�D�^�%�?�           x�@                           �?��y����?�           ��@                           �?q,mҏZ�?�            @t@������������������������       �(f da�?Y            �a@������������������������       �j��fw��?t            �f@                           @�fi}]�?           �x@������������������������       �H�z���?�             n@������������������������       �
�V`���?b            �c@
                           @4�fJ�(�?�            �t@                           @2�ʫK:�?�            �s@������������������������       �9��v���?             I@������������������������       ���'�1,�?�            �p@������������������������       �X�3�R�?             3@                            @l�bGa�?           V�@                           �?d��ú��?�           L�@                           @zX�	�"�?"           H�@������������������������       �D��?���?�            �x@������������������������       �{[y�(�?#           �}@                            �?�"��s�?�           ��@������������������������       �{�Ic �?.           @�@������������������������       ������?�             p@                           �?��M���?           ��@                          �6@S>{@h��?Y            �b@������������������������       ����iL�?0            �S@������������������������       �����L��?)            �Q@                           �?Vq���K�?�           �@������������������������       ��uE���?�            pr@������������������������       ���x,�?�            �y@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @h@     �G@     �B@      >@     �^@     ��@      <@     ��@      1@      .@     �R@      O@     ��@     ��@      4@      p@     @P@      @      (@      1@      :@     �f@      @     �l@      @      @      :@      8@     �j@     �c@      "@     �R@      E@      @       @      *@      *@     �_@      @     �a@      �?              .@      2@     �e@     �Y@      @     �I@      1@              @       @      $@      J@      �?     @R@      �?              @      &@     �L@     �I@      @      :@      @              @              @      ?@              >@      �?              @      &@      2@      2@              .@      *@              @       @      @      5@      �?     �E@                                     �C@     �@@      @      &@      9@      @      �?      @      @     �R@      @     �Q@                       @      @     �\@      J@      @      9@      (@      @              �?      �?     �K@      @      F@                      @      @     @Q@     �A@       @      @      *@       @      �?      @       @      3@              :@                      @      �?      G@      1@       @      3@      7@              @      @      *@     �L@       @     @U@       @      @      &@      @     �D@      L@       @      8@      7@              @      @      (@     �K@       @     @T@       @      @      &@      @     �D@     �F@       @      7@      $@                              �?      @       @      *@                       @               @      @               @      *@              @      @      &@      H@              Q@       @      @      "@      @     �@@      D@       @      5@                                      �?       @              @                                              &@              �?      `@      E@      9@      *@     @X@     P~@      6@     Ȋ@      ,@      (@     �H@      C@     �@     pw@      &@     �f@     �V@      <@      1@      &@     @T@     @v@      1@     x�@      (@       @     �D@      >@     �u@     �q@      $@     �a@     �I@      *@      &@      @     �I@      f@      "@     @k@      @       @      &@      ,@     @\@      \@      @     �S@      8@      @      "@      @      8@     �S@      �?      ]@       @       @      "@      $@      F@      A@              @@      ;@      "@       @              ;@     @X@       @     �Y@      @               @      @     @Q@     �S@      @      G@     �C@      .@      @      @      >@     �f@       @     Ps@      @      @      >@      0@     �m@      e@      @     @P@      >@      *@       @      @      .@     �b@      @      p@      @              0@      $@     @f@     �`@      @     �F@      "@       @      @              .@      =@       @     �I@              @      ,@      @      N@      B@      @      4@     �C@      ,@       @       @      0@      `@      @     �t@       @      @       @       @     �c@     �W@      �?      C@      &@               @              @      9@      @     �B@                                      <@      8@              ,@      @              �?                      ,@      @      6@                                      $@      @              ,@      @              �?              @      &@              .@                                      2@      1@                      <@      ,@      @       @      &@      Z@       @     Pr@       @      @       @       @     @`@     �Q@      �?      8@      6@      @      @              @     �E@       @     @Z@              �?      @              I@     �@@      �?      ,@      @       @       @       @      @     �N@             �g@       @      @      �?       @      T@     �B@              $@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJU�nhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @Xs}|�o�?�	           ��@       	                    �?�8z���?�           ڥ@                           �?=���r�?           ��@                           �?��+���?g             f@������������������������       �
U��6��?*             Q@������������������������       �jko���?=            @[@                          �=@�w
�vk�?�           8�@������������������������       �n���Fx�?�           ��@������������������������       ����|���?             F@
                            �?Z��}BD�?�           ��@                           @������?�           `�@������������������������       ��E���?M           H�@������������������������       ���Fԛn�?�            �m@                           @����n��?�            `u@������������������������       ���[��?�            Pq@������������������������       �����?+            @P@                           �?�u����?�           p�@                           �?�5N����?t            �g@                           @e���KY�?B            @\@������������������������       �t̳|���?7            �U@������������������������       �z�<p��?             :@                          �3@��?�'��?2             S@������������������������       �(��&y��?             =@������������������������       ��o�?            �G@                           �?>+ 	���?5           ��@                          �0@D>��?�             z@������������������������       ��.�?�P�?	             .@������������������������       �#��{���?�            y@                          �2@X��`�?@           �@������������������������       �6�cm�?W            ``@������������������������       �H(t�\��?�            �w@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �l@      8@      A@      @@     �]@     �@      <@     ȑ@      2@      @     �P@     �N@     ��@     �}@      &@     p@     �e@      3@      6@      >@     �W@      �@      5@     �@      (@      @     �M@     �H@     �}@     �v@      $@     �j@      T@       @      4@      .@      M@     �m@      $@     �q@      @      @      ?@      <@      j@      d@       @     �^@      "@      @       @      @      (@      3@       @      L@      �?              &@       @      9@      0@              .@      @              �?              @       @              :@                      @       @      @      $@              @      @      @      �?      @      @      1@       @      >@      �?              @              3@      @              &@     �Q@      @      2@      &@      G@      k@       @     `l@      @      @      4@      :@      g@      b@       @     �Z@     @Q@      @      2@      &@      E@      k@       @     �i@      @      @      4@      :@      f@     �a@       @     @Z@       @                              @      �?              7@                                      @      @               @     �W@      &@       @      .@      B@     �q@      &@      |@      @      �?      <@      5@     �p@     �h@       @      W@     �Q@      "@      �?      *@      4@     `l@      "@     `w@      @              ,@      &@     �j@     �b@       @      N@     �P@      @      �?      &@      0@      f@       @     �q@       @              (@      $@     `f@     �_@             �E@      @       @               @      @     �I@      �?     �W@      �?               @      �?      A@      8@       @      1@      9@       @      �?       @      0@     �J@       @      S@      @      �?      ,@      $@     �K@     �H@              @@      5@       @      �?       @      "@      H@       @      N@      @      �?      $@      $@      B@      G@              9@      @                              @      @              0@                      @              3@      @              @     �K@      @      (@       @      9@     �g@      @     Py@      @      �?      @      (@      l@     �]@      �?     �E@      @              @              @      >@      �?     �M@                      @      �?      A@     �@@              "@      @              @              @      7@              =@                      @      �?      4@      4@              @      @              @               @      2@              0@                      @      �?      2@      1@              @                                      @      @              *@                                       @      @                       @              @               @      @      �?      >@                                      ,@      *@              @       @               @              �?       @      �?      &@                                      @                      @                      �?              �?      @              3@                                       @      *@                     �H@      @      @       @      2@      d@      @     �u@      @      �?      @      &@     �g@     �U@      �?      A@      @@       @      @      �?      (@     �T@      @      `@      @      �?      @      @     �Q@     �G@              5@       @                                      �?              �?                                      @      @              @      >@       @      @      �?      (@     �T@      @     �_@      @      �?      @      @     �P@     �E@              2@      1@      @       @      �?      @     �S@      @     @k@      �?                       @     @^@     �C@      �?      *@      @                      �?              3@              C@                              �?     �I@      (@              @      &@      @       @              @     �M@      @     �f@      �?                      @     �Q@      ;@      �?      $@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�>hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �:@�;v>��?�	           ��@       	                     @NR
�	��?#           �@                           �?��K�~�?�           ��@                          �9@]"�Mz�?�           Ȑ@������������������������       �Y��j��?�           �@������������������������       ��q�q\�?              H@                          �0@��y���?G           ��@������������������������       �ln��s��?2            �S@������������������������       �^�lӶ��?           T�@
                          �0@�=d��s�?;           h�@                           @��'s�	�?             A@������������������������       �V-��?             9@������������������������       ������H�?             "@                          �2@2�~�}�?$           X�@������������������������       �ꍂ;p��?�            �p@������������������������       ��=^1}�?�           �@                            @���g�.�?t           0�@                          �;@�0Ҳ;��?�            �x@                           �?&�R�G}�?<            �X@������������������������       �0Rb�+��?             =@������������������������       ��a����?*            @Q@                           @���/b��?�            �r@������������������������       ��X��b�?�            �i@������������������������       �ʴ�(?�?:            �W@                          �=@"љl��?x             g@                           �?��
ц��?E             Z@������������������������       ��j��=�?            �E@������������������������       �0�R^=d�?-            �N@                           �?�ڬre�?3            @T@������������������������       �N[]G�?            �C@������������������������       ��Q���f�?             E@�t�b�K     h�h4h7K ��h9��R�(KKKK��h��B�        l@      9@      C@      6@     @[@     �@     �@@     4�@      3@      $@     @R@     �N@     X�@     �~@      0@      q@     @h@      0@      A@      4@     �X@     ��@      <@     ��@      0@      @     �Q@      L@     ��@     �z@      ,@      n@     `d@      "@      <@      0@      S@     �z@      5@     ��@      ,@      @     �I@     �G@     pz@     �t@      ,@      h@      U@      @      1@      "@      D@      j@      ,@      j@      $@      �?      0@      @@     @h@     �a@      @      V@     �T@      @      1@      @      D@     �g@      *@     �i@      "@      �?      .@      @@     �g@      a@      @      U@       @                      @              5@      �?      @      �?              �?              @      @              @     �S@      @      &@      @      B@     �k@      @     �v@      @       @     �A@      .@     �l@     �g@      @      Z@      $@                       @              .@              *@                       @       @      3@      $@              @     @Q@      @      &@      @      B@     �i@      @      v@      @       @     �@@      *@     @j@     `f@      @     �X@      ?@      @      @      @      7@     `d@      @     �s@       @      @      3@      "@     �i@     @Y@              H@      �?                              @      @      �?      3@                      �?              �?       @              @                                              �?              2@                      �?              �?       @               @      �?                              @       @      �?      �?                                                              �?      >@      @      @      @      4@      d@      @     `r@       @      @      2@      "@     �i@     �X@             �F@       @               @      @      @     �E@             �S@                       @      @     �T@      1@              ,@      6@      @      @              ,@     @]@      @      k@       @      @      $@      @     @^@     �T@              ?@      ?@      "@      @       @      $@     @T@      @     �j@      @      @      @      @     �]@      M@       @      @@      3@       @       @       @      @      K@      @     ``@       @      �?      @      @     �U@     �E@      �?      <@      @                       @       @      @      �?      :@              �?              �?      <@      3@               @      �?                      �?                              @                                      0@      @              �?       @                      �?       @      @      �?      7@              �?              �?      (@      (@              @      0@       @       @              @     �G@      @     @Z@       @              @      @     �M@      8@      �?      4@      .@       @       @              @      >@      @      Q@       @              @       @      =@      0@      �?      4@      �?                                      1@             �B@                              �?      >@       @                      (@      �?       @              @      ;@             �T@      �?      @              �?      @@      .@      �?      @      @      �?       @                      3@             �J@                                      $@      (@              @                      �?                      @              ;@                                      @      @               @      @      �?      �?                      .@              :@                                      @      @               @      "@                              @       @              >@      �?      @              �?      6@      @      �?               @                              �?      �?              *@                              �?      &@      @      �?              �?                               @      @              1@      �?      @                      &@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�j�&hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?��R��?�	           ��@       	                   �=@�����^�?E           ��@                          �5@�|��d�?           D�@                          �0@`p�����?{           H�@������������������������       ���Cf��?C            �Y@������������������������       �r�&3[��?8           �@                          �8@^�z+��?�           @�@������������������������       �Lj�:!�?�            Pu@������������������������       ���^�U
�?�            0q@
                          �?@���@�c�?5            �U@                            @�q�q�?             H@������������������������       �N�St$�?             9@������������������������       �J��LQ�?             7@                           �?����U�?             C@������������������������       �      �?             8@������������������������       �������?
             ,@                            @}��#*�?l           D�@                           @�r~���?�           ��@                            �?0~�w�?�           Ȅ@������������������������       ���k���?J           �@������������������������       �R�砄��?c            �c@                            �?d�:Fq�?4           @�@������������������������       �|:�L��?�           ��@������������������������       �����?n            �f@                           @��F�e�?�           �@                           �?-k��^?�?g           8�@������������������������       �զ\�L��?�            �y@������������������������       ��S��7�?h            �e@                          �9@�4���c�?$             M@������������������������       ���m(�9�?            �E@������������������������       ��q�q�?	             .@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@      ?@     �G@      ?@      a@     ��@      ;@     d�@      6@      $@     �P@     �Q@     `�@     �~@      4@     �o@     �Y@      2@     �A@      ,@      V@     �s@      *@     �w@      *@      @      ;@      >@      r@      m@      @     �`@     �V@      2@     �A@      ,@     @S@     Ps@      *@     �u@      *@      @      ;@      >@      q@     @l@      @     �`@      P@      *@      :@      @     �O@     @g@      &@     �j@      &@      @      4@      :@     �a@     @_@      @     @U@      @       @       @      �?      $@      (@      @      1@       @       @       @      @      2@      $@      �?      "@      N@      &@      8@      @     �J@     �e@      @     �h@      "@      @      2@      5@     @_@     �\@      @      S@      ;@      @      "@       @      ,@     �^@       @     �`@       @       @      @      @      `@     @Y@       @     �G@       @              @       @      @     �Q@      �?      R@       @       @      @      @     �U@      K@       @      5@      3@      @       @      @      "@      J@      �?      O@                      @              E@     �G@              :@      (@                              &@      @              >@                                      0@      @              @      @                              &@      �?              0@                                      (@      @               @                                      @                      $@                                      @       @               @      @                              @      �?              @                                       @      �?                      "@                                      @              ,@                                      @      @              �?      @                                      @              @                                      @      �?              �?      @                                                       @                                              @                     �[@      *@      (@      1@      H@     �u@      ,@      �@      "@      @      D@      D@     �~@     Pp@      ,@      ^@     @V@      &@      @      *@     �C@      o@      (@     �{@       @       @      C@      >@     `s@     �i@      (@     @X@     �J@      @      @      @      4@     �X@      @     `f@      @               @      2@     �c@     �R@      @      A@      A@      @       @      @      (@      V@      @     �b@      @              @      "@      _@      J@      �?      4@      3@              @      �?       @      $@              >@                      @      "@      @@      7@      @      ,@      B@       @       @      "@      3@     �b@      @     �p@      @       @      >@      (@     @c@     ``@       @     �O@      :@      @      �?      @      &@      _@      @     �m@      @              3@      "@      `@     �X@      @      E@      $@      @      �?       @       @      ;@              <@      �?       @      &@      @      9@     �@@      @      5@      5@       @      @      @      "@      X@       @     @l@      �?      �?       @      $@     �f@     �K@       @      7@      2@      �?      @      @      "@      T@       @     �i@      �?      �?       @      @     �e@      J@       @      5@      *@      �?      @      @      @     �K@       @     �a@      �?      �?      �?      @     �Z@     �F@       @      5@      @               @              @      9@              O@                      �?             �P@      @                      @      �?                              0@              5@                              @       @      @               @      @                                      @              4@                              @      @       @               @              �?                              &@              �?                                      �?      �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJO� hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?;L����?�	           ��@       	                   �<@1y�C`%�?b            �@                            @��Q8>�?           0�@                           @�p'��_�?�           ,�@������������������������       ��x�n�?�           ��@������������������������       �;&����?9             W@                          �6@tD퟉��?.           |@������������������������       ��S�����?�             s@������������������������       � 4gd��?^             b@
                           @�Ezu��?L             _@                           @��>`���?<            �W@������������������������       ���6���?/             Q@������������������������       �p������?             ;@                          @@@����5�?             =@������������������������       �����>4�?
             ,@������������������������       ����ĳ��?             .@                           @#��.���?}           �@                            @a�mv��?e           ��@                           @�;<�)�?�            �@������������������������       ��aW��?S           �@������������������������       �t�y_sj�?h            `d@                           �?]:yȶw�?�             q@������������������������       ��q��D�?h            �d@������������������������       ��!�����?B             [@                           @�j��?           ,�@                          �<@�(��?�           ��@������������������������       ����bX�?�           ��@������������������������       ��βMV:�?I            �]@                            �?{[����?             C@������������������������       �A��?�?             ;@������������������������       �>;n,��?             &@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @j@      ?@      E@      =@     @Y@     p�@      C@     t�@      .@      $@      Q@     �R@     0�@      �@      .@     `o@     �Z@      1@      <@      &@     �N@     0r@      5@     0{@       @      @      A@     �D@     r@      o@      @     �`@     �W@      1@      :@      &@     �L@     �q@      5@     @x@       @      @      @@     �D@     �p@      m@      @      `@     �Q@       @      ,@      $@     �F@     @k@      .@     @p@       @      @      5@     �A@     �e@     �e@      @     �Y@      Q@       @      (@      $@     �D@      j@      ,@      m@       @      @      5@      A@     �c@     �c@      @      W@       @               @              @      $@      �?      ;@                              �?      1@      1@              &@      9@      "@      (@      �?      (@     �O@      @      `@               @      &@      @     �V@     �L@              :@      .@      @      "@      �?      "@      C@      @     @W@               @      "@      @      O@      >@              5@      $@      @      @              @      9@       @     �A@                       @              =@      ;@              @      (@               @              @      $@             �G@                       @              9@      1@              @      @               @              @      $@              C@                       @              4@      @              @      @               @              @      $@              >@                       @               @       @              @       @                                                       @                                      (@      @                      @                                                      "@                                      @      $@                      @                                                      @                                      @      �?                       @                                                      @                                              "@                     �Y@      ,@      ,@      2@      D@     �t@      1@     P�@      @      @      A@     �@@     P|@     �r@      $@     @]@     �O@      @      @      $@      .@      a@      @     `s@      @      @      *@      &@     `l@     �W@      @      H@      K@      @      @       @      &@     �Z@      @     @i@      @              $@      $@      b@     @R@      @      D@     �J@      @       @      @      &@     �T@      @     `a@                      "@      @     �Z@      N@      @      <@      �?               @       @              7@             �O@      @              �?      @      C@      *@              (@      "@              �?       @      @      ?@              [@              @      @      �?     �T@      6@               @      @              �?       @      �?      6@             �P@              @      @      �?      C@      1@               @      @                              @      "@             �D@                                      F@      @                      D@      &@      "@       @      9@     @h@      ,@     @w@      @       @      5@      6@     @l@     �i@      @     @Q@      C@      $@      "@       @      8@     @g@      ,@     �v@      @       @      5@      6@     `k@      h@      @     �P@      B@      $@      "@       @      8@      e@      ,@      s@       @       @      3@      4@     �h@     �g@      @      N@       @                                      2@             �O@      �?               @       @      4@      @              @       @      �?                      �?       @              @                                      @      &@              @      �?      �?                      �?      @              @                                      @      @              @      �?                                      @                                                              @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ+�)NhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx                              @E���5�?�	           ��@       	                    @1m��7��?�           L�@                           �?\<����?B           �@                           @'�Kgå�?�            w@������������������������       �47׀��?�            @r@������������������������       ����	 ��?-            @S@                          �1@�sog��?f           2�@������������������������       �paRC4%�?           �y@������������������������       �^8�xL��?X           �@
                          �;@b� <`i�?�            �q@                           �?�՗Q]�?�            @m@������������������������       �D^�����?            �@@������������������������       ������c�?�             i@                           �?n���?             I@������������������������       ��b�=y�?             9@������������������������       ��+e�X�?             9@                           @Es1mZ�?�           ��@                           �?����@Z�?�           D�@                          �9@���G�\�?           0{@������������������������       �c{���?�            �u@������������������������       ����&���?6            @V@                          �<@<�Q��?�           ��@������������������������       �`���?^           ؀@������������������������       �����?*            �P@������������������������       ��Kh/���?             2@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @h@      ?@      B@      7@     �Y@     ��@      =@     �@      ,@      @     �R@      Q@     ��@     ��@      ,@     �l@     �b@      9@      9@      3@      W@     �@      4@     h�@      &@      @     �P@      N@     p~@      y@      *@     �g@     �a@      9@      5@      2@     @U@     @}@      3@     8�@      "@      @     �N@      K@     `{@     �v@      *@     �e@      0@      �?      @      �?       @      L@       @     �W@                      0@      @     @T@     �H@      @     �A@      .@      �?      @               @     �E@              Q@                      ,@      @     @R@      A@      �?      <@      �?                      �?              *@       @      :@                       @               @      .@       @      @     �_@      8@      1@      1@     @S@     �y@      1@     H�@      "@      @     �F@     �I@     Pv@     �s@      $@     @a@      6@      @      @      @      "@      W@      @     �R@      �?      �?      @      ,@      Q@     �Q@      @      ;@     @Z@      4@      (@      ,@      Q@      t@      (@     �@       @       @      C@     �B@     r@     @n@      @     �[@      @              @      �?      @      E@      �?     �Y@       @              @      @     �H@     �C@              2@      @              @      �?      @     �B@      �?     �R@       @              @      @      B@     �B@              2@      �?              �?              �?      @              0@                                      &@                              @              @      �?      @      A@      �?     �M@       @              @      @      9@     �B@              2@                                              @              ;@                      �?       @      *@       @                                                              @               @                      �?       @      @       @                                                                              3@                                      @                              F@      @      &@      @      &@     �b@      "@     �z@      @      @      @       @     �i@      `@      �?      D@      F@      @      &@      @      &@     �a@      "@     Pz@      @      @      @       @     �i@     @_@      �?      D@      :@      @       @              @     �N@      @      d@       @      �?      @      @      S@     �J@              5@      1@      @      @              @      L@      @     �\@       @      �?      @      @     �N@      E@              3@      "@               @                      @             �F@                                      .@      &@               @      2@      �?      @      @      @     �T@       @     Pp@      �?      @       @      @      `@      R@      �?      3@      1@      �?      @      @       @      Q@       @     �l@                       @      @      ]@      R@      �?      2@      �?                               @      ,@             �@@      �?      @                      (@                      �?                                              @              @                                              @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�^thG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @Z�(��?�	           ��@       	                     @q�X�k��?g           �@                            �?J��k�?#           ��@                           @?����?_           ��@������������������������       ���bM>��?�           ؅@������������������������       ���^�J�?�            �o@                           @����[,�?�            �r@������������������������       ��Y+���?a            �b@������������������������       ���'j���?c             c@
                           �?I���})�?D           ��@                          �6@��L���?�            �r@������������������������       ��wB��|�?v            `f@������������������������       �;��v�?F            @]@                          �0@/�Y�f�?�            �m@������������������������       �"pc�
�?             &@������������������������       ���U&#�?�             l@                           �?7Q���b�?E           ��@                          �;@X�f�f��?=           �@                          �3@��-���?           H�@������������������������       � F>DK�?�            @t@������������������������       ����H��?2           P~@                           @�����?7             V@������������������������       �r3�M�e�?#             M@������������������������       �贁N�?             >@                           �?
?H���?           8�@                          �1@��T���?_           ��@������������������������       ��D̏S�?            �I@������������������������       �    P�?B            �@                           @�v�D{��?�           ؄@������������������������       �� '���?s            @h@������������������������       �r�I$?�?6           �}@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@     �@@      ?@      <@     @[@     0�@      ?@     ��@      6@      "@      T@     @R@     ��@     @      6@      p@     @[@      &@      9@      2@     �H@     �r@      &@     @~@       @      @      ?@     �@@     `w@      i@      @     @_@      W@      "@      3@      0@     �D@     �k@      @     Ps@       @      �?      4@      ?@     `m@     �a@      @     �X@      L@       @      (@      $@      5@      g@      @      p@      @              .@      3@     �g@     �Y@      @      P@      H@       @      "@      @      1@     �`@      @     `e@                      (@      .@     @a@     �U@             �J@       @              @      @      @      J@             @U@      @              @      @     �J@      1@      @      &@      B@      �?      @      @      4@      C@       @     �J@      @      �?      @      (@      F@      D@             �A@      1@      �?      @      @      ,@      @              >@      �?              @      @      6@      7@              4@      3@              @       @      @      ?@       @      7@       @      �?       @       @      6@      1@              .@      1@       @      @       @       @     @S@      @     �e@              @      &@       @     `a@      M@              :@      $@              @       @      @      F@      �?      \@              @      @      �?     �N@      @@              1@      @               @       @      �?     �A@      �?     �J@                       @              E@      7@              (@      @               @              @      "@             �M@              @       @      �?      3@      "@              @      @       @       @              @     �@@      @     �O@                      @      �?     �S@      :@              "@                                               @              "@                                                                      @       @       @              @      ?@      @      K@                      @      �?     �S@      :@              "@     @V@      6@      @      $@      N@     �w@      4@     �@      ,@      @     �H@      D@     �u@     �r@      3@     �`@     �E@      *@      @       @     �A@     �e@      $@      n@       @      @      .@      0@      `@     �_@      (@     @P@     �@@      &@      @       @      A@     �d@      $@     �j@       @      @      ,@      0@     @\@     �\@      &@     �K@      2@      @       @              $@     �I@      @     �V@      �?       @      @      (@      F@      E@      @      @@      .@      @       @       @      8@      ]@      @     �^@      @      �?      "@      @     @Q@     @R@      @      7@      $@       @                      �?      @              <@                      �?              0@      (@      �?      $@       @       @                      �?      @              6@                      �?              @      @      �?      @       @                                                      @                                      &@      @              @      G@      "@       @       @      9@     �i@      $@     �x@      @      �?      A@      8@     �k@      e@      @      Q@      7@      �?      �?      @      (@     �[@       @      f@      @      �?      $@      $@     �X@     �Q@      @      8@       @                              @      @              8@                              �?      @       @       @      @      5@      �?      �?      @      "@      Z@       @      c@      @      �?      $@      "@      W@     @Q@       @      5@      7@       @      �?       @      *@     �W@       @     `k@      �?              8@      ,@     @^@     �X@      @      F@      @       @                      @      9@             �Q@                      @      @     �G@      5@              0@      4@      @      �?       @      $@     @Q@       @     �b@      �?              4@      &@     �R@     @S@      @      <@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��UhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B         
                     @~6�K���?�	           ��@       	                    !@X�>]�?�           �@                          �2@xl�wM	�?�           ƥ@                           @����V�?�           (�@������������������������       ��Ib �2�?a           0�@������������������������       ��$���?�            �k@                            �?���2���?�           ��@������������������������       �>.F3���?�           ��@������������������������       ���ĝ�{�?4           �}@������������������������       �     @�?	             0@                          �:@����S�?�           X�@                           @zX%bB��?E           ��@                           @a�V���?<            �@������������������������       ��ہ2���?�           �@������������������������       ��@�l}�?�            p@������������������������       ��P�n#�?	             1@                           @֚����?y             h@                           �?��b����?k            `e@������������������������       �h���I�?             7@������������������������       ���X��?Z            �b@                           �?�7�A�?             6@������������������������       �r�q��?             (@������������������������       �{�G�z�?             $@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@     �@@      C@      ?@     @\@     ��@     �A@     Ȑ@      .@      @     �T@     �N@     ��@     ��@      7@     pq@     �b@      .@      9@      :@      W@     �~@      @@     p�@      $@      @     @R@      I@      @     �x@      4@     �l@     �b@      .@      9@      :@      W@     �~@      =@     p�@      $@      @     @R@      I@      @     �x@      4@     �l@      O@       @      $@      @      3@     �b@      @      d@              �?      8@      5@      c@      ^@      ,@     �M@      F@       @      @      @      &@     �\@      @      ]@                      2@      2@      ]@      T@      (@     �B@      2@              @               @      A@       @      F@              �?      @      @      B@      D@       @      6@     �U@      *@      .@      5@     @R@     @u@      6@     p�@      $@      @     �H@      =@     �u@     0q@      @      e@      Q@       @      &@      5@      B@     �q@      ,@     0z@      @              C@      1@     �p@      h@      @     �^@      2@      @      @             �B@     �M@       @     �Z@      @      @      &@      (@     �S@     �T@      �?      G@       @                                      @      @                                                      @               @     �G@      2@      *@      @      5@     �e@      @     @x@      @       @      $@      &@      m@     @`@      @     �H@      D@      *@      "@      @      1@     @b@      @     pr@       @       @      $@      "@      i@     �]@      �?      G@      D@      *@      "@      @      1@     �a@      @     `r@       @       @      $@      "@     @h@      ]@      �?      E@      >@      @      "@      @      &@      [@      @     �h@       @       @      @       @      `@     �X@      �?      A@      $@       @               @      @     �A@             @X@                      @      �?     @P@      2@               @                                              @              �?                                      @      @              @      @      @      @              @      ;@             @W@      @                       @      @@      &@       @      @      @       @       @              @      3@             @V@       @                       @      >@      "@       @      @      �?               @              �?      @              @                                       @      @                      @       @                      @      .@             �T@       @                       @      <@      @       @      @              @       @                       @              @      �?                               @       @                              @       @                      @              �?                                       @      �?                                                              @              @      �?                                      �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��UhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�C~֊�?�	           ��@       	                   �1@$g��?&           ��@                            �?���1���?�            Pt@                          �0@|�����?l            �f@������������������������       �e�A�$��?(            �P@������������������������       ��}�c���?D            @]@                            @�<�i�x�?S            �a@������������������������       �`�3�9�?3            @V@������������������������       ��2+��?�?             �J@
                           �?�U�Z���?g           ��@                           �?��Q�&�?z            �h@������������������������       ��������?-             R@������������������������       �w�x��?M            @_@                            @�x��C��?�           ��@������������������������       �j%���4�?           p�@������������������������       ��:Y����?�            `u@                            @�9-~���?a           6�@                            �?~@؜���?�           $�@                          �;@\��0�?           X�@������������������������       ���JA�?�           ��@������������������������       �鵂O�?f            @e@                          �1@�]�i��?�            0w@������������������������       ��Zk����?#             O@������������������������       �Im����?�            Ps@                          �;@��>-��?t           ��@                          �5@�Z��e+�?>           �@������������������������       ���F|Y��?�            �q@������������������������       �Rg0���?�             l@                          @@@[����?6            �T@������������������������       �zDن��?%             K@������������������������       ���>�Q�?             =@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @g@      E@     �@@     �A@      [@     �@      >@     t�@      5@       @     @V@      J@     p�@     �@      3@     @q@      Y@      6@      7@       @     �I@     �s@      ,@     �z@      *@      @      E@      =@     �q@      l@       @     @c@      5@              @              *@      M@      @      L@               @      .@      "@      F@      J@      @     �C@      .@              @              @      9@      @      @@                      @      @      >@      C@       @      .@                      �?              @      $@      @      @                              @      (@      3@              @      .@               @               @      .@       @      9@                      @       @      2@      3@       @      $@      @              @               @     �@@              8@               @      $@       @      ,@      ,@       @      8@       @              �?              @      8@              &@               @      @      �?      $@      @       @      1@      @               @              �?      "@              *@                      @      �?      @       @              @     �S@      6@      1@       @      C@     �o@       @      w@      *@       @      ;@      4@     �m@     �e@      @     �\@      @      �?              @      "@      >@             �O@       @              @              C@      3@              ,@      �?      �?                      @      @              :@      @               @              &@      "@              "@      @                      @      @      8@             �B@      @              @              ;@      $@              @     �R@      5@      1@      @      =@      l@       @     s@      @       @      5@      4@     �h@     @c@      @     @Y@      O@      1@      *@      @      4@     `d@      @     `h@       @      �?      ,@      2@     �`@     @\@      @     �T@      (@      @      @      �?      "@      O@      @     �[@      @      �?      @       @     @P@     �D@              2@     �U@      4@      $@      ;@     �L@     �v@      0@     ��@       @      @     �G@      7@     `{@     �q@      &@     �^@     �R@      1@       @      2@      J@     `p@      0@     �z@      @      @      G@      2@     �s@     @l@      $@     �[@     �L@      ,@      �?      &@      9@     `k@      *@     �v@      @              =@      &@     �n@     �d@      @      R@      J@      &@      �?      @      7@     �f@      (@     �r@      @              <@      $@      l@      c@      @     �L@      @      @              @       @      B@      �?     �O@      @              �?      �?      7@      &@              .@      2@      @      @      @      ;@     �E@      @     �N@              @      1@      @     �Q@      O@      @      C@      @               @      @              0@              @                      @      @      @      .@      �?      �?      .@      @      @       @      ;@      ;@      @      K@              @      *@      @     @P@     �G@      @     �B@      &@      @       @      "@      @     �X@             �p@      �?      �?      �?      @     @^@      K@      �?      (@      $@      @       @      "@      @     �R@             @l@      �?              �?      @     �[@     �J@      �?      (@      @               @      "@       @      B@              a@      �?                       @      J@      A@              @      @      @                      �?      C@             @V@                      �?      @     �M@      3@      �?      @      �?                               @      9@             �E@              �?                      $@      �?                                                              6@              ;@                                      @      �?                      �?                               @      @              0@              �?                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJO��-hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @M-�=��?�	           ��@       	                     �?���Ϭ��?�           ��@                           @��&�ޏ�?-           L�@                            �?mI��Õ�?�           З@������������������������       �s��^��?�           ��@������������������������       �v�S�:!�?�           ��@                          �@@O��FA�?\           ��@������������������������       �T����6�?T           �@������������������������       �6�h$��?             .@
                          �0@�HZ��?�           �@                           @6��D��?             E@������������������������       �      �?              @������������������������       �d��E���?             A@                           �?�~�F5��?�           ��@������������������������       �t}:k��?}            �i@������������������������       ���4���?           @z@                           �?8�Rp~x�?�           �@                           @���ð��?:           �@                           @��)t��?           �z@������������������������       ��'���?�            @w@������������������������       �2��t��?&            �L@                           �?"J��:�?4            @T@������������������������       �,R�n��?             B@������������������������       ���`d�k�?            �F@                           @j2t�C[�?�           @�@                           @y1�R��?8           �@������������������������       �Ϝ����?            z@������������������������       �'�Tk��?5            �V@                           @��B�(��?\            �a@������������������������       ��J�fj�?L            �[@������������������������       ��8���?             =@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      ?@      F@      6@      Y@     �@      E@     @�@      5@       @     �T@     @Q@     І@     ��@      :@     p@     @b@      5@      <@      1@     �T@     �|@     �A@     H�@      1@      @     @R@      M@     �}@     �x@      6@      i@     �[@      .@      4@      .@     �K@     0v@      8@     ��@       @       @     �F@      E@     �w@     0q@      *@      `@     �U@      "@      .@      *@      I@     �q@      .@     �{@      @             �A@      >@     �o@     `f@      &@      X@      >@      �?      �?      @      4@      a@      (@      n@      @              &@      1@     @`@      U@      @     �B@     �L@       @      ,@      @      >@     `b@      @      i@      @              8@      *@     @_@     �W@      @     �M@      8@      @      @       @      @      R@      "@     �c@       @       @      $@      (@     �_@      X@       @     �@@      8@      @      @       @      @     �Q@      "@     `c@       @       @      $@      &@     �_@     @U@       @     �@@                                               @              �?                              �?              &@                     �A@      @       @       @      <@     �Z@      &@     @]@      "@      @      <@      0@     @X@      ^@      "@      R@      �?                              �?      (@      �?      @                              @      @      ,@              �?                                      �?      @                                              @              �?                      �?                                      "@      �?      @                                      @      *@              �?      A@      @       @       @      ;@     �W@      $@     @\@      "@      @      <@      *@      W@     �Z@      "@     �Q@      ,@       @      �?       @      $@      :@              =@      @      �?       @      @      B@      F@      @      :@      4@      @      @              1@     @Q@      $@      U@       @      @      :@      $@      L@      O@      @     �F@     �N@      $@      0@      @      1@     �e@      @     px@      @       @      $@      &@     �o@      a@      @      L@      C@      @      &@      �?      &@     �R@      @     `b@      �?       @       @      @      X@     @P@      �?     �B@      ?@       @      $@      �?      &@     �N@      @      ^@      �?               @      @     �U@      N@      �?      <@      :@       @      $@      �?      $@     �L@      @     �Y@                       @      @      R@     �I@              8@      @                              �?      @      �?      1@      �?                              ,@      "@      �?      @      @      @      �?                      *@      @      ;@               @                      $@      @              "@      @      �?      �?                       @              0@               @                      @       @              �?       @      @                              &@      @      &@                                      @      @               @      7@      @      @      @      @     @Y@             �n@      @               @      @     �c@      R@      @      3@      5@       @      @      @      @      O@              i@                      �?      @     @a@      H@              1@      0@       @       @      @      @     �G@              e@                      �?      @     �]@     �B@              1@      @              @               @      .@              @@                               @      4@      &@                       @       @                      �?     �C@              F@      @              �?      �?      2@      8@      @       @       @      �?                      �?      @@              C@                              �?      2@      .@      @                      �?                              @              @      @              �?                      "@               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�<�
hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @�Z��{�?�	           ��@       	                     @�~��s�?8           ��@                          �?@*9��?��?           ��@                           �?����?�           �@������������������������       ���T�q3�?�            �q@������������������������       �|0L����?<           ��@                           �?�Z=;n�?             F@������������������������       ��(��0�?             9@������������������������       ���a_j�?             3@
                          �2@�iJ��?+           P�@                           �?D����?�            �q@������������������������       �݃QNZ��?O             _@������������������������       ��Q`؈��?^            �c@                          �;@����?~           x�@������������������������       �.؂-��?7            ~@������������������������       ����@��?G            �[@                            @��O¿}�?�           ��@                          �;@���4���?�           ��@                            �?�֙��9�?�           h�@������������������������       ���\��?F           �~@������������������������       ���:��?b            @d@                          �@@�T�6|��?=             Z@������������������������       �l �&��?7             W@������������������������       �r�q��?             (@                           �?�hZ_�?�             p@                           @ �͜�%�?A            @Z@������������������������       ��3ot`�?2            @T@������������������������       ���8��8�?             8@                          �4@S��X�?Z             c@������������������������       �L�/�V�?             �J@������������������������       ��Q����?:             Y@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @i@      >@      F@      5@     @_@     (�@      :@     ��@      5@      "@     �R@     �Q@     ȇ@     �~@      .@     �o@     @e@      .@      @@      ,@      Z@     ~@      1@     ��@       @      @     �N@      E@     @�@      u@      (@     @g@     �`@      &@      6@      "@     �T@     @v@      &@      �@      @      @     �I@     �C@     �v@     �o@      (@     �b@     ``@      &@      6@      "@     �T@     �u@      &@     �~@      @      @     �I@      C@     �v@     �o@      "@     �b@      (@      �?      �?      �?      1@      C@              Q@                      .@      @     �I@      C@      �?      B@     �]@      $@      5@       @     �P@     ps@      &@     pz@      @      @      B@     �@@     �s@      k@       @     �\@       @                                      @              9@      �?                      �?      @      �?      @      �?      �?                                      @              3@                                      �?                              �?                                      @              @      �?                      �?       @      �?      @      �?     �B@      @      $@      @      5@     @_@      @     �s@      @       @      $@      @     @k@     @T@             �A@      "@              @      @      @      C@             �T@                       @       @      X@      ;@              (@      @              @              @      8@              7@                       @      �?      C@      0@              @      @              �?      @       @      ,@              N@                              �?      M@      &@              @      <@      @      @       @      ,@     �U@      @     �l@      @       @       @      �?     �^@      K@              7@      8@      @      @       @      "@     �S@      @     �e@      @               @             @Y@      H@              4@      @              @              @       @              M@               @              �?      5@      @              @      @@      .@      (@      @      5@     �d@      "@     �r@      *@      @      ,@      <@      f@     `c@      @     �P@      ;@      "@      $@      @      3@     �[@       @      j@      @       @      *@      7@     �`@     @^@       @      M@      ;@      "@      $@      @      2@     �X@       @     �c@      @       @      (@      6@     @\@     �Z@       @     �K@      4@      "@      @      @      ,@      T@      @      `@      @       @      @      $@     @V@     �Q@              D@      @              @              @      2@      �?      =@      @              @      (@      8@     �A@       @      .@                                      �?      (@             �I@                      �?      �?      4@      .@              @                                      �?      (@             �H@                      �?              4@      @              @                                                               @                              �?              "@                      @      @       @               @      K@      �?     �U@      @      �?      �?      @      F@      A@      �?       @      @       @       @              �?      3@      �?      D@      @      �?              @      .@      &@              @      @       @       @                      *@      �?     �A@      @      �?              @       @       @               @      �?                              �?      @              @                                      @      @              �?      �?      @                      �?     �A@             �G@      @              �?       @      =@      7@      �?      @               @                      �?      $@              7@                      �?              &@      @                      �?       @                              9@              8@      @                       @      2@      2@      �?      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�c&hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @ْ�p?��?�	           ��@                           �?nH-Z�?�           ��@                           @
W�ٮ�?�           ��@                            �?˪Z���?�           \�@������������������������       �)3u��?�             x@������������������������       �خ�TQ�?�           ��@������������������������       ��ˠT�?             &@                            �?�Ɨ~�{�?�           p�@	       
                    !@�������?
           ��@������������������������       ������?           ��@������������������������       �X�<ݚ�?             "@                           @@5�&��?�            �v@������������������������       ���v���?�            �k@������������������������       �J �f32�?Z            @b@                           �?��{8��?�           ,�@                           �?b�P.�?0           �@                          �1@y
�=?�?n            �f@������������������������       �^�:|z�?             5@������������������������       �
³a8{�?b            @d@                          �<@��:��r�?�            Pt@������������������������       ���]���?�            `q@������������������������       ��o[��?            �G@                           @h����?z           x�@                           @u����?�            �w@������������������������       �������?�            �u@������������������������       �     ��?             @@                           �?7u�׃��?�            @j@������������������������       �l� {�/�?             A@������������������������       ��4_���?r             f@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      9@      H@      4@     �[@     ��@     �B@     (�@      6@      (@      W@     �M@     Ȇ@     @@      0@     pq@     `c@      2@     �A@      ,@     �T@     �~@      >@     ��@      1@      "@      T@     �I@     �~@     �w@      0@     �m@     �Q@      &@      9@       @      M@     �j@      ,@     �o@      (@      @     �@@      ?@     @g@      b@      @      ]@     �Q@      &@      9@       @     �K@     �j@      *@     �o@      (@      @     �@@      ?@     @g@     �a@      @     @\@      1@      �?       @      @      *@     @S@      @      Y@      �?              @      ,@     �Q@     �F@       @      =@      K@      $@      7@      @      E@      a@      "@      c@      &@      @      :@      1@     �\@      X@      @      U@                                      @      �?      �?                                                      @              @      U@      @      $@      @      8@     `q@      0@     0|@      @      @     �G@      4@     @s@     �m@      "@     �^@      K@      @      @      @      0@     �l@      (@      x@      @              8@      .@     0p@     �e@      @      Q@      K@      @      @      @      0@     �k@      (@     x@      @              8@      .@     0p@     �e@      @      Q@                                              @              �?                                               @                      >@      �?      @               @     �H@      @     @P@              @      7@      @     �H@     �N@      @      K@      :@      �?      @              @     �A@      �?     �B@              @       @      @     �B@      @@       @      7@      @              @              �?      ,@      @      <@               @      .@      �?      (@      =@      @      ?@     �H@      @      *@      @      =@      e@      @     �x@      @      @      (@       @     `m@      ^@             �D@      D@      @      @              1@     �U@      @      c@      �?      �?      @      @     @Y@     �L@              9@      1@       @      @              @      A@      @      A@                      @      �?      I@      7@              "@       @               @                      $@                                                      @                      �?      .@       @      �?              @      8@      @      A@                      @      �?      F@      7@               @      7@      @      @              *@      J@       @     �]@      �?      �?      @       @     �I@      A@              0@      (@      @      @              "@     �I@       @      X@              �?      @       @     �G@     �@@              ,@      &@                              @      �?              7@      �?                              @      �?               @      "@       @      @      @      (@     �T@       @     @n@      @       @      @      @     �`@     �O@              0@      @      �?       @      @      @      D@             `d@      �?       @      @             @Z@      ?@              0@      @      �?       @      @      @     �C@             `a@      �?       @      @             �X@      ?@              0@      �?                                      �?              8@                                      @                              @      �?      @              @     �E@       @     �S@      @               @      @      =@      @@                      @              @              @      �?       @      &@                                      @      @                       @      �?                              E@              Q@      @               @      @      :@      ;@                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJgH�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @e��o\u�?�	           ��@       	                     �?Xs>u��?           Υ@                            �?����]��?Q           ��@                          �;@l��"�?�           L�@������������������������       �3���N�?R           ��@������������������������       �@�
L���?R             `@                          �0@^��z�?�           ܐ@������������������������       �t�û��?(            @Q@������������������������       ����6��?�           ��@
                          �1@<A�С~�?�           �@                           @���+m��?W            �`@������������������������       �\l�<,U�?*            �N@������������������������       ���[�?-            �R@                           �?8��]Q�?Y           ��@������������������������       �������?�            �l@������������������������       ��l$Y�Q�?�            �r@                           �?%��B���?�           ��@                           @T[�_�
�?7           �}@                           @���E�?�            0t@������������������������       �>��l���?�            �m@������������������������       ���$��?4            �U@                           @֙N���?h            �c@������������������������       �<#��cl�?T            @^@������������������������       ���˰"��?            �A@                          �@@?�-Ƈ��?�           �@                           @���^��?�           ��@������������������������       ��3x���?'           �|@������������������������       �b�a��?e             e@������������������������       �*D>��?             *@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        f@      ;@     �C@      5@     �[@     ��@      ?@     ��@      :@      $@     @V@      P@     H�@     (�@      3@      o@     `a@      2@      =@      4@     @V@     �@      9@     ��@      4@      "@     �Q@     �K@     �}@     �w@      3@     �i@     @Z@      (@      8@      0@      M@      y@      4@     H�@      *@       @     �L@     �B@     �w@     �o@      .@     �a@     �L@       @      @      (@      <@     �h@      &@     `s@      @              *@      1@     `h@     `a@      @     �E@      K@       @      @      (@      8@     �f@      $@     �o@      @              "@      1@     �e@     @_@      @     �A@      @                              @      1@      �?      L@      �?              @              5@      ,@               @      H@      @      5@      @      >@     �i@      "@     0q@       @       @      F@      4@     @g@     �\@      &@     �X@       @              @               @      "@              @       @              @       @      6@       @               @      G@      @      1@      @      <@     `h@      "@     �p@      @       @     �D@      2@     �d@     �Z@      &@     �V@      A@      @      @      @      ?@     @[@      @      a@      @      @      ,@      2@     @X@     �_@      @     @P@      "@      @      �?              �?      A@      �?      $@               @      @      @      ,@      ?@       @      3@      �?      @                      �?      3@              @                       @      @      @      @       @      *@       @              �?                      .@      �?      @               @      �?      �?       @      8@              @      9@      @      @      @      >@     �R@      @     �_@      @      @      &@      *@     �T@     �W@       @      G@       @      �?      �?       @      &@     �C@       @     �J@      @       @      @       @      >@     �H@      �?      .@      1@       @      @       @      3@      B@       @     �R@      �?      @       @      @     �J@      G@      �?      ?@     �B@      "@      $@      �?      5@     �f@      @     `y@      @      �?      2@      "@     `m@     @a@              E@      5@      @       @              (@     @R@      @     �a@      @              "@      @     �Z@      Q@              8@      1@              @              "@      M@       @      T@                      @       @     �S@      E@              5@      ,@              @              @      C@       @     @P@                      @             �N@      ;@              ,@      @                              @      4@              .@                               @      2@      .@              @      @      @      �?              @      .@       @      O@      @              @       @      ;@      :@              @      @      @      �?               @      ,@       @      E@      @                       @      3@      9@              @              �?                      �?      �?              4@                      @               @      �?                      0@      @       @      �?      "@     �[@       @     �p@       @      �?      "@      @      `@     �Q@              2@      .@      @       @      �?      "@     �[@       @     0p@       @      �?      "@      @     �^@     �Q@              2@      *@      �?       @      �?      @     �P@       @     `i@       @      �?      @      @      W@      F@              1@       @      @                       @     �E@              L@                       @       @      >@      :@              �?      �?                                                      @                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��'hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx                             �?�����?�	           ��@       	                    @�y����?L           h�@                           �?�۰���?@           �@                           �??���l��?t           ��@������������������������       ��@��B��?�            p@������������������������       �6��w��?�            `u@                           �?˱C;��?�           ��@������������������������       �l�~Oh�?           �z@������������������������       ���(x���?�           �@
                          �5@�KM�]�?             3@������������������������       �F]t�E�?             &@������������������������       �      �?              @                            @@�ZҶ��?V           ޠ@                           !@`�eG
q�?�           ��@                           @�Z���o�?�           ��@������������������������       ��:SZ΋�?�           ��@������������������������       ����qs��?�            @x@������������������������       ��'}�'}�?             .@                          �5@8<KQ��?�           ��@                           @o=��ڛ�?�            �s@������������������������       ��Z��t�?�            �j@������������������������       �������?@            @X@                           @SCp�j��?�            �s@������������������������       ��C����?�            �q@������������������������       �ݾ�z�<�?             :@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@      =@      =@      9@      U@     X�@     �F@     (�@      4@       @     @R@     @P@     ��@     �@      .@     �p@     �Z@      0@      7@      ,@      J@     �u@      9@     �y@      (@      @     �A@      >@     0s@      l@       @     `a@     �Z@      0@      7@      ,@     �I@     Pu@      7@     �y@      (@      @     �A@      >@     0s@     �k@       @     �`@     �@@      @      .@       @      3@     �[@      @     `d@      @      �?      3@      @     @W@      O@       @      L@      $@              @      �?       @      B@      �?     @S@      @              .@      @     �I@      6@       @      5@      7@      @       @      �?      &@     �R@      @     �U@      @      �?      @      �?      E@      D@             �A@     @R@      "@       @      (@      @@     �l@      1@     �n@      @      @      0@      :@     �j@     �c@      @     �S@      ?@      @      �?      $@      .@     �V@      @      R@       @       @      @      "@     @S@     @Q@       @     �@@      E@      @      @       @      1@     �a@      $@     �e@      @       @      &@      1@      a@     �V@      @     �F@      �?                              �?      @       @                                                      @              @                                              @       @                                                       @              @      �?                              �?      @                                                              �?              �?     �Z@      *@      @      &@      @@     �t@      4@     ��@       @      @      C@     �A@     �{@     �q@      @      `@     @W@      &@      @      @      =@     �n@      2@     �{@      @      �?      B@      >@     �q@     �j@      @      [@     @W@      &@      @      @      =@     `m@      2@     �{@      @      �?      B@      >@     �q@     @j@      @     �Z@      T@      @      @      @      2@     `f@      0@      s@      @      �?      <@      4@     �k@     �e@      @      P@      *@      @      �?       @      &@      L@       @     `a@                       @      $@     �N@     �A@       @     �E@                                              "@               @                                              @              �?      *@       @       @      @      @     �V@       @     @n@       @       @       @      @      d@     @Q@      �?      5@      @      �?       @      @      �?      F@       @     �Y@       @                      @      W@      C@              &@      @               @      @      �?      :@             �O@       @                       @     �R@      9@              "@       @      �?                              2@       @     �C@                               @      2@      *@               @      @      �?                       @     �G@             �a@               @       @      �?     @Q@      ?@      �?      $@       @                               @      D@             ``@               @       @      �?     @P@      >@      �?      $@      @      �?                              @              "@                                      @      �?                �t�bub�     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��"hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?����}�?�	           ��@       	                     @�3��%�?N           ��@                           �?�g��Zr�?
           ��@                          �0@o�l�5�?c            �a@������������������������       �      �?              @������������������������       ��k%���?]            �`@                          �;@|�e�d�?�           h�@������������������������       �N���m�?n           ��@������������������������       �d��Ü�?9            �V@
                          �<@�F1'
U�?D           8�@                           @�ձ�'k�?*           �}@������������������������       �����~�?�             x@������������������������       ���l�!�?8            @W@                           @�p=
ף�?             D@������������������������       �d���?             ;@������������������������       �.y0��k�?             *@                           @`xע���?Q           2�@                           �?MZ���~�?8           ��@                            @�^��ڊ�?`           H�@������������������������       ��!/��3�?           �{@������������������������       ���꟣��?[            �a@                            @@ժ�U�?�            `u@������������������������       ��j�"�?�            �l@������������������������       ��a�����?G            �\@                           !@v@Rܧ��?           �@                           @���1��?           ��@������������������������       ��T�x?��?�            �@������������������������       � �����?W           X�@������������������������       ��.�?��?
             .@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      C@      C@      <@     �Y@      �@      7@     ��@      *@      @      V@     @P@     (�@      �@      1@     q@     �X@      .@      6@      *@      M@     Ps@      .@     �y@       @      @      H@      A@     �q@     �n@      @      a@     �P@      $@      1@      *@      F@     �i@      *@     �p@      @      @      B@      <@     �g@     �e@      @     @[@      $@               @      �?      @      $@      @     �D@      @              "@       @      6@      2@              .@                      �?              �?                                                              �?      @                      $@              �?      �?      @      $@      @     �D@      @              "@       @      5@      *@              .@     �L@      $@      .@      (@      D@     `h@      "@     �l@       @      @      ;@      :@      e@     �c@      @     �W@     �J@       @      ,@      (@     �A@     `g@      "@     `h@       @      @      7@      :@     �c@     �a@      @     �T@      @       @      �?              @       @              A@                      @              "@      *@              &@      @@      @      @              ,@      Z@       @     �a@      �?              (@      @      X@     @R@              ;@      >@      @      @              (@     @Y@       @     �^@                      (@      @     �V@     �Q@              :@      8@      @      @              "@     �U@      �?     �U@                      $@       @     �S@     �M@              6@      @      �?                      @      .@      �?      B@                       @       @      (@      &@              @       @                               @      @              4@      �?                       @      @      @              �?      �?                               @      @              "@      �?                       @      @       @              �?      �?                                                      &@                                              �?                     �X@      7@      0@      .@     �F@     �t@       @     X�@      @       @      D@      ?@     p|@     �p@      &@      a@     �G@      &@       @      @      :@     �`@      �?     �r@              �?      @      &@     �l@     �V@      @      J@      >@      @      @       @      .@     �T@              g@                      @       @     @b@      Q@      @      B@      <@      @      @      �?      (@     �Q@             �^@                      @       @      Z@      I@      @      @@       @                      �?      @      &@             �N@                                      E@      2@              @      1@       @      @      �?      &@      J@      �?      ]@              �?      @      @     �T@      7@       @      0@      *@       @      @      �?       @      B@      �?      P@                       @       @      M@      0@       @      ,@      @               @              @      0@              J@              �?      �?      �?      9@      @               @     �I@      (@       @      (@      3@     �h@      @     �y@      @      �?      A@      4@     @l@     @f@      @     @U@     �I@      (@       @      (@      3@     �g@      @     �y@      @      �?      A@      4@      l@     @f@      @     @U@     �A@      @      @      @      .@     �]@      @     �m@      @              .@      $@     �X@     �W@      @     �H@      0@      @      �?      @      @     @Q@      @     �e@      �?      �?      3@      $@     �_@     �T@              B@                                              "@              @                                      �?                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJr��8hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�d�ۀ�?�	           ��@       	                     @���pW/�?;           0�@                           @3ā�H�?           ��@                          �?@�����?�           �@������������������������       �ח�<��?�           ��@������������������������       �zv�X�?             6@                           @�_JB2�?7            �W@������������������������       �>M\kz��?1            @U@������������������������       ��������?             $@
                           @P��h�?,           �~@                           �?�l>ĕ��?�            �t@������������������������       ����1�N�?5            @T@������������������������       �fj�!��?�            @o@                           @�}�s��?Z            �c@������������������������       �0�|���?-            �S@������������������������       ��{E��?-            �S@                           �?������?g           ��@                          �3@���e�?�            pu@                          �0@�F��<�?Q            �^@������������������������       �s
^N���?
             ,@������������������������       ���}*_��?G             [@                            �?ƵHPS!�?�            �k@������������������������       �|��U�=�?)            �P@������������������������       ��M�=��?a            `c@                          �;@��$����?�           ��@                            @�N����?�            �@������������������������       �d�eH��?�           ��@������������������������       �CbΊ��?            }@                           @I���?�            �k@������������������������       ��U6A3x�?z            �g@������������������������       ���QN�?             ?@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @i@      ?@      C@      >@     @Z@     0�@      7@     А@      0@       @      S@      R@     ȇ@     �@      2@     �m@      Y@      6@     �A@      1@     �Q@     0u@      (@     Py@      (@      �?      C@      B@     �r@     `l@      @     �]@      O@      ,@      <@      1@      N@      n@      "@      p@      "@              @@      ?@     �j@     �e@      @     �X@      O@      ,@      :@      1@     �L@      m@      @      l@       @              @@      >@     �h@      c@      @     �V@      N@      ,@      :@      1@     �L@     �l@      @     �j@       @              @@      >@     �h@     `b@      @     �V@       @                                      @              &@                                              @                                       @              @      "@       @     �@@      �?                      �?      .@      5@               @                       @              @       @              @@      �?                      �?      ,@      3@              @                                              �?       @      �?                                      �?       @              @      C@       @      @              $@     �X@      @     `b@      @      �?      @      @     �V@      K@              3@     �A@      @      @              @     �R@       @     �T@      @      �?      @      @      L@     �C@              (@      "@              �?              @      7@              ,@                      @              *@      *@               @      :@      @      @              @     �I@       @      Q@      @      �?              @     �E@      :@              $@      @       @      �?              @      8@      �?     @P@                      @              A@      .@              @       @      �?                               @              C@                                      6@      @              @      �?      �?      �?              @      0@      �?      ;@                      @              (@      $@              @     �Y@      "@      @      *@     �A@     0w@      &@     ��@      @      �?      C@      B@     �|@      r@      (@      ^@      2@       @              �?       @      N@      �?     �T@                      @      �?     �R@     �N@      @      9@      $@                              @      *@      �?     �A@                      @              =@      ,@      @      &@      @                                       @              �?                                      @       @               @      @                              @      &@      �?      A@                      @              :@      (@      @      "@       @       @              �?      @     �G@             �G@                      @      �?     �F@     �G@              ,@      @                               @      1@              4@                                      (@      @              @      @       @              �?      @      >@              ;@                      @      �?     �@@      D@              "@      U@      @      @      (@      ;@     ps@      $@     h�@      @      �?      ?@     �A@     x@     `l@      "@     �W@      T@      @      @      (@      :@     Pp@      "@     �~@      �?      �?      ;@      ?@     �u@      k@      @     @V@      N@      @      @      "@      8@     �g@       @     �r@      �?      �?      7@      ;@     �m@     `e@      @     @S@      4@       @              @       @     �Q@      �?     �g@                      @      @     �[@     �F@              (@      @                              �?      I@      �?     @Y@      @              @      @     �A@      &@       @      @      @                              �?      I@      �?     �S@      @               @      @      ?@      $@       @      @                                                              7@                       @      �?      @      �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�BhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�2-��x�?�	           ��@       	                   �:@/�����?�           ��@                           �?0YX��?�           ��@                            �?vĥ�
��?�           ��@������������������������       �~�ቌ�?�            �u@������������������������       ���LL���?�           ��@                          �0@�l�4@��?V           ��@������������������������       �@�(ݾ��?2            �S@������������������������       ��C��?$           l�@
                          �<@�8��8��?�             x@                           @樈/H}�?p            �f@������������������������       ���J(�'�?M            ``@������������������������       �R���
�?#            �H@                           �?&5DSb�?�            �i@������������������������       ������q�?            �E@������������������������       ���+7��?f             d@                           �?ܶ����?�           ȑ@                          �1@-s�[")�?J           @�@                           @���<U"�?0            �S@������������������������       �     ��?&             P@������������������������       ��|�j��?
             .@                          �=@<�*���?           �}@������������������������       ���eJ���?           �z@������������������������       �|z3���?             E@                           @,_t'�}�?p           P�@                          �?@��t���?           |@������������������������       �)�dU��?	           �z@������������������������       ��Q����?             9@                          �=@d�5����?W             a@������������������������       ��#��?N            @^@������������������������       �     ��?	             0@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      ?@      E@      ;@     @X@     P�@      B@     ԑ@      4@      $@     �Q@      O@     H�@     H�@      6@     @o@      e@      7@     �@@      8@     @T@     p{@      <@     ��@      ,@      "@      K@     �J@     P@     @x@      2@     �j@      c@      2@      ?@      4@     �R@     �w@      ;@     �@      &@      "@     �F@      I@     �y@     0v@      0@     �g@      Q@      $@      9@      @     �H@      f@      &@     �m@      &@      @      0@      ?@     �e@      b@      @     �W@      6@      �?      @      �?      .@      N@      �?     @Y@       @              @      *@     �L@      G@      �?      5@      G@      "@      6@      @      A@      ]@      $@      a@      "@      @      *@      2@     �]@     �X@      @     �R@      U@       @      @      *@      9@     �i@      0@     �v@               @      =@      3@     @m@     `j@      "@     �W@      @                      �?              4@              &@                      �?      @      0@      $@               @     @S@       @      @      (@      9@      g@      0@     @v@               @      <@      .@     @k@      i@      "@     �U@      1@      @       @      @      @     �M@      �?     �^@      @              "@      @      W@     �@@       @      9@      &@      @              @      @      :@      �?     �H@       @               @              L@      $@              "@      @      @              @      @      4@              ?@                       @              G@      "@              @      @                              �?      @      �?      2@       @                              $@      �?              @      @      �?       @              �?     �@@             @R@      �?              @      @      B@      7@       @      0@      @                                      &@              "@                      �?      �?      @      @              @      @      �?       @              �?      6@              P@      �?              @       @      >@      1@       @      $@      J@       @      "@      @      0@     `f@       @     �y@      @      �?      0@      "@     �n@     �`@      @      B@      A@      @      @      �?      &@     �X@      @     �d@      @              *@      @     @[@      O@       @      <@      @      �?                      @      (@       @      4@                      @      �?      @      "@              .@      @                              @       @              0@                      @              @      @              .@              �?                      �?      @       @      @                              �?               @                      >@      @      @      �?      @     �U@      @     `b@      @               @      @     �Y@     �J@       @      *@      4@      @      @      �?      @     �T@      @     �`@      @               @       @     �W@     �I@              *@      $@                               @      @              (@       @                      �?       @       @       @              2@       @      @       @      @     @T@       @     �n@      �?      �?      @      @     �`@     �Q@       @       @      ,@      �?      @       @      @     �H@       @     �i@              �?       @      @     �Y@     �H@               @      (@      �?      @       @       @      H@       @     �g@                       @      @     @Y@     �H@               @       @                              @      �?              0@              �?                       @                              @      �?                              @@              D@      �?              �?       @      @@      6@       @              @      �?                              >@              >@                      �?       @      =@      6@       @                                                       @              $@      �?                              @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ;�>whG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @�#��ܛ�?�	           ��@       	                   �;@pƩ��?�           �@                           �?���.�?7           ʣ@                          �1@��"7���?�           �@������������������������       �n+,����?�            0p@������������������������       �w2o�]s�?<           �@                           �?�;�Č��?^           ��@������������������������       �,�kW�M�?           �{@������������������������       ��n�W���?A           @�@
                           @��X����?�            @r@                          �?@�ګH9�?�            �j@������������������������       �/�~�@�?l            �c@������������������������       �������?              L@                           @�f醇�?2            �S@������������������������       ���҂��?+            @Q@������������������������       �z�G�z�?             $@                           �?�A��_\�?�            �@                          �@@ݝ�9+��?�           ؃@                           �?�';���?�           p�@������������������������       ��d/�ď�?�            �o@������������������������       �,���@��?�            �v@������������������������       �$�q-�?             *@                          �2@@z�����?           P|@                          �1@l(�����?b             c@������������������������       �`��NF<�?4            �T@������������������������       ��l%�|�?.            @Q@                          �4@}�W�{��?�            �r@������������������������       �C��j��?/            �P@������������������������       ����W$�?�            `m@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �f@      >@     �F@      9@      a@     p�@     �D@     ؐ@      :@      @      T@      K@     ��@     `@      8@     @n@      a@      8@      ?@      1@     �Z@     �~@      C@     x�@      7@      @     @R@      G@     �@     Pw@      7@     �i@     �`@      6@      =@      .@     �Y@     0{@      B@     ��@      5@      @      P@     �F@     �|@     �u@      5@      g@     �O@      &@      0@      "@     �K@     �h@      1@     @m@      1@       @      A@      3@     �i@      d@      *@     @Y@      (@       @      @              .@      @@      @      @@      @      �?       @       @     �J@     �H@      @      B@     �I@      "@      $@      "@      D@     �d@      ,@     @i@      *@      �?      :@      1@     @c@      \@      "@     @P@     �Q@      &@      *@      @      H@     �m@      3@     @w@      @       @      >@      :@      p@     �g@       @      U@      7@      �?      @       @      2@      V@      @     @^@       @              @      .@      X@     �B@      �?      6@     �G@      $@       @      @      >@     �b@      0@     `o@       @       @      7@      &@      d@      c@      @      O@      @       @       @       @      @     �L@       @     @\@       @              "@      �?     �I@      6@       @      3@       @       @       @              @      C@       @     �V@                      "@              <@      2@       @      0@       @       @       @              @      7@      �?     �M@                      "@              9@      ,@              0@                                              .@      �?      ?@                                      @      @       @               @                       @              3@              7@       @                      �?      7@      @              @       @                       @              3@              .@       @                      �?      5@      @              @                                                               @                                       @                              G@      @      ,@       @      =@     @h@      @     pv@      @      @      @       @      n@      `@      �?      C@     �@@      @      (@      @      2@     �Y@       @      k@      @      @      @      @     @]@      U@      �?      6@      @@      @      (@      @      2@     �Y@       @     �i@      @      @      @      @     @]@      U@      �?      6@      8@      @      @              @     �G@      �?     �Q@      @       @       @       @      D@      D@      �?      @       @              @      @      (@      L@      �?     �`@              �?       @      @     @S@      F@              .@      �?                                                      (@                                                                      *@      @       @      �?      &@     �V@      �?     �a@                      @       @     �^@     �F@              0@      @                      �?      @      9@      �?      D@                      �?      �?      K@      (@              @      @                              @      0@      �?      6@                              �?      2@      "@              @      �?                      �?              "@              2@                      �?              B@      @                      @      @       @               @     �P@             �Y@                       @      �?     @Q@     �@@              "@      @      �?      �?              @      3@              6@                       @      �?      @      @               @       @       @      �?              @     �G@              T@                                      P@      <@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ!�eyhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �<@���,%o�?�	           ��@       	                     @vW�6��?	           z�@                           �?��>����?t           f�@                            �?�a,����?�           ��@������������������������       �u���D�?2           �@������������������������       �Vq�����?�            �s@                           @����@�?�           �@������������������������       �(i�޼*�?�           ��@������������������������       �;u�}11�?�           H�@
                          �2@�~�z�J�?�           (�@                           �?϶��@�?�            q@������������������������       �4���D�?S            @]@������������������������       �f����?_            �c@                           @ZD�6�?�           ȇ@������������������������       ��Teݕ�?�            Pu@������������������������       �(0����?           @z@                            @���>�V�?�            �p@                            �?WY>��?m            �c@                           �?�`���?+            �P@������������������������       �>;n,��?             &@������������������������       �/����?$             L@                            �?ܳ�����?B            �V@������������������������       �2�{�y�?.            �M@������������������������       �     p�?             @@                          �@@PE=l18�?B            �[@                           �?(��&y��?6            �U@������������������������       �      �?	             0@������������������������       �T/e	w�?-            �Q@������������������������       �h�d0ܩ�?             7@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      <@     �I@      7@     �[@     H�@      B@     �@      7@      "@     �P@      N@     0�@     �@      &@     0p@      h@      :@      I@      7@     �Z@     ��@      B@     X�@      2@       @     �O@      K@     ��@     @@       @      o@      c@      5@     �@@      5@      V@     �{@      <@     ��@      .@      @      H@      H@     �{@     Pw@       @     �h@     @S@      ,@      :@       @     �K@      k@      1@      p@      $@      @      3@      8@     @h@     @f@      @     @Y@      K@       @      5@      @     �A@      f@      .@      i@      @      @      0@      ,@     �c@      \@      @      Q@      7@      @      @      �?      4@      D@       @      M@      @       @      @      $@      C@     �P@       @     �@@     �R@      @      @      *@     �@@     `l@      &@     �z@      @      �?      =@      8@      o@     `h@      @     �W@     �C@      @       @       @      0@     @V@             �f@      @              $@      (@      `@     �O@             �C@      B@      @      @      @      1@     @a@      &@     @o@      �?      �?      3@      (@      ^@     �`@      @      L@      D@      @      1@       @      2@     `d@       @     `v@      @      �?      .@      @     `k@     �_@              J@      (@      �?      @       @      @     �C@      �?      V@                       @      �?     �R@      7@              *@      @      �?      �?      �?      @      4@      �?      =@                       @      �?      ?@      $@               @      "@              @      �?      @      3@             �M@                                     �E@      *@              @      <@      @      (@              (@      _@      @     �p@      @      �?      @      @      b@      Z@             �C@       @              "@              @      E@      @      a@                      @      �?      N@      G@              5@      4@      @      @              @     �T@      @     �`@      @      �?              @     @U@      M@              2@      .@       @      �?              @     �E@             �[@      @      �?      @      @     �H@      *@      @      &@      @       @      �?              �?      4@             �P@      @              @      @     �A@      "@              &@      �?                                      "@              B@      �?                              *@      @               @                                              @              @                                              �?                      �?                                      @              ?@      �?                              *@      @               @       @       @      �?              �?      &@              >@       @              @      @      6@      @              "@               @      �?              �?      $@              .@       @               @      �?      ,@      @              @       @                                      �?              .@                       @       @       @                       @      (@                              @      7@             �F@       @      �?              @      ,@      @      @               @                              @      7@              ?@       @      �?              @      "@      @      @                                              �?      @              @                              @       @                               @                               @      0@              <@       @      �?                      @      @      @              @                                                      ,@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ`e8hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?�u���?�	           ��@       	                     @	�����?�           L�@                            �?�p��}C�?<           `�@                            �?Y����?�           ��@������������������������       �(���v��?           �z@������������������������       ����'_�?�            Pv@                           @�����?K            �^@������������������������       ��q�q,�?9             X@������������������������       �fw���?             ;@
                           @<f���m�?�           8�@                           �?d�i*��?�           Ȃ@������������������������       ���'���?�             n@������������������������       ����ы~�?�            �v@                          �:@�=��h��?             G@������������������������       ��paRC4�?             A@������������������������       �      �?             (@                           @a�+���?�           l�@                          �?@e�f���?x           (�@                           �?S�[���?k           ��@������������������������       ��#�f���?           �{@������������������������       �[�1���?L           ��@������������������������       ��������?             4@                            @��2��?T           D�@                            �?R����"�?�           ��@������������������������       ��UL�;��?�            @r@������������������������       �w�.��?           ��@                           @��,�s�?�             n@������������������������       �д>��C�?H             ]@������������������������       ���x[��?J            @_@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �e@      @@     �D@      <@     �Z@     Ȅ@      F@     ��@      3@      &@      W@     �H@     �@     0@      2@     �q@     �S@      ,@      3@      0@     �A@     �o@      ,@     P|@      $@      @     �E@      2@     �p@      h@       @     ``@     �F@      "@      *@      (@      7@     �b@      $@     @l@      @              @@      *@      a@     @^@      @     �Y@      E@      @      (@      (@      6@      a@       @     �j@       @              :@      *@     �[@     @Y@      �?     @T@      4@      @      @      @      (@     �T@      @     �_@      �?              ,@       @      P@      J@      �?      ;@      6@      @       @      @      $@      K@      @     @U@      �?              (@      @      G@     �H@              K@      @      @      �?              �?      ,@       @      ,@      @              @              ;@      4@      @      5@      @      @      �?              �?      *@       @      @       @              @              9@      &@      @      3@                                              �?              "@      @                               @      "@      �?       @      A@      @      @      @      (@     @Y@      @     `l@      @      @      &@      @      `@      R@      �?      =@      A@      @      @      @      (@     @X@      @     �i@      @      @      &@      @     �^@     �M@      �?      =@      8@      @      @              @      B@      �?      P@       @       @      "@      �?     �H@      9@              *@      $@      �?      �?      @      @     �N@      @     �a@      �?       @       @      @     �R@      A@      �?      0@                                              @              7@                                      @      *@                                                              @              ,@                                      @      *@                                                                              "@                                      @                              X@      2@      6@      (@      R@     �y@      >@     ��@      "@      @     �H@      ?@     p@      s@      $@      c@     �G@      @      @      @      :@     @f@      (@     `o@      �?      �?      ,@      @      p@     �b@       @      B@     �G@      @      @      @      9@      f@      (@     �m@      �?      �?      ,@      @     p@     `b@       @     �A@      9@      @      @       @      3@     �W@      &@     �T@      �?              @      �?     @W@      T@      �?      6@      6@       @      @      �?      @     @T@      �?     �c@              �?      $@      @     �d@     �P@      �?      *@                                      �?       @              *@                                      �?       @              �?     �H@      (@      .@      "@      G@     `m@      2@     �w@       @      @     �A@      9@     �n@     �c@       @     @]@     �H@       @      .@       @     �D@     �h@      1@     �q@       @      @      <@      7@     `h@     @`@       @      Z@      &@      �?               @      @     �K@      @     @X@       @               @      @      N@      ;@      @      2@      C@      @      .@      @      B@     �a@      (@      g@      @      @      :@      3@     �`@     �Y@      @     �U@              @              �?      @     �B@      �?     �W@                      @       @      I@      ;@              *@               @                      �?      2@             �J@                       @              >@      @              @               @              �?      @      3@      �?     �D@                      @       @      4@      7@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�6�FhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?�%��.��?�	           ��@       	                   �?@�3�H�h�?]           ��@                          �1@����r�?F           ,�@                            �?������?�            �t@������������������������       �Us�k���?q            �e@������������������������       ��&;����?`            @d@                            @���]<�?u           ��@������������������������       ��"��!��?f           Ў@������������������������       �%rj���?           0z@
                          �@@��Ze��?            �A@                           �?���H�?             9@������������������������       ��)x9/�?
             ,@������������������������       �                     &@������������������������       ���Q��?             $@                          �;@|T���	�?N           ��@                            @1�g�4�?�           t�@                            �?GӇc���?J           ��@������������������������       �z7�b�E�?c           h�@������������������������       ��ۊ>@t�?�            �v@                          �9@����3I�?Z           (�@������������������������       �� �)�?7           �~@������������������������       �*x9/��?#             L@                            @f�<86�?�            �o@                          �@@Z?`���?r            �d@������������������������       ��6�J�?g            �a@������������������������       �ŕ�(�?             5@                          �@@�`Y5J��?8            �V@������������������������       ��P��#�?-            �Q@������������������������       �
ףp=
�?             4@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      =@     �B@      =@     @U@     8�@      H@     ��@      4@      $@     �W@     �P@     P�@     �@      *@      s@     �Y@      0@      ;@      *@     �L@     �s@      ?@     `x@      &@      @      G@      H@     @t@     �k@      @      d@     �X@      0@      ;@      *@     �L@     ps@      ?@     w@      "@      @      G@      H@      t@     �k@      @      d@      0@      @      "@       @      *@     �K@      ,@     �G@       @              "@      *@     �K@      N@      �?     �A@      *@              @       @      @      A@      @      7@       @               @      @      <@      ?@      �?      ,@      @      @      @               @      5@      @      8@                      @      "@      ;@      =@              5@     �T@      *@      2@      &@      F@      p@      1@      t@      @      @     �B@     �A@     �p@     `d@      @     @_@     �I@      "@      *@      $@      >@     �g@      .@      h@      @      @      ;@      =@     �e@     �]@      @     �[@      ?@      @      @      �?      ,@     @P@       @      `@              �?      $@      @     �V@     �F@      �?      .@      @                                      @              5@       @                              @                              �?                                       @              1@       @                              @                              �?                                       @              @       @                              @                                                                                      &@                                                                      @                                      �?              @                                      �?                             �]@      *@      $@      0@      <@     �t@      1@     Є@      "@      @      H@      2@     `z@     �q@      @      b@     �\@      *@      $@      .@      :@     �q@      ,@     ��@      @      @     �E@      .@     �w@     �p@      @     �`@     �V@      "@       @      (@      4@     �i@      ,@     �u@      @      @     �D@      *@     �n@     �j@      @     @Z@      O@      @      �?      $@      .@     �d@      (@     �q@       @              0@      @      h@     ``@      @     �Q@      <@      @      @       @      @      D@       @     @Q@      �?      @      9@      @     �K@     @T@      �?     �A@      8@      @       @      @      @      T@             �j@       @               @       @      `@     �J@      �?      <@      8@      @       @      @      @      R@             �h@       @               @       @     �Z@     �F@      �?      9@              �?                               @              ,@                                      6@       @              @      @                      �?       @     �H@      @     �Y@      @       @      @      @      G@      3@      �?      &@      @                      �?              =@      @     �J@      @              @      @      A@      2@      �?      $@      @                      �?              4@      @     �J@      @              @      �?      ?@      *@      �?       @                                              "@                                               @      @      @               @      �?                               @      4@              I@      �?       @                      (@      �?              �?                                       @      4@             �B@      �?       @                      @      �?              �?      �?                                                      *@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��rhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @�3����?�	           ��@       	                     �?����?�           ��@                           �?:�B��?           �@                          �?@Y��Em�?�           ��@������������������������       ��I����?�           ��@������������������������       �H�7�&��?             .@                           @M%�f'��?2           <�@������������������������       �\i��W��?�           x�@������������������������       ��v:��U�?N            �@
                          �;@Ҝ�b��?�           (�@                           �?w��78�?�           ��@������������������������       �:*9�<d�?�            �s@������������������������       �ڪ�����?�            �u@                           �?<,Ԛ��?$             I@������������������������       �k��\��?             1@������������������������       ��rW���?            �@@                           �?�6���?�           ؑ@                          �0@w�����??           0�@������������������������       ��|�j��?	             .@                          �<@E�0�]��?6           p@������������������������       �l�?�\{�?           0|@������������������������       ��`��"�?!             J@                           @[5�I.�?�           ��@                          �;@�o�n�?&           �|@������������������������       ��5�S8��?           py@������������������������       ����.H;�?#            �H@                           @�3_�?b             e@������������������������       �;�\�?W            @b@������������������������       �D��2(�?             6@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@     �D@      B@      5@      ]@     ��@      ;@     ��@      3@       @     �U@      N@     0�@     H�@      6@      o@     `c@      ?@      =@      2@     �X@     �}@      7@     ��@      *@      @     @S@     �H@     �@     y@      3@     `i@     �Y@      .@      5@      .@      O@     0x@      .@     ��@       @      �?      G@      ;@     �x@     �q@      $@     ``@     �F@      �?      (@      "@      7@      `@      @     �l@       @              2@      0@     �a@     @T@      @     �J@     �F@      �?      (@      "@      7@      `@      @     @k@       @              2@      0@     �a@     @T@      @     �J@                                              �?              (@                                       @                              M@      ,@      "@      @     �C@      p@      (@     �s@      @      �?      <@      &@      p@      i@      @     �S@      D@       @      @      @      =@     �b@       @     �g@      @              2@       @     �`@     �Z@      @      J@      2@      @      @      �?      $@     �[@      $@     �^@       @      �?      $@      @     �^@     @W@      @      :@      J@      0@       @      @     �B@     �U@       @      `@      @      @      ?@      6@     �Z@      ^@      "@      R@     �I@      0@       @      @     �B@     �T@      @     @Z@      @      @      ?@      5@     @Y@     @\@      @     @Q@      4@      &@      @       @      5@     �C@      @     �H@      @      @       @      ,@     �C@      L@       @      B@      ?@      @      @      �?      0@     �E@       @      L@               @      7@      @      O@     �L@      @     �@@      �?                                      @      �?      8@                              �?      @      @      @      @      �?                                      �?               @                                      �?      @                                                              @      �?      0@                              �?      @      �?      @      @     �E@      $@      @      @      1@     �k@      @      y@      @       @      $@      &@     �m@      ^@      @      G@      :@       @      @      �?      &@     �[@       @      d@      �?      �?      @      @      W@     @P@      �?      9@      �?                                               @                               @       @      @       @              �?      9@       @      @      �?      &@     �[@              d@      �?      �?      @       @     �U@     �O@      �?      8@      0@       @      @      �?      $@     @Z@             �a@              �?      @       @      T@      L@              7@      "@                              �?      @              3@      �?                              @      @      �?      �?      1@       @      @       @      @     �[@       @      n@      @      �?      @      @     @b@     �K@       @      5@      *@      �?      @       @      @     �P@       @     �g@      @      �?       @      @      ]@     �A@              *@      &@      �?      @       @       @      N@       @     @d@      @               @      @     �[@     �@@              (@       @                               @      @              <@              �?                      @       @              �?      @      �?                       @      F@              I@       @              �?      @      >@      4@       @       @      @      �?                       @      D@             �C@                              @      >@      2@       @      @                                              @              &@       @              �?                       @               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJE��MhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @%��灜�?�	           ��@       	                    �?T�6`��?�           2�@                           @2����?           ��@                            �?��¨���?�           @�@������������������������       �;h����?�            �y@������������������������       ��s�/t �?�           ��@                          �7@����7��?=             W@������������������������       ��h�+�(�?&            �J@������������������������       ���Y� ��?            �C@
                           @�4�?�?�           ��@                          �;@���w�?s           p�@������������������������       ���yU��?,           �@������������������������       ��(y��i�?G            @[@                            �?�J��k�?k           ��@������������������������       �''Mp�F�?�             y@������������������������       �t���?r            �e@                           �?�>���?�           ��@                           �?F�����?o            �f@                          �6@I:�1�?2            �U@������������������������       �j\�A�
�?            �F@������������������������       �;j����?             E@                          �4@+�6g�?=            @W@������������������������       ��=��C�?            �F@������������������������       �      �?             H@                           @9��`�?0           ��@                           @7��EL�?e           ��@������������������������       �������?.           P|@������������������������       ����{���?7            �V@                          �;@.�%ݕ1�?�            �u@������������������������       �GW d��?�             r@������������������������       �N2t��E�?%            �M@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      @@     �F@      7@     �_@     H�@      4@     H�@      5@      (@     �U@      N@     �@     �~@      1@     pr@     �b@      9@      B@      5@     @[@     0~@      0@     ؅@      3@      @     �R@     �J@     �@     �w@      0@     �n@     @Q@      (@      <@      *@     �Q@     �l@      @     �o@      (@      @      =@      =@     �i@      c@      "@      a@     @P@      (@      :@      *@     �P@     �k@      @     �k@      (@      @      =@      <@     �h@     `a@      "@     @^@      1@      @      @      @      *@     @T@       @      Z@       @              .@      &@      P@      I@             �C@      H@       @      7@      $@     �J@     �a@      @      ]@      $@      @      ,@      1@     �`@     @V@      "@     �T@      @               @              @       @      �?      @@                              �?      $@      ,@              .@      @               @              @      @      �?      &@                              �?      @      *@              @                                               @              5@                                      @      �?              &@      T@      *@       @       @      C@     �o@      "@     �{@      @      @      G@      8@     �r@     `l@      @      [@      N@      "@      @      @      5@     �c@      @     �p@       @      @      :@      (@     @i@     �d@      @      O@     �K@      @      @      @      4@      b@      @      l@       @      @      :@      $@      g@      c@      @     �K@      @      @                      �?      *@              G@                               @      1@      (@       @      @      4@      @      @      @      1@     �W@      @      f@      @              4@      (@     @Y@     �O@       @      G@      "@      @       @      @      @     �P@      @      b@      @              $@      @     �S@      A@       @      ;@      &@              �?      �?      (@      <@      @      ?@                      $@      @      6@      =@              3@      I@      @      "@       @      1@     �d@      @     py@       @      @      (@      @     �k@      [@      �?     �I@      ,@              @               @      <@              K@                      @              @@      =@              ,@       @                                      1@              5@                      @              4@      &@              @      @                                      @              (@                      @              $@      �?              @      @                                      $@              "@                                      $@      $@                      @              @               @      &@             �@@                                      (@      2@              @      @              @              �?      �?              *@                                      @      @              @                      �?              �?      $@              4@                                      @      &@                      B@      @      @       @      .@     @a@      @     v@       @      @      "@      @     �g@     �S@      �?     �B@      <@      @      @       @      $@     @R@      @      j@               @      @      �?     @a@      F@              5@      2@      @      @       @      $@      K@      @      f@               @      @              ^@      D@              0@      $@                                      3@              ?@                       @      �?      2@      @              @       @      @      �?              @     @P@      �?      b@       @      @      @      @     �J@     �A@      �?      0@       @      @      �?              @     �G@      �?     @]@              @      @      @      G@     �A@              ,@                                      �?      2@              <@       @                              @              �?       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJq�DFhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�sw{�?�	           ��@       	                    �? �qJV��?�           ��@                          �1@W���q�?           ��@                           @]�b8��?�             q@������������������������       �(>�����?F            �Z@������������������������       �5M�4M��?Z             e@                           @00Ef;�?r           ��@������������������������       ��,��P#�?2           0@������������������������       �P��9"�?@            ~@
                            �?��5���?�           ܗ@                          �=@������?�           8�@������������������������       ��������?�            �@������������������������       �ɔLɔL�?4            �S@                          �=@�}��
�?�            �v@������������������������       ��4ؖ��?�            u@������������������������       ��������?             8@                          �=@z�����?�           ��@                          �4@��=�8��?�           (�@                           @��� ��?E           �}@������������������������       �[�b��?�            �s@������������������������       �"�	³a�?v            @d@                          �;@'�f��?Z           `�@������������������������       �O�!J[��?2           �~@������������������������       �     �?(             P@                           @��(@J�?8            @X@                           �?Fp�u=q�?             G@������������������������       �b���i��?             6@������������������������       �9��8���?             8@                           �?��S���?            �I@������������������������       ��4_�g�?             6@������������������������       �hha�H��?             =@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@      =@     �@@      6@      ^@     ��@      D@     ��@      0@      @     �S@      M@     8�@     �@      2@      p@     �c@      7@      9@      2@     @W@     �{@     �@@     h�@      (@      @     @P@      I@     @     @y@      1@      k@     @R@      &@      3@      (@      M@     `i@      0@     �q@      @      @      <@      <@      k@     �e@      @      ]@      2@      @      @      @      1@      F@      @     �B@               @      @      @     �K@      E@       @     �A@      @       @      @              @      2@      @       @                      �?              =@      2@      �?      &@      &@      �?              @      *@      :@              =@               @      @      @      :@      8@      �?      8@     �K@       @      .@      "@     �D@     �c@      *@      o@      @      @      7@      8@     @d@     @`@      @     @T@      =@      @       @      @      6@      X@      @     ``@      @      @      .@      *@      S@      G@      �?     �D@      :@      @      @       @      3@     �O@      "@     �]@      @               @      &@     �U@      U@       @      D@     @U@      (@      @      @     �A@     `n@      1@     �z@      @       @     �B@      6@     �q@      m@      (@     @Y@      M@      "@      @      @      3@     �h@      &@     �v@      @              0@      0@     �k@      e@      @      Q@      L@      "@      @      @      3@      f@      &@      v@       @              .@      .@      i@      d@      @     �N@       @                                      4@              .@      �?              �?      �?      7@       @              @      ;@      @      @      @      0@      G@      @      P@      @       @      5@      @     �L@     �O@       @     �@@      ;@      @      @      @      0@      G@       @      I@      @       @      4@      @     �L@     �O@      @      ?@                                                      @      ,@                      �?      �?                       @       @     �A@      @       @      @      ;@      g@      @     �y@      @              ,@       @     �n@      a@      �?     �D@      <@      @       @      @      2@     �e@      @     w@       @              ,@       @     @k@      a@      �?     �D@      ,@      @      @      @      (@     �Q@      @     �f@      �?              "@      @     �Y@     �G@              5@       @      �?      �?      @      @      I@             �[@      �?              @       @     @T@      ?@              *@      @      @       @              @      5@      @     �Q@                       @      @      6@      0@               @      ,@      �?      @              @     �Y@      @     �g@      �?              @      @     �\@     @V@      �?      4@      *@      �?      @              @     �U@      @     �d@      �?              @      @     @[@     �S@      �?      0@      �?               @                      1@              8@                                      @      $@              @      @                              "@      &@             �C@       @                              <@      �?                      @                              @       @              6@      �?                              "@      �?                                                      @      �?              @      �?                               @                              @                              �?      �?              .@                                      �?      �?                       @                              @      "@              1@      �?                              3@                               @                              @       @               @                                      @                                                                      @              "@      �?                              (@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ#�@hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �0@ܰ�[^��?�	           ��@       	                    @Чu�g�?�            @j@                           �?�WV��?f            �c@                            �?��	"P7�?6             S@������������������������       ����$��?             �G@������������������������       �Ĝ�-�?             =@                           @���(\O�?0             T@������������������������       �uH�����?             ?@������������������������       ���Z��?            �H@
                           @໑ɒ��?%             K@                            �?B����?             E@������������������������       ����(\��?             4@������������������������       �}��7�?             6@������������������������       ��8��8��?             (@                            @"8�X#f�?	           �@                           �?��ײ���?l           t�@                          �<@Y[���l�?�           �@������������������������       ��;1qp�?�           ��@������������������������       ���f��J�?)            �P@                           �?���0j�?�           ��@������������������������       ������?*            ~@������������������������       �"qq���?w           ��@                          �=@"�����?�           ��@                          �2@�W���?u           h�@������������������������       �=�+���?�             n@������������������������       ��g����?�           ��@                           �?)\���h�?4             T@������������������������       �������?             >@������������������������       ��e��a��?$             I@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `k@      9@     �A@      8@     �[@     ��@      @@     `�@      0@      @      T@     �O@     (�@     (�@      8@     `o@      0@                      @      @     �D@      @      =@                      @       @     �D@      B@      �?      5@      &@                      @       @      B@      @      4@                      @      @      B@      3@              .@      �?                      �?       @      1@       @      (@                       @      @      0@      2@              �?                              �?       @      ,@       @      @                              �?       @      ,@                      �?                                      @              @                       @      @       @      @              �?      $@                       @              3@       @       @                       @       @      4@      �?              ,@                                              "@              @                               @      *@      �?              @      $@                       @              $@       @      @                       @              @                      &@      @                              @      @      �?      "@                               @      @      1@      �?      @      @                                      @      �?       @                               @      @      0@      �?      �?       @                                      @              @                               @      @      @              �?       @                                       @      �?      @                                      �?      &@      �?              �?                              @                      �?                                      �?      �?              @     `i@      9@     �A@      5@     @Z@     H�@      ;@     �@      0@      @      S@     �K@     ��@     ~@      7@     �l@     �c@      1@      8@      1@     �S@     �y@      8@     ��@      *@      @     �P@     �G@     �~@     v@      7@     �h@     �R@      "@      2@       @     �E@      g@      ,@      q@      @      @      :@      8@     @g@     �c@      *@     @Z@     @R@      "@      0@       @     �C@     `f@      ,@      o@      @      @      3@      8@     �f@     �a@      *@     @Y@       @               @              @      @              7@                      @              @      1@              @     �T@       @      @      "@     �A@     �l@      $@      z@      @      �?      D@      7@      s@     `h@      $@     @W@      =@      �?       @       @      &@     @P@      �?     �b@      �?              @      ,@     �]@     �K@      �?      <@     �J@      @      @      @      8@     �d@      "@     �p@      @      �?     �B@      "@      g@     �a@      "@     @P@      G@       @      &@      @      ;@     @e@      @     �x@      @              $@       @     @n@      `@              @@      D@       @      &@      @      3@     @c@      @     �v@       @              $@       @     �k@      `@              ?@       @              @       @      @      C@             �R@                      @      �?      Q@     �@@              @      @@       @      @       @      ,@      ]@      @     Pr@       @              @      @      c@     �W@              :@      @                               @      0@              :@      �?                              6@                      �?      @                              @       @              @                                      "@                      �?      �?                               @      ,@              3@      �?                              *@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ>%8mhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @��-ƀ�?�	           ��@       	                   �?@�^n0~�?(           ަ@                          �1@�%�Y���?           X�@                            �?;�*���?9           �@������������������������       ��55��?N            �`@������������������������       ���:j��?�            �w@                          �3@&���m�?�           T�@������������������������       �g���hO�?x           @�@������������������������       ��E-\��?P           ��@
                           @ ȥ=���?'            �P@                           �?���u�?            �@@������������������������       �&���^B�?             2@������������������������       �����2�?
             .@                           @RC4%�?             A@������������������������       �P�|�@�?             1@������������������������       ��������?
             1@                            @��qn�?n           Ў@                           @ �CM���?�           ��@                          �7@vl]���?]           X�@������������������������       �G�n#0�?�            �w@������������������������       ��ϋj�0�?n             f@                          �0@�������?l             e@������������������������       ��n���?             2@������������������������       �����S��?`            �b@                           �?����?�            pp@                          �;@M:�f@�?b            �b@������������������������       �L����{�?K            @\@������������������������       �ޯ�f��?             C@                           @�Cc}h��?C             \@������������������������       �06eg�w�?,            �Q@������������������������       �q\�yQ�?            �D@�t�b��     h�h4h7K ��h9��R�(KKKK��h��B�        f@      D@     �G@      4@      \@     ��@      >@     ��@      ;@      (@     @U@     �R@     h�@     �~@      <@     �l@     �`@      ;@      C@      3@     �W@     �~@      3@     H�@      1@       @     �K@     �K@     8�@     �t@      3@     �g@     �`@      ;@      C@      3@     �W@     `~@      .@     H�@      1@       @     �K@     �K@     ��@     �t@      2@     �g@      A@      �?      @       @      1@     �Y@      @      ]@               @      $@      $@     �Z@     �K@      @      D@      $@               @              @      1@      �?     �F@                              @      ;@      0@               @      8@      �?      @       @      *@     �U@      @     �Q@               @      $@      @      T@     �C@      @      @@     �X@      :@      @@      1@     @S@     �w@      $@     ��@      1@      @     �F@     �F@     �|@     `q@      (@     �b@      :@      @      @      @      7@      S@       @     �j@              �?      ,@      "@     �]@     �M@      @      <@     @R@      7@      =@      ,@      K@     0s@       @     �}@      1@      @      ?@      B@     @u@     `k@      @      ^@       @                              �?      @      @      @@                                      2@      �?      �?      �?      �?                              �?                      5@                                       @              �?      �?      �?                                                      *@                                      @                                                              �?                       @                                      @              �?      �?      �?                                      @      @      &@                                      $@      �?                                                              @      @      @                                      �?      �?                      �?                                      �?              @                                      "@                             �D@      *@      "@      �?      1@      e@      &@     �q@      $@      @      >@      3@     �d@      d@      "@     �D@     �@@      $@      @      �?      .@     @^@       @     @h@      $@       @      :@      .@     �\@      _@      @     �B@      :@       @      @      �?       @     @X@       @     �b@      $@       @      3@      (@     �W@      V@      @      8@      7@       @      @      �?      @     �P@       @     @U@      $@              "@      $@     @R@     �L@      @      ,@      @                              @      >@              P@               @      $@       @      6@      ?@              $@      @       @       @              @      8@             �F@                      @      @      4@      B@       @      *@      �?                              �?      �?               @                                              $@              @      @       @       @              @      7@             �E@                      @      @      4@      :@       @      $@       @      @       @               @     �G@      @     @W@               @      @      @     �I@      B@      @      @      @               @              �?      4@              N@               @              �?     �@@      3@      @      @      @               @              �?      "@             �E@               @              �?      ;@      1@      @      @       @                                      &@              1@                                      @       @                       @      @                      �?      ;@      @     �@@                      @      @      2@      1@              �?       @      �?                      �?      .@      @      8@                      �?      @      &@      "@              �?               @                              (@              "@                      @              @       @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJPhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@ɺO*���?�	           ��@       	                    �?�`��@��?�           "�@                           @H��=e�?�           ��@                          �1@�)�Z�?G           ��@������������������������       ��f�� �?�            �p@������������������������       ��38�F�?�           ��@                            �?RD���v�?�            �m@������������������������       �	$N�G��?^             a@������������������������       ���A�x�?>            �X@
                           �?B"���?�           ��@                            �?iA� �?�            �q@������������������������       ��3��b�?3            �S@������������������������       �ɦj��?�            @i@                           @�mQzT�?�           T�@������������������������       �9>���?           �@������������������������       ���V�Q�?�           ��@                           �?+1�o'��?           �{@                            �?������?t             f@                           @5_�g���?             F@������������������������       ��}��?            �@@������������������������       �b���i��?             &@                           �?���¨k�?V            �`@������������������������       �,R�n��?/             R@������������������������       �AHa*�?'            �N@                           @G��3yT�?�            pp@                           @j��и<�?�             l@������������������������       �c��v��?0            �S@������������������������       ���(�?Y            `b@                           @ԍx�V�?             C@������������������������       �      �?	             (@������������������������       ��N��N��?             :@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �m@     �A@     �B@      ;@     �]@     ��@      =@     (�@      5@      &@      P@     @R@     h�@     (�@      7@     �n@     �j@      >@     �A@      :@      \@     P�@      ;@     ��@      0@      &@      L@      Q@     ��@     �}@      1@     �k@     @Z@      5@      :@      (@     �P@      q@      1@     `v@      $@       @      <@     �@@     �p@     �k@      "@     �]@      W@      2@      7@      $@      F@     �m@      .@     �r@      $@      @      9@      =@      m@      g@      "@     @X@      1@      @      "@              *@      D@      @     �D@      @      �?      @      &@     �H@     �F@      @      7@     �R@      ,@      ,@      $@      ?@     �h@      &@     `p@      @      @      5@      2@      g@     `a@      @     �R@      *@      @      @       @      6@      A@       @     �K@               @      @      @     �A@      B@              6@      (@               @      �?      *@      :@      �?      =@               @              @      4@      (@              .@      �?      @      �?      �?      "@       @      �?      :@                      @              .@      8@              @     @[@      "@      "@      ,@      G@     �q@      $@     ��@      @      @      <@     �A@     pz@     �o@       @     �Y@      0@               @      �?       @      @@      �?     �P@                       @      �?      S@      J@      @      3@      @                      �?       @      0@      �?      8@                                      2@       @              @      (@               @              @      0@             �E@                       @      �?      M@      F@      @      .@     @W@      "@      @      *@      C@     @o@      "@     �~@      @      @      :@      A@     �u@     `i@      @     �T@     �H@      @      @       @      .@     @^@      @     �p@      @      �?      &@      2@     �i@     @]@       @      @@      F@      @      @      @      7@      `@      @     @l@      �?       @      .@      0@     �a@     �U@      @     �I@      9@      @       @      �?      @     @R@       @     @f@      @               @      @      M@      E@      @      7@      3@               @              @      0@              R@       @              @       @      4@      7@       @      $@                                      @      @              7@                      �?              @       @              @                                      @      @              4@                      �?                      �?              @                                                              @                                      @      �?              @      3@               @                      &@             �H@       @              @       @      0@      5@       @      @      ,@               @                      @              9@       @              @       @      @      $@       @      �?      @                                      @              8@                                      (@      &@              @      @      @              �?      @     �L@       @     �Z@      @               @      @      C@      3@      @      *@      @      @                      @      F@       @     �W@       @               @      @      :@      3@      @      *@       @      @                      �?      0@       @      5@                      �?       @      ,@      @       @      @      @                              @      <@             �R@       @              �?      �?      (@      (@       @       @                              �?              *@              &@      �?                              (@                                                      �?              �?              @                                      @                                                                      (@              @      �?                               @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���2hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @	�4�Fb�?�	           ��@       	                   �0@�<i���?�           Х@                            �?+sI�v�?t            �f@                           �?�]�W��?S            @^@������������������������       ���O"�?!            �G@������������������������       �em��7��?2            �R@                           @��Ɉ�?!            �M@������������������������       ��8��8��?             (@������������������������       ��W+J���?            �G@
                            �?W��'A��?�           h�@                            �?ci��e�?�           �@������������������������       �0����?Q           ��@������������������������       �ٚ#	���?�           ��@                           �?��C"���?�           ��@������������������������       �xz�,C�?#             I@������������������������       �<ݚu�?s            �@                          �<@��v>��?�           ��@                           @�.��u"�?u           P�@                           �?�<�h2�?%           H�@������������������������       �m��?�            `w@������������������������       �H7Ȫ%�?3           0}@                           �?�$�N%�?P             `@������������������������       ���O"�?            �G@������������������������       ��{���?2            �T@                           �?��_���?S            �b@                           @T�r
^N�?             L@������������������������       ��|Ӭ��?            �A@������������������������       �:/����?
             5@                          �=@��$j�R�?5            �W@������������������������       �0���?             7@������������������������       �r�q��?(             R@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `h@      4@      @@      5@     @[@     ��@     �B@     �@      0@      .@     �Q@      P@     X�@     0@      3@     `p@     @b@      0@      9@      1@     @U@     �@      8@     x�@       @      &@      N@      L@     �@     �v@      2@     @l@       @      �?      @      �?      "@      @@      �?      ?@      �?      @      @      @      9@      B@      @      7@                      @      �?      @      3@      �?      9@      �?               @      �?      2@      ;@              2@                       @      �?       @      (@      �?      @      �?               @              @      ,@              @                      �?              @      @              4@                              �?      ,@      *@              .@       @      �?                      @      *@              @              @      �?      @      @      "@      @      @                                      @      @                                              @                               @       @      �?                      �?      $@              @              @      �?              @      "@      @      @      b@      .@      6@      0@      S@     �}@      7@     ��@      @      @     �L@     �I@     @~@     pt@      .@     `i@     �X@      .@      &@      *@     �I@     �w@      1@     p�@      @       @      E@      @@      x@     �k@      *@     `a@     �J@      @      @      @      5@     �d@      @     �q@      �?              2@      (@      g@      ]@      @     �G@      G@      $@       @      @      >@      k@      $@     @q@      @       @      8@      4@      i@     @Z@       @      W@     �F@              &@      @      9@     �W@      @     @`@       @      @      .@      3@     �X@     �Z@       @      P@      @              @      �?              @              @      �?              �?              $@      @              (@      E@              @       @      9@     @V@      @     �_@      �?      @      ,@      3@      V@     �X@       @      J@     �H@      @      @      @      8@     �f@      *@     �z@       @      @      $@       @     �i@      a@      �?      B@     �E@      @      @      @      3@     �c@      *@     �u@      @      @      $@      @      g@      `@      �?      A@     �B@      @      @      @      1@      _@      $@     0s@      @      @      "@      @      e@     @\@      �?      =@      7@      @      @              &@     @P@      @     �\@      �?      @      @       @     �R@      H@              .@      ,@                      @      @     �M@      @      h@      @              @      @     �W@     @P@      �?      ,@      @      �?      �?      �?       @      A@      @     �E@                      �?      �?      0@      .@              @      @                              �?      (@              &@                      �?      �?       @      @              �?              �?      �?      �?      �?      6@      @      @@                                       @      "@              @      @                              @      8@             �S@      @      �?              �?      5@       @               @      @                                      @              A@       @                      �?      @      @              �?      @                                       @              1@       @                      �?      @      @              �?       @                                       @              1@                                                                      �?                              @      4@             �F@       @      �?                      0@      @              �?                                               @              $@                                              @              �?      �?                              @      (@             �A@       @      �?                      0@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJi�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@�[���?�	           ��@       	                    �?�^����?�           �@                           �?ŗ��,�?�           |�@                            @)xI:�?�             j@������������������������       �S���?O             _@������������������������       �nт4��?3            @U@                           @�])��G�?X           8�@������������������������       ���y��;�?�           @�@������������������������       ������?�            �s@
                           @b��7�?�           \�@                           �?�؉����?            �@������������������������       ������?T           ��@������������������������       ��:�N�?�            �r@                          �6@�ⲣga�?�           \�@������������������������       ����[�?�           (�@������������������������       ��#ʌ�?�             s@                           �?A����?           0}@                          �?@[14�T��?t            �g@                          �=@�� ����?V            �a@������������������������       ���-1�#�?=            �Y@������������������������       ����Դ�?             C@                          @@@4�\9���?            �H@������������������������       �dT!)��?             3@������������������������       �(}�'}��?             >@                           �?�k��X��?�            Pq@                          �>@��n���?              I@������������������������       �     ��?             @@������������������������       �0�����?             2@                            �?�;X��w�?�            `l@������������������������       ��
�'��?+            @P@������������������������       �V"�R<�?`            @d@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        j@      B@      G@      7@      X@     �@      <@     T�@      0@      @     �V@      M@     І@     ��@      .@     q@     �f@      @@     �F@      7@     �T@     ؁@      :@     ��@      $@      @      T@      K@     ��@     �~@      .@     `o@      U@      2@      >@      (@     �J@     �r@      .@     �v@      "@      @      B@      8@     pq@     �i@       @     �_@      $@      @      @              @     �B@             �P@      @              @              D@      2@              .@       @      @      @              @      4@              ?@      @              @              ;@      @              &@       @                              �?      1@             �A@                       @              *@      &@              @     �R@      .@      ;@      (@      G@     �p@      .@     `r@      @      @      >@      8@     �m@     �g@       @     �[@      N@      (@      5@      (@     �E@     �j@      @      j@       @      @      7@      .@     �h@      a@      @     �T@      ,@      @      @              @      J@      "@     @U@      @       @      @      "@      D@     �I@      @      =@     �X@      ,@      .@      &@      >@     �p@      &@     x�@      �?       @      F@      >@     �w@     �q@      @     @_@     �I@      @      @      @      &@     �\@             �o@      �?              *@      &@     �h@      Y@       @     @P@      B@              @      @      @     �R@             �b@      �?              @      "@      `@     �R@      �?     �D@      .@      @      @              @      D@             �Y@                      @       @     @Q@      :@      �?      8@      H@      &@      "@      @      3@     `c@      &@     0s@               @      ?@      3@     �f@      g@      @      N@     �C@      @      @      @      (@     @]@       @     �j@              �?      4@      "@      [@      b@      @      H@      "@      @      @      �?      @      C@      @     @W@              �?      &@      $@      R@     �C@      �?      (@      :@      @      �?              *@     �Q@       @     �g@      @              $@      @     @R@     �F@              6@      2@      @      �?              $@      6@             �P@      �?              @              ?@      5@              (@      ,@      @      �?              $@      0@             �D@                      @              =@      .@               @      @      @      �?              @      0@              ?@                      @              7@       @              @      @                              @                      $@                                      @      @              �?      @                                      @              :@      �?                               @      @              @      �?                                      �?              ,@      �?                               @                              @                                      @              (@                                              @              @       @      �?                      @     �H@       @     �^@      @              @      @      E@      8@              $@      @      �?                       @      @              *@                               @      $@       @              @      @      �?                              @               @                               @      "@      @                      �?                               @       @              @                                      �?      @              @      @                              �?     �E@       @     �[@      @              @       @      @@      0@              @       @                                      @              @@      �?               @              *@      "@              �?       @                              �?      C@       @     �S@      @              @       @      3@      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJXU<DhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@��C�c�?�	           ��@       	                    @m��w�?�           8�@                           �?����1_�?^           :�@                           �?��I�?�           ��@������������������������       ������?�            �n@������������������������       �
�����?           @�@                          �3@�����?�           ��@������������������������       ����5��?u           ��@������������������������       �%��||�?0           x�@
                          �3@�������?#           ��@                            @׷����?             y@������������������������       ��jo��?�            Pv@������������������������       �����l�?             �F@                          �7@����pn�?#           �~@������������������������       �L���?�            �t@������������������������       �(���?^            �d@                           @x1���X�?           �z@                           �?tt�J"�?�            �v@                           �?o,x���?`            �c@������������������������       ��v�[o�?2            @T@������������������������       ���L���?.            �R@                           @��]�<�?�            @j@������������������������       �U@$���?=            �W@������������������������       �-�n#�?Q            �\@                           �?vY5I�?!            �O@������������������������       ���!pc�?             &@                           �?~e�.y0�?             J@������������������������       ��q�q�?             8@������������������������       ��S�r
^�?             <@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @j@      A@      B@      5@     @X@     (�@      :@     ��@      0@      *@     �P@      O@     �@     �~@      3@     @o@     �f@      <@     �@@      4@     �V@      �@      8@      �@      *@      &@      L@     �M@     ȅ@     �|@      1@     �k@     ``@      4@      8@      .@     �J@     �}@      5@     ��@      "@       @      E@      C@     (�@     �u@      (@     �b@     �K@      .@      ,@      $@     �@@     �l@      *@     �m@      "@      @      $@      7@     @h@     �b@      @      T@      "@       @      @      @      (@     �A@      �?     �R@      @              @      @     �E@      7@              7@      G@      *@      &@      @      5@     �h@      (@     @d@      @      @      @      1@     �b@     �_@      @     �L@      S@      @      $@      @      4@     `n@       @     �|@               @      @@      .@     0v@     �h@      @     @Q@     �D@              @      @      @      X@      @     �d@                      .@      @     @f@     @S@      @      9@     �A@      @      @       @      ,@     `b@      @     Pr@               @      1@      $@      f@     @^@      �?      F@     �I@       @      "@      @     �B@     @a@      @     �p@      @      @      ,@      5@     �b@     @[@      @      R@      >@              @      @      0@     �O@       @     �_@      �?      @      $@      @     �E@      K@       @     �B@      ;@              @      @      0@     �I@       @     �Y@      �?      @      $@      @     �D@      J@       @     �A@      @                      �?              (@              7@                                       @       @               @      5@       @      @              5@     �R@      �?     �a@      @              @      .@     @Z@     �K@      @     �A@      .@      @      @              3@      K@      �?     �T@      �?              @      (@     �O@     �A@      @      =@      @      @      �?               @      5@             �M@       @                      @      E@      4@              @      <@      @      @      �?      @     @P@       @      d@      @       @      &@      @     �R@     �@@       @      =@      <@      @      @      �?      @      O@       @     @^@      @       @      $@       @     �L@     �@@       @      ;@      3@      @      @              @      .@             �G@                      @              6@      7@              ,@      (@      @       @              @      @              ;@                      @              @       @              "@      @              �?                      &@              4@                                      0@      .@              @      "@      @              �?      @     �G@       @     �R@      @       @      @       @     �A@      $@       @      *@       @      @              �?      @      3@       @      8@               @      �?       @      2@      @      �?       @      �?                              �?      <@              I@      @               @              1@      @      �?      @                                              @             �C@                      �?      �?      1@                       @                                                              @                                      @                       @                                              @              A@                      �?      �?      *@                                                                       @              (@                      �?      �?       @                                                                      �?              6@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJmn!hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @������?�	           ��@       	                    @V*�]��?           `�@                           @�/���?B           ��@                           �?]�ƭ�?           �@������������������������       �# ����?L           ��@������������������������       �E����?�           |�@                          �:@R1t4]2�?'            �Q@������������������������       �RM�ı��?!             M@������������������������       �r�q��?             (@
                          @@@d������?�           ؆@                           !@O�L ���?�           p�@������������������������       �@"���?�           ��@������������������������       ��)O�?             2@������������������������       �&�q-�?             *@                           �?�=d���?�           d�@                           @V��;e��?           `{@                          �3@����$�?�            Pu@������������������������       ��� �?M            @]@������������������������       �$I�$IR�?�             l@                          �4@wv~ثT�?:            @X@������������������������       ����|��?            �H@������������������������       �r�qG�?             H@                           �?����H2�?�           �@                          �6@����i�?9             U@������������������������       �p��$a��?#            �I@������������������������       �ogH���?            �@@                           �?R�o�?U           x�@������������������������       �W-��d�?�            @t@������������������������       �*4�+��?�            `i@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        l@      <@      D@      7@      Y@     �@      ?@     X�@      4@      @     �Q@      O@     ��@     �@      <@     �p@      f@      4@      A@      6@      T@     �|@      :@     ��@      4@      @      P@      L@     @�@     @y@      <@     �l@     �a@      ,@      :@      5@     �P@     @v@      ,@     (�@      *@      @     �F@      D@     �x@     �o@      3@     �e@     �a@      ,@      :@      4@     @P@     pu@      ,@     (�@      *@      @     �F@     �B@     Px@      o@      3@     �d@      P@      @      3@      .@      E@     `d@      @      k@       @       @      8@      4@     �b@     �[@      (@     �U@     �S@       @      @      @      7@     �f@      "@     �r@      @      @      5@      1@     �m@     @a@      @     �S@                              �?       @      *@              @@                              @      @      @              $@                              �?              *@              7@                               @      @      @              $@                                       @                      "@                              �?                                      A@      @       @      �?      *@     �Y@      (@     `e@      @      �?      3@      0@     �_@     �b@      "@      K@      @@      @       @      �?      *@     �Y@      (@     `e@      @      �?      3@      ,@     �_@     �a@      "@      K@      ?@      @       @      �?      (@     �W@      $@     `e@      @      �?      3@      ,@     �^@     �a@      "@      K@      �?                              �?       @       @                                              @      @                       @                                      �?                                               @               @                      H@       @      @      �?      4@     �f@      @     `x@                      @      @     `m@     @Z@              B@      <@      @      @              ,@     @U@      @      `@                      @       @     �U@      L@              6@      6@      @      @              &@     @Q@       @     �V@                      @       @     @S@      C@              4@      @      @                       @      0@              E@                       @      �?      9@      1@              @      2@      �?      @              "@     �J@       @      H@                      �?      �?      J@      5@              .@      @       @                      @      0@      �?     �C@                                      $@      2@               @      @       @                      @      @      �?      8@                                      @      @              �?       @                                      "@              .@                                      @      ,@              �?      4@       @      @      �?      @     �X@       @     Pp@                      @      @     �b@     �H@              ,@      @              @               @       @      �?      C@                                      1@      @              @      @              @              �?      @      �?      2@                                      "@      @              @                                      �?       @              4@                                       @       @                      *@       @              �?      @     �V@      �?     �k@                      @      @     ``@      F@              &@       @      �?              �?      @     �L@      �?      a@                       @       @      R@      =@              $@      @      �?                             �@@             �U@                      �?       @     �M@      .@              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��/3hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �0@�}�|Q��?|	           ��@                            @���3Q�?|            �i@                           @�?����?e            �d@                            �?}�/*B�?[            `b@������������������������       ��.+K�j�?            �H@������������������������       �;����t�?=            �X@������������������������       ���Q��?
             4@       	                    �?�^v�]�?            �B@������������������������       ���� =�?
             1@
                           �?ffffff�?             4@������������������������       �r�q��?             (@������������������������       �      �?              @                            @�Q�/1u�? 	           ��@                           @������?X           B�@                          �>@*��k��?}           �@������������������������       ���9~��?P           ��@������������������������       ��`����?-            @S@                            �?D����?�           8�@������������������������       ��ev���?�            �i@������������������������       �&�2�7r�?Z           Ѐ@                           �?�Ԟ�&�?�           p�@                          �1@�V�1��?,           �@������������������������       �Nj�
9��?            �H@������������������������       ����-%��?           �|@                           �?�����?|           ��@������������������������       �v�{�+�?6            �V@������������������������       ��{�҉�?F            �@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @j@     �B@      E@      D@     �Z@     (�@      B@     t�@      2@      @     �Q@     �P@     ��@     P@      4@     `n@      *@      �?       @      @      @     �E@       @      >@      �?      @      @      @     �D@     �A@              &@      &@      �?       @      @      @      C@              2@      �?      @       @      @     �C@      =@              @      &@      �?       @      @      @      9@              0@      �?      @       @      @     �B@      :@              @      �?                      @       @      @              "@                                      4@      @              @      $@      �?       @       @      @      2@              @      �?      @       @      @      1@      7@              @                                              *@               @                                       @      @                       @                                      @       @      (@                       @       @       @      @              @       @                                      �?       @                               @       @      �?      @              @                                              @              (@                                      �?      @                                                                              "@                                      �?       @                                                              @              @                                              �?                     �h@      B@      D@     �A@     @Y@     Ѓ@      A@     ��@      1@       @     �P@     �M@     P�@      }@      4@      m@      b@      :@      ?@      <@      T@     P|@      9@     (�@      *@       @      M@     �H@     }@      u@      3@      g@     �W@      7@      3@      4@     �H@     �t@      5@     ~@      &@      �?     �E@      ?@     `t@      q@      &@     �]@     @W@      7@      3@      4@      H@     �s@      1@     `|@      &@      �?      D@      =@     t@     `p@      $@     �Z@      �?                              �?      (@      @      ;@                      @       @      @      $@      �?      &@     �I@      @      (@       @      ?@     �^@      @     �h@       @      �?      .@      2@     `a@     �P@       @     �P@       @       @              @      @      ?@      �?     �S@      �?              �?       @      C@      .@      @      $@     �E@      �?      (@      �?      9@      W@      @     @]@      �?      �?      ,@      0@     @Y@     �I@      @      L@      J@      $@      "@      @      5@     �f@      "@     �y@      @              "@      $@      k@      `@      �?      H@      :@      @      @       @      (@     @X@      @     �c@      �?              "@      @     �V@     �N@              ?@      �?      �?                       @      0@              &@                              �?      @      @              @      9@      @      @       @      $@     @T@      @     `b@      �?              "@      @     �U@     �K@              8@      :@      @      @      @      "@      U@       @     �o@      @                      @     �_@     �P@      �?      1@      @              @              @      @      �?     �E@                                      (@      ,@              @      7@      @      �?      @      @     �S@      �?      j@      @                      @     �\@     �J@      �?      (@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��!hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@8A�?xi�?�	           ��@       	                   �:@(�UT��?�           �@                           �?e�!e��?5           �@                           �?v��#��?�           �@������������������������       �$C����?"           �{@������������������������       ���j���?�           4�@                           @��6��?�           ��@������������������������       �&#�X��?           `�@������������������������       �Hd:�?           ��@
                           @�v)'���?O            �`@                            �?P&�to@�?>            @Z@������������������������       �� ��t��?"            �L@������������������������       ��8��8��?             H@                            �?�Cc}h��?             <@������������������������       ���ˠ�?	             &@������������������������       ���U�(�?             1@                           @�C�p��?           0}@                           �?��;�OF�?�             w@                           �?���y�?,            �S@������������������������       ���8��8�?             8@������������������������       �b���i��?            �K@                           @?�����?�            0r@������������������������       ���Ģ���?B            �Z@������������������������       �ܳ�����?r             g@                            �?X������?3            @X@                           �?H�z�G�?             N@������������������������       ��]^m>��?             7@������������������������       �e��3��?            �B@                          �=@*7��?            �B@������������������������       �r�q��?             8@������������������������       ��(ݾ�z�?             *@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@      =@     �C@      8@     @W@     ��@      ?@     T�@      5@      $@     @P@      M@     X�@     ȁ@      1@      n@     �e@      9@      C@      5@     �U@     ��@      ?@     �@      1@      "@      L@      J@     ��@     @�@      ,@     �k@     @e@      3@     �B@      2@     @T@     ��@      <@     ��@      1@      "@      L@     �I@     H�@     �@      ,@     �k@     �R@      &@      4@      $@      K@     �p@      .@     pu@      (@      @      <@      =@     �p@     �k@      @      \@      6@              "@       @      0@     �R@       @     �\@       @       @      &@      @     �N@     �N@              K@      J@      &@      &@       @      C@     `h@      *@     �l@      @      @      1@      8@     `i@     @d@      @      M@      X@       @      1@       @      ;@     �r@      *@     8�@      @       @      <@      6@     v@     �q@      @     @[@      H@      @      ,@      @      &@      \@      @     Pp@                      @       @     �f@      [@      �?      I@      H@      @      @      @      0@     �g@      $@      r@      @       @      7@      ,@     �e@     @f@      @     �M@      @      @      �?      @      @      9@      @      ?@                              �?      D@      &@               @      @       @      �?      @      @      .@       @      6@                              �?      C@      $@              �?      @                      @       @      @       @      $@                              �?      <@      @              �?      �?       @      �?              @      (@              (@                                      $@      @                              @                              $@      �?      "@                                       @      �?              �?                                                      �?      @                                       @      �?              �?              @                              $@              @                                                                      2@      @      �?      @      @     �Q@              g@      @      �?      "@      @     �V@     �H@      @      2@      *@      @      �?              @      L@             �c@       @      �?      "@      @      N@     �B@      @      0@      @      �?                              3@              :@                      @       @      @      &@              @       @      �?                               @              @                      @       @      @       @              �?      @                                      1@              6@                                      �?      "@               @      @      @      �?              @     �B@             @`@       @      �?      @      @     �J@      :@      @      *@              �?      �?              @      "@             �D@       @      �?      �?       @      :@      $@      �?      @      @       @                       @      <@             @V@                      @       @      ;@      0@       @      @      @                      @              .@              <@       @                              >@      (@               @      @                      @              ,@              $@      �?                              3@       @                      @                                      @              @                                      @       @                                              @              &@              @      �?                              0@                                                                      �?              2@      �?                              &@      @               @                                                              *@                                       @      �?               @                                              �?              @      �?                              @      @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ&��hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @v�܋6��?	           ��@       	                     �?����?�           ��@                           @�F�ا�?           N�@                           �?�VpMc��?H           Ȍ@������������������������       �+��<F�?           �{@������������������������       ��6����?*           �}@                           @������?�           8�@������������������������       ���c�
}�?�           ��@������������������������       ��o^M<+�?            �F@
                           �?j�@����?�           ��@                           @�6��a��?�            pv@������������������������       �_([3��?�            �t@������������������������       �      �?             <@                           @p3)���?�            �v@������������������������       �;������?�            �q@������������������������       ��߿�|��?4            �U@                           @�]�4���?�           0�@                           �?ʄ^�}�??           �@                           �?�ܭei��?�            `o@������������������������       ��(�B'�?            �@@������������������������       �glq���?�            @k@                           @�l�c�Z�?�            �o@������������������������       �b��~��?�            �k@������������������������       �`)P�W
�?            �@@                           @r;�v�?l           ��@                          �:@)O��?b            �@������������������������       ����U`�?           �|@������������������������       �����W�?F            @]@������������������������       ��)O�?
             2@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        k@     �A@     �B@      B@     �W@     h�@      @@     <�@      3@      "@     @X@     �P@     `�@     0�@      &@     �m@     �d@      5@      >@      =@     �T@     �{@      ;@     @�@      2@       @     �S@     �M@      @     �z@      &@      i@     �\@      &@      5@      <@      D@      v@      7@     ��@       @      �?      E@     �C@      x@     @s@       @     �a@      M@       @      (@      0@      4@     �d@      "@     �m@       @              7@      1@     �h@     �Y@      @      L@      @@       @      &@      "@      0@     @U@      @      X@      �?              .@      $@      W@      F@       @      =@      :@              �?      @      @     @T@      @     �a@      �?               @      @      Z@      M@      �?      ;@     �L@      "@      "@      (@      4@     @g@      ,@     �t@      @      �?      3@      6@     �g@     �i@      @      U@      L@      @      "@      (@      4@     `f@      (@      t@      @      �?      3@      6@     �f@      h@      @     �S@      �?      @                              @       @      @                                      @      ,@              @     �I@      $@      "@      �?      E@     �V@      @      b@      $@      @     �B@      4@      \@     �^@      @     �N@      5@      @      @              ;@      F@       @      S@      @      @      $@      $@     �M@     �M@      �?      :@      5@      @      @              ;@     �E@       @     �N@      @      @      $@      $@      M@     �I@      �?      9@                      �?                      �?              .@      �?                              �?       @              �?      >@      @      @      �?      .@     �G@       @     @Q@      @      @      ;@      $@     �J@      P@       @     �A@      ;@      @      @      �?      $@     �C@       @     �M@               @      3@      @     �G@      B@      �?      9@      @                              @       @              $@      @      �?       @      @      @      <@      �?      $@      I@      ,@      @      @      (@     @f@      @     px@      �?      �?      2@       @     �o@     �]@             �B@      5@      @      @      @      @     �O@             �f@              �?      $@      @     �a@      I@              2@      ,@      @      @      �?      @     �D@             @P@                      @      �?     @Q@      ?@              *@      �?              �?                      &@              @                                      @      @              @      *@      @       @      �?      @      >@              M@                      @      �?     �O@      <@              "@      @              �?       @      @      6@              ]@              �?      @      @      R@      3@              @      @              �?       @      @      5@             �X@              �?      @              P@      2@              @      �?                                      �?              2@                              @       @      �?                      =@      &@      @      @      @     �\@      @     @j@      �?               @      @     �[@     @Q@              3@      =@      &@      @      @      @     �[@      @     �i@      �?               @      @     �[@      O@              1@      6@      @      @      @      @     @S@      @     @c@      �?               @      @     �X@     �L@              0@      @      @                      �?     �@@             �J@                                      &@      @              �?                                              @              @                                      �?      @               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJU�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@���_�}�?�	           ��@       	                   �0@�jK����?k           �@                            @ғj,v��?�             k@                           �?�n�tv�?r            �f@������������������������       ��z�<p�?>             Z@������������������������       �У1���?4             S@                           �?�^v�]�?            �B@������������������������       �����X�?             5@������������������������       �     ��?             0@
                           �?_1ϱ��?�           V�@                          �8@�����?�           ܖ@������������������������       ���k��!�?	           ��@������������������������       ���-�W��?|            �i@                            @�
�e��?]           Л@������������������������       �"b�����?!           ��@������������������������       �'�`d�?<           ��@                           �?�Cs��?           P|@                           @&y=d�Z�?q            �e@                            @�g\��?G             Z@������������������������       �     8�?-             P@������������������������       �ףp=
��?             D@                           @��M���?*             Q@������������������������       ��8��8��?             8@������������������������       �fP*L��?             F@                            @�~�[��?�            �q@                           @(H� ʱ�?v            `h@������������������������       ������*�?I            @^@������������������������       ��a��^�?-            �R@                           �?n:*G��?7            �U@������������������������       �ڍ�Ç�?$             M@������������������������       �4և����?             <@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        g@      ;@      B@      =@     �\@     ��@      9@     h�@      6@      @     �U@      O@     (�@     X�@      1@     �p@     `d@      8@      A@      :@     �Z@     @�@      8@     P�@      3@      @      S@     �M@     ��@     �~@      .@     `m@      "@       @              @       @      A@      @      >@      �?              @       @     �F@      F@      @      .@      @       @              @      @     �@@      @      5@      �?              @      @     �C@      A@      @      *@       @       @              @      @      5@      @      ,@      �?              �?       @      7@      0@      @      @      @                      @              (@              @                      @      @      0@      2@              @      @                               @      �?      �?      "@                       @      �?      @      $@               @      @                               @              �?                               @      �?      @      @               @                                              �?              "@                                      @      @                     @c@      6@      A@      3@     �X@     0�@      4@     `�@      2@      @     @Q@     �I@     X�@     �{@      (@     �k@     �Q@      ,@      4@      @     �J@     pq@      &@     @u@      *@       @      @@      2@     �p@      j@      @     @^@     �P@      ,@      3@      @     �I@     �k@      "@     �r@      (@       @      >@      2@      m@     `e@      @     @Y@      @              �?       @       @     �M@       @      E@      �?               @             �A@     �B@              4@      U@       @      ,@      (@      G@     �p@      "@     ��@      @      �?     �B@     �@@     �u@     �m@      @     �X@     �P@      @      @      "@     �E@     `h@       @     0v@      @      �?      A@      9@     `m@      f@      @     @U@      1@      @      @      @      @      S@      �?     �j@       @              @       @      ]@     �N@              ,@      5@      @       @      @       @     �S@      �?      f@      @      �?      &@      @     @S@      A@       @      =@      *@      �?       @              @      9@              L@      �?              @      �?      9@      4@       @      *@      @      �?       @              @      5@             �A@      �?              @      �?      (@      $@       @       @              �?       @              �?      3@              3@                      @              @       @               @      @                              @       @              0@      �?                      �?      @       @       @              @                               @      @              5@                                      *@      $@              &@                                               @              @                                      @      �?              $@      @                               @       @              ,@                                      "@      "@              �?       @       @              @      �?      K@      �?      ^@       @      �?      @       @      J@      ,@              0@      @       @              @      �?      D@      �?     �R@                      @       @      A@      $@              0@      @       @              @              <@      �?      A@                      @       @      3@      @              0@                                      �?      (@              D@                       @              .@      @                      �?                                      ,@              G@       @      �?                      2@      @                      �?                                      (@             �A@              �?                      @      @                                                               @              &@       @                              (@      �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJt��uhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�>A���?�	           ��@       	                    �?�^?�-/�?X           <�@                            �?���a$��?�           p�@                           �? ��lG�?s            �g@������������������������       ��2^���?8            �V@������������������������       �� m>�?;            �X@                            @��u���?            {@������������������������       ���aP{��?p            �d@������������������������       ������?�            �p@
                           @�BU�n>�?�           ��@                            @���	R@�?�           l�@������������������������       �ؐ�y�l�?           @�@������������������������       �JD<7j�?�            `j@                           @�7F0���?1            �Q@������������������������       ��
GJ>�?*            �M@������������������������       �*L�9��?             &@                            @ֽ���?O           ��@                            �?�SR���?�           t�@                          �>@�Rs���?�           ؒ@������������������������       �U�I���?�           <�@������������������������       ��T���6�?            �C@                          �0@hp�f��?�            pv@������������������������       ��q�q�?             8@������������������������       ������?�            �t@                           @��>�ʁ�?}           �@                           @*)����?�            @x@������������������������       ��c�[Ư�?�            @q@������������������������       ������?F             \@                          �;@�y]6���?�             k@������������������������       �{������?y            `g@������������������������       �&�X�%�?             >@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@     �H@     �B@      9@     @_@     ��@      =@     ��@      2@      (@     �S@     �P@      �@     (�@      3@     �m@     �Y@      <@      ;@      *@      R@     Pt@      0@     y@      $@      @      D@      =@     �s@     @n@      (@     @Y@     �A@      *@      2@      �?      9@      Z@      @      e@      �?       @      ,@      @     �X@      W@      �?     �B@      "@       @      @      �?      @      9@      @      P@                      @      @      ?@      5@      �?      $@      @       @                      �?      @       @      @@                      @      @      .@      (@              @      @              @      �?      @      2@      @      @@                       @       @      0@      "@      �?      @      :@      &@      .@              3@     �S@              Z@      �?       @      @       @      Q@     �Q@              ;@      @      @      (@              &@     �@@              ;@      �?              @              6@      6@              4@      4@      @      @               @      G@             @S@               @      �?       @      G@     �H@              @     �P@      .@      "@      (@     �G@     �k@      &@      m@      "@      @      :@      6@     �k@     �b@      &@      P@     �P@      .@       @      (@      E@     @j@      "@     �j@      "@      @      :@      6@     �j@     �`@      &@     �L@     �O@      "@      @      &@      C@     �e@      @      c@      "@      @      5@      4@     �d@     �Z@      &@      E@      @      @      �?      �?      @     �B@      @     �N@                      @       @      G@      :@              .@                      �?              @      &@       @      4@                                      @      1@              @                      �?              @       @              4@                                      @      *@              @                                      �?      @       @                                                      @              �?      Z@      5@      $@      (@     �J@     �u@      *@     `�@       @      @      C@     �B@     Pz@     0q@      @     �`@     �T@      .@       @       @      F@      o@      $@     `|@      @      @      B@      ?@     �q@     �j@      @     �[@      M@      $@       @       @      8@     �h@      $@     x@      @              8@      5@      m@     @e@      @      L@      M@      $@       @       @      8@      h@       @     �w@      @              8@      2@     �k@     @d@      @      J@                                              @       @      @                              @      &@       @              @      9@      @      @              4@     �I@             @Q@      @      @      (@      $@     �J@      F@      @      K@      @                                       @              �?                               @              $@                      6@      @      @              4@     �E@              Q@      @      @      (@       @     �J@      A@      @      K@      5@      @       @      @      "@     �X@      @     �l@      �?       @       @      @     �`@     �N@              9@      $@      @      �?      @      @     �F@              c@               @      �?      @     @Z@      C@              2@      @              �?      @      @      =@             �Z@               @      �?      �?     �T@      :@              0@      @      @              �?      �?      0@              G@                               @      7@      (@               @      &@      @      �?              @     �J@      @     �S@      �?              �?      @      >@      7@              @      &@      @      �?              @     �E@      @     �M@                      �?      @      >@      7@              @                                              $@              3@      �?                                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJZ�BhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @'G`bn��?�	           ��@       	                     �?���7(�?�           &�@                          �1@�U�h���?K           �@                           �?��Gd���?�            @w@������������������������       �h�)�?q            @h@������������������������       �l��A�,�?w            @f@                            �?��U��?c           �@������������������������       ��);b�"�?#           X�@������������������������       ��p�E7�?@           ��@
                           @ H�Y���?�           �@                           @⽟8���?}           ��@������������������������       �*������?�            �u@������������������������       �G���?�             p@                           @L�a��?#            �O@������������������������       �r�q��?             8@������������������������       ��o��o��?            �C@                           �?W�'�~��?�           ؐ@                           @�\ ��?|            �h@                           �?�}�BU�?r            �f@������������������������       �F���j��?8            �W@������������������������       �mweȫ�?:            �U@������������������������       �     ��?
             0@                          �2@��c�D�?;           ��@                          �1@&�7Ë��?�             h@������������������������       ���#ʆA�?F            �Z@������������������������       �bΊx��?:            �U@                           �?��a �?�           x�@������������������������       ���Dl�|�?�             r@������������������������       �B
f
ε�?�            �x@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@     �A@     �D@      4@     @Y@     �@      <@     �@      1@      &@     @U@     �S@     ؇@      �@      4@     �q@      f@      7@      >@      3@     @T@     �{@      6@     `�@      *@      @     �S@     @P@     ��@     �x@      4@     `n@      `@      0@      1@      0@      N@     �w@      ,@     @�@      $@              J@      E@     @z@     �q@      $@     �d@      8@              @      �?      *@     @Q@      @     �S@                      @      @      P@     �R@       @      <@      "@              @      �?      *@      @@      @     �@@                              @      ?@      F@       @      4@      .@                                     �B@      �?     �F@                      @      @     �@@      ?@               @     @Z@      0@      ,@      .@     �G@     `s@      $@     �}@      $@             �G@      B@     @v@      j@       @     @a@     �F@       @      @      @      .@     �b@      @     �n@      @              .@      (@     �h@     �\@       @     �F@      N@       @      $@      (@      @@     �c@      @     `l@      @              @@      8@      d@     @W@             @W@      H@      @      *@      @      5@      P@       @     �`@      @      @      ;@      7@     �\@     @\@      $@     @S@     �F@      @      $@      @      5@     �K@       @     �[@      @      @      3@      7@     �[@      Y@      $@     �R@      5@      @      @      @      &@     �D@      @     �P@      @      @      "@      @      I@     @P@      "@     �E@      8@       @      @              $@      ,@       @      F@               @      $@      0@     �N@     �A@      �?      ?@      @              @                      "@              5@                       @              @      *@              @      @              �?                       @              @                      �?               @      @              �?                       @                      �?              1@                      @              �?      "@               @      C@      (@      &@      �?      4@     �d@      @     �y@      @      @      @      *@     �l@      ]@             �D@      2@              @              $@      A@      �?     �O@                                      ?@      9@              *@      2@              @              "@      =@      �?      K@                                      >@      9@              *@       @              �?              @      0@              7@                                      4@      ,@              "@      $@               @              @      *@      �?      ?@                                      $@      &@              @                                      �?      @              "@                                      �?                              4@      (@       @      �?      $@     �`@      @     �u@      @      @      @      *@     �h@     �V@              <@      @      �?       @      �?      @      =@      �?      N@                      �?       @     �N@      4@              @      @      �?      �?               @      4@      �?     �A@                      �?       @      8@      &@              @      �?              �?      �?      �?      "@              9@                                     �B@      "@              @      ,@      &@      @              @     �Y@      @     �q@      @      @      @      &@      a@     �Q@              6@      $@      @      @              @      F@       @     �Y@      @      @      @      @      L@      B@              $@      @      @                       @     �M@       @      g@      �?       @      �?       @     @T@     �A@              (@�t�bub�     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�Y�fhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?}��� ��?�	           ��@       	                    �?{z>�?           ��@                          �0@���\+�?w           �@                           @�m��1�?             :@������������������������       ��&5D�?
             1@������������������������       ��2�tk~�?             "@                            @*}��?g           8�@������������������������       ����ٽp�?�            �t@������������������������       �4"�L'T�?�            �o@
                          �0@��k���?�           �@                           �?R����?            �@@������������������������       ��s�n_�?             *@������������������������       �333333�?             4@                          �<@�閴y�?t           �@������������������������       �:��d+��?"           �@������������������������       �Yo���-�?R             `@                            @�M�r��?�           ʡ@                            �?��́�
�?�           (�@                           �?K;l�?��?1           ԓ@������������������������       ��7���#�?�           x�@������������������������       �R�����?�           0�@                           �?ͪ�%\u�?S           ��@������������������������       ����{ �?m             g@������������������������       ��}{���?�            �u@                           �?^���W�?#           �}@                          �2@�#Y9���?[             c@������������������������       �I�7�&��?&             N@������������������������       ��1�e,�?5            @W@                           @Y��r��?�             t@������������������������       �H�%s��?W            �a@������������������������       ��~�~�?q            �f@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      B@     �A@     �@@     @V@     P�@      H@     �@      2@      @     @S@     �Q@     x�@     ؀@      *@     �p@     �W@      .@      9@      0@     �B@     �o@      &@     (�@      &@      @     �@@      2@     0r@     �i@      @     �X@     �A@      @      5@      @      7@      W@       @     @d@      @      �?      4@      @     �W@      V@       @      F@                                      �?      �?                                      �?      @      @      &@               @                                                                                      �?      �?      @       @                                                      �?      �?                                               @              @               @     �A@      @      5@      @      6@     �V@       @     @d@      @      �?      3@      @     �U@     @S@       @      E@      2@       @      &@      @      &@     �K@      �?     �T@      @              1@      @      G@     �B@      �?     �@@      1@      @      $@              &@      B@      �?     �S@      @      �?       @             �D@      D@      �?      "@     �M@      $@      @      "@      ,@     `d@      "@     0v@      @      @      *@      (@     �h@      ]@      @     �K@       @                                      &@              @                                      "@      @              @       @                                      @              �?                                      @      �?               @                                               @               @                                      @      @              �?     �L@      $@      @      "@      ,@      c@      "@      v@      @      @      *@      (@     �g@     �[@      @      J@     �J@      "@      @      "@      ,@     @^@      @     �r@      @              *@       @      e@      Z@      @     �F@      @      �?                              ?@       @     �I@              @              @      3@      @              @     @Z@      5@      $@      1@      J@     �x@     �B@     ��@      @      @      F@      J@     �|@     �t@      @     �d@     �V@      .@      @      .@      F@     ps@      A@      z@      @      @     �C@     �G@     pu@     �q@      @     �a@     �L@      (@      @      &@      9@     �l@      7@      u@      @       @      1@      B@     �p@      d@      @     @S@     �B@      @      @      @      1@     �\@      .@     @`@      �?       @      $@      3@      `@     �V@       @      C@      4@      @      �?      @       @     @\@       @     �i@      @              @      1@     @a@     �Q@      @     �C@      A@      @      �?      @      3@     �T@      &@      T@              �?      6@      &@      S@     �^@       @      P@      0@              �?      @      @      ;@      @      5@                      @      @      @@      H@              4@      2@      @                      .@      L@       @     �M@              �?      2@      @      F@     �R@       @      F@      ,@      @      @       @       @      U@      @     �b@      �?              @      @     @]@      J@              9@      "@       @                       @      :@       @     �A@                      �?      �?     �E@      5@              &@       @                                      @              2@                                      <@      @               @      @       @                       @      4@       @      1@                      �?      �?      .@      1@              "@      @      @      @       @      @      M@      �?     �\@      �?              @      @     �R@      ?@              ,@       @              @       @      @      ,@              O@                                     �A@      *@              @      @      @                       @      F@      �?     �J@      �?              @      @     �C@      2@              "@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ4��/hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?}�����?�	           ��@       	                    @����?^           ��@                           �?J�2Q��?�           ��@                            �?�kL1���?�            �y@������������������������       �p��:9��?K            @^@������������������������       �6��?�?�            0r@                            @H���j��?�           ��@������������������������       �&���^�?q            �@������������������������       �yA+�R�?e            �c@
                           @�K�tF�?�           x�@                           @�7W��5�?}           ��@������������������������       �9�G�V^�?�             q@������������������������       �����i��?�            pt@������������������������       �r�q��?             8@                            @�;����?X           Ġ@                          �0@��맃��?�           ܗ@                            �?)O���?1             R@������������������������       �'y�Y�?#             K@������������������������       �����K�?             2@                            �?ү��gr�?�           ��@������������������������       �������?�           ��@������������������������       ���H�N��?�            �t@                           @��a�8(�?�           X�@                           @&R����?&           �}@������������������������       �2(�D�"�?�            Pv@������������������������       ����B�?D            �\@                          �3@<9�۸,�?_            `b@������������������������       �v�)�Y7�?            �B@������������������������       �>���	��?G            �[@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        k@     �A@      >@      4@     �Z@     ؄@     �@@     ��@      .@      @     �U@     �O@     ��@     �@      ?@     �o@      Z@      7@      5@      @     �M@     �s@      5@     �{@       @      @      F@      C@     �r@     @m@      3@      `@     @S@      $@      ,@      @     �G@     `h@      @     �r@      @       @      @@      9@     �k@     �`@      @     �Q@      9@      @      "@      �?      &@     �M@       @      _@      @              1@       @      N@     �K@       @      =@      @                      �?      @      0@              I@                      @      @      *@      (@       @      "@      4@      @      "@               @     �E@       @     �R@      @              ,@      �?     �G@     �E@              4@      J@      @      @      @      B@      a@      �?     �e@       @       @      .@      1@      d@      T@      @     �D@      G@       @      @      @      A@      [@             �^@       @       @      $@      1@     �^@     @P@      @      A@      @      @      �?               @      <@      �?      I@                      @              C@      .@              @      ;@      *@      @       @      (@     �]@      2@     �b@      �?       @      (@      *@     �S@     �X@      ,@      M@      ;@      *@      @       @      (@      ]@      *@      b@      �?       @      (@      *@     �R@      X@      ,@     �I@      3@      @      @      �?       @      I@      @      M@              �?       @      @      B@      I@      @      6@       @      @      �?      �?      @     �P@      @     �U@      �?      �?      $@      $@     �C@      G@      $@      =@                                               @      @      @                                      @      @              @     @\@      (@      "@      *@      H@      v@      (@     �@      @              E@      9@     �z@      q@      (@     @_@     �V@      $@      @      $@      C@     �o@      (@      {@      @             �D@      4@     �q@     �j@      $@     �Y@      @                      �?              9@              "@                      �?      �?      &@      @              (@      @                                      2@              "@                      �?      �?      "@      @              $@       @                      �?              @                                                       @      @               @     @U@      $@      @      "@      C@     �l@      (@     pz@      @              D@      3@      q@      j@      $@     �V@     �O@       @      @       @      5@      f@      @     v@      @              .@       @     �m@      d@       @     �H@      6@       @      @      �?      1@      J@      @     �Q@      �?              9@      &@      A@      H@       @     �D@      7@       @      @      @      $@     @Y@             @n@       @              �?      @     �a@     �M@       @      7@      2@      �?      @      @      @     �O@              i@                      �?      @      [@     �F@              3@      $@      �?      @      @      @      J@             �a@                      �?      @     �U@      A@              1@       @                                      &@             �N@                                      6@      &@               @      @      �?                      @      C@             �D@       @                       @     �A@      ,@       @      @      @                              @      @              @                                      .@      @                      �?      �?                             �@@              A@       @                       @      4@      &@       @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�l#*hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�gD���?�	           ��@       	                   �;@�h��?�           ��@                          �0@L�b�a�?&           &�@                           �?@DE�"��?n            �d@������������������������       ����!��?>            �U@������������������������       �ףp=
W�?0             T@                            �?�8v��?�           ء@������������������������       �������?=           x�@������������������������       �a�W���?{           p�@
                           �?�:����?�            ps@                           �?!��wy��?U            @a@������������������������       ��8��8��?             8@������������������������       ���8='n�?J            �\@                           @x�����?p            �e@������������������������       ���HHI�?J            �[@������������������������       �z8,���?&             O@                           �?�Ĩb�C�?�           ��@                           @�C�A�6�??           �@                          �>@�O�[^�?           �y@������������������������       �DӵX?�?�            px@������������������������       ���(\���?             4@                           @_�-J��?<            �W@������������������������       �ȖLy�r�?*            �P@������������������������       �����>�?             <@                           @�t�8�?�           (�@                           �?]�M�?�            �x@������������������������       �@��5-�?�            �o@������������������������       �zD94_�?]             b@                           @�-7���?�            �n@������������������������       �z�����?q            `g@������������������������       ��P�a�r�?%             N@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @j@      @@      C@      9@      ^@     x�@      >@     �@      .@       @     �S@     �L@     �@     �@      .@     �m@      d@      8@      =@      5@      Y@     0|@      9@     `�@      &@      @      P@     �J@     8�@     �w@      *@     @h@     �b@      3@      <@      4@     �W@     �y@      6@     ��@      "@      @     �M@      H@     �|@     �u@      *@     �e@      @      �?      @       @      &@     �C@      @      8@               @       @      @      ;@      8@      �?      1@       @      �?      @              &@      1@      @      $@               @       @              *@      &@      �?      $@      @                       @              6@              ,@                              @      ,@      *@              @     �a@      2@      9@      2@     �T@     Pw@      2@     ��@      "@      @     �L@     �E@      {@     0t@      (@     �c@     �X@      ,@      (@      .@      G@     `r@      .@      }@      @      �?      F@      7@     �t@      l@       @     �X@     �F@      @      *@      @     �B@     �S@      @      Z@      @       @      *@      4@     @Y@     �X@      @      M@      (@      @      �?      �?      @     �C@      @      _@       @              @      @      M@      >@              4@       @      @      �?              @      .@             �H@                       @              6@      2@              ,@                                              @              0@                       @                      �?              �?       @      @      �?              @      &@             �@@                                      6@      1@              *@      @       @              �?              8@      @     �R@       @              @      @      B@      (@              @      @       @              �?              1@      @     �B@       @                      @      <@       @              @                                              @              C@                      @       @       @      @                      I@       @      "@      @      4@     �i@      @      w@      @      @      ,@      @     �q@      `@       @     �F@      =@       @      @      @      (@      Z@      @     �a@      �?       @      "@       @      X@     @Q@       @      5@      9@      @      @      @      &@     @V@       @     �Y@      �?              @       @      U@      L@       @      3@      5@      @      @      @      &@     @U@       @      X@                      @             �T@      L@              3@      @                                      @              @      �?                       @      �?               @              @      @                      �?      .@      �?     �C@               @       @              (@      *@               @      @      @                      �?      (@              7@               @                       @      (@              �?                                              @      �?      0@                       @              @      �?              �?      5@              @      �?       @      Y@       @     `l@      @      �?      @       @     `g@     �M@              8@      .@              @      �?      @     �D@              c@      �?      �?       @      �?      `@      ;@              2@      $@               @      �?      @      <@             �W@      �?      �?       @      �?      R@      4@              2@      @              �?              @      *@             �M@                                     �L@      @                      @               @               @     �M@       @     �R@       @              @      �?      M@      @@              @      @               @               @      F@       @     �H@                              �?     �I@      9@              @                                              .@              9@       @              @              @      @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJF�dhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�"��@j�?�	           ��@       	                     �?�a�H`��?�           �@                          �=@�yoֲ��?L           ֠@                           �?֯IQ��?           ��@������������������������       �0�{��I�?:           P�@������������������������       ��ݓ��?�           ̑@                          �@@(Qq����?I            �[@������������������������       ���rm��?9            �U@������������������������       �36�v[�?             7@
                           @��x9��?�           �@                          �4@+��R��?w           0�@������������������������       �0�\[
�?�            ps@������������������������       �e�MgHR�?�            �r@                           @�I��I��?$             N@������������������������       �O�mL�?            �E@������������������������       �� =[y�?             1@                           �?
4�F��?�           �@                           �?��$jD�?%           �{@                          �2@���^B��?g             b@������������������������       ��qǱ�?"             H@������������������������       �������?E             X@                          �0@\#Y�z��?�            �r@������������������������       ��������?             .@������������������������       �>�w��V�?�            �q@                          �;@©s�7R�?�           �@                          �9@�5�K��?X           ��@������������������������       ��f��)��?2           �~@������������������������       �Z�N���?&            �P@                           @:��C#�?/            �T@������������������������       �ʬJ�h�?            �G@������������������������       ��Hx�5�?             B@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      >@      @@      4@     �Z@     p�@     �E@     ȑ@      1@      &@     �M@     �J@     H�@     �@      6@     �p@     �c@      7@      ;@      2@      V@     �@     �B@     ��@      (@      "@      I@      H@     �~@     �w@      3@     �k@     @]@      .@      6@      0@     �O@     Py@      <@     ��@      @       @      ?@      9@     `x@      q@      &@      c@      ]@      ,@      6@      0@     �M@     �x@      :@     Ȁ@      @       @      >@      8@     �w@     �p@      &@     �b@      K@      @      2@      $@     �A@     @h@      *@     �g@      @       @      4@      (@     `c@     �[@      @      T@      O@      "@      @      @      8@     �h@      *@     �u@       @              $@      (@     �k@     @c@      @     @Q@      �?      �?                      @      (@       @     �M@      �?              �?      �?      ,@      $@              @      �?      �?                      @      $@       @      J@      �?              �?              &@       @               @                                               @              @                              �?      @       @               @      E@       @      @       @      9@      [@      "@     @`@      @      @      3@      7@     @Z@     @[@       @     @Q@     �C@       @      @       @      9@      W@      "@     @[@      @      @      2@      7@      X@     @Z@       @      P@      4@      @      �?      �?      ,@     �K@       @     �B@              @      ,@      0@      B@     �N@       @      C@      3@      @      @      �?      &@     �B@      @      R@      @       @      @      @      N@      F@              :@      @                                      0@              5@      �?              �?              "@      @              @      @                                      *@              ,@      �?              �?               @      �?               @                                              @              @                                      �?      @              @     �F@      @      @       @      3@     �e@      @     �y@      @       @      "@      @     @k@     ``@      @      E@      <@      @      @              *@     @Q@      @     �`@      @      �?      @      @     �U@     �J@      @      =@      "@      �?       @               @      9@      �?      >@                      @      �?      A@      4@              .@      @               @                      (@              $@                                      0@      @               @      @      �?                       @      *@      �?      4@                      @      �?      2@      1@              *@      3@      @       @              &@      F@      @      Z@      @      �?      @       @      J@     �@@      @      ,@      �?                                       @       @                               @              @                      @      2@      @       @              &@      E@      �?      Z@      @      �?      �?       @      H@     �@@      @      $@      1@      @      �?       @      @      Z@       @     `q@       @      �?       @       @     �`@     �S@              *@      0@      @      �?       @      @     �T@       @     �l@       @               @       @      _@     �R@              *@      0@      @      �?       @      @     @S@       @      j@       @               @       @     @Y@      N@              &@                                              @              6@                                      7@      .@               @      �?                              �?      6@             �G@              �?                       @      @                      �?                              �?       @             �B@              �?                      @                                                                      4@              $@                                      @      @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�@@hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@M��xp�?�	           ��@       	                     @��l.��?�           �@                            �?�?J$���?9           J�@                          �0@kB��G~�?�           T�@������������������������       �< G58m�?Q             _@������������������������       ����b�?g           d�@                          �4@RCXh"��?�           ��@������������������������       ����O���?�            �s@������������������������       ��Cٗ�K�?�             q@
                           @J��f�?a           �@                          �5@.j��[�?V           ��@������������������������       ���jw�?f           ��@������������������������       �F�;�
�?�            �w@������������������������       �$�ɜoB�?             1@                           �?�r$a,��?           |@                            �?);�h�?j            �d@                          �=@�"��U>�?             ?@������������������������       �I�O���?             7@������������������������       �      �?              @                            @[y�����?U             a@������������������������       ��.��6i�?2            �S@������������������������       ���9 �"�?#            �L@                          �@@��U��?�            �q@                          @@@<��E��?�            �o@������������������������       ��/K�]l�?�             m@������������������������       �"�����?
             5@                             @��>�Q�?             =@������������������������       �<+	���?             .@������������������������       �T�r
^N�?	             ,@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@     �A@      C@      8@     �\@     �@      F@     ��@      4@      &@     �P@      L@     ��@     ��@      3@      n@     `e@      =@     �A@      7@     �X@      �@      D@     ��@      0@      $@      N@     �I@     Є@     P@      .@     �j@      a@      1@      :@      .@     @T@      {@      ?@     X�@      (@      $@     �H@     �C@      |@     �v@      ,@     @e@     @Z@      (@      .@      .@     �I@     pv@      7@     �@      @              <@      ;@     @v@     �o@      $@      [@      @              �?       @       @      5@              *@      �?                      @     �@@      <@              $@     �Y@      (@      ,@      *@     �E@      u@      7@      @      @              <@      7@     0t@      l@      $@     �X@      ?@      @      &@              >@     �R@       @     �[@      @      $@      5@      (@     �W@     �\@      @      O@      6@      �?      @              &@     �H@      @      H@              @      .@      "@      C@     �P@      @      D@      "@      @      @              3@      :@      @      O@      @      @      @      @      L@      H@              6@     �A@      (@      "@       @      1@     �a@      "@     0u@      @              &@      (@      k@     �`@      �?     �F@     �A@      (@      "@       @      1@     �`@      "@      u@      @              &@      (@     �j@     ``@      �?     �F@      3@       @      @       @      0@      R@      @     �j@      @              &@      $@     �]@     �R@              >@      0@      @       @              �?      O@      @     �^@      �?                       @     �W@     �L@      �?      .@                                               @              �?                                      @      @                      2@      @      @      �?      0@     @P@      @     �e@      @      �?      @      @     �U@      ?@      @      9@      $@      @      @              @      3@              J@                      @             �@@      3@       @      (@                                       @      @              .@                      �?              @      �?              �?                                      �?      @              $@                      �?              @                      �?                                      �?                      @                                      �?      �?                      $@      @      @              @      ,@             �B@                      @              ;@      2@       @      &@      @      @       @              �?      &@              .@                      @              1@      &@               @      @              �?              @      @              6@                                      $@      @       @      @       @                      �?      "@      G@      @     �^@      @      �?       @      @     �J@      (@       @      *@      @                      �?      "@      G@      @      [@      @      �?       @      @     �E@      &@       @      $@      @                      �?       @     �E@      @     �Y@       @               @      @     �E@      &@              $@                                      @      @              @       @      �?                                       @              �?                                                      ,@                                      $@      �?              @                                                              @                                      @      �?              @      �?                                                       @                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��51hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             @��|k�?�	           ��@       	                    �?=�4�h�?           �@                           �?�l�P��?�           ��@                          �9@��#m�?�           ��@������������������������       ������?]           0�@������������������������       �g�vPا�?2            �R@                          �;@Z���ll�?9           �@������������������������       ���^$ʔ�?           �{@������������������������       ������?(            �N@
                           �?"�Ɔ[��?@           ��@                          �<@��9�C�?�            �l@������������������������       �u�L]���?�            �j@������������������������       �{�/��>�?
             1@                          �3@��z�r�?�           �@������������������������       �H�2�E�?            {@������������������������       ��a�?�           P�@                           @h��n�W�?�           ��@                          �0@�p],�?J           �@������������������������       �\���(\�?             4@                          �<@]+���??           �~@������������������������       ��2\G�?            {@������������������������       �ϊF�y�?'             N@                           @�U��"\�?d           ��@                           @��#��?�           `�@������������������������       ���C��0�?*           �}@������������������������       �Qf����?`            �a@                          �:@�-�I��?�             u@������������������������       �fx��R%�?�            `p@������������������������       ��6<�v$�?-            �R@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@     �A@      F@      <@      U@     ��@      A@     L�@      (@      @     �S@     �P@     �@     �~@      3@     �n@     @a@      1@      A@      1@     �P@     pz@      2@     8�@       @       @      G@      A@     ��@     Pp@      $@      d@      O@      (@      ?@      "@      F@      k@      @     �p@      @      �?      6@      0@      l@     �`@      @      U@     �D@      "@      1@       @      3@      [@      @     @a@      @      �?      ,@      $@      ]@     �R@      @      M@     �A@      "@      1@      @      3@      Y@      @      \@      @      �?      (@      "@     �W@      R@      @      I@      @                      �?               @              :@                       @      �?      5@       @               @      5@      @      ,@      �?      9@      [@             �_@      �?               @      @      [@      M@      �?      :@      3@      �?      &@      �?      8@     �W@             �X@      �?               @      @     @Y@      K@      �?      9@       @       @      @              �?      *@              <@                                      @      @              �?      S@      @      @       @      7@     �i@      (@     �y@      @      �?      8@      2@     s@      `@      @      S@      (@       @                      @     �@@             �H@                      @      @     �P@      7@              ;@      &@       @                      @      ;@              G@                      @      �?     �P@      7@              :@      �?                               @      @              @                              @      �?                      �?      P@      @      @       @      1@     �e@      (@     �v@      @      �?      1@      ,@     �m@     �Z@      @     �H@      2@                      @      @     �P@      @     ``@                      @      "@     �]@      J@       @      4@      G@      @      @      @      *@      [@      "@     `m@      @      �?      (@      @     �]@      K@      @      =@     �P@      2@      $@      &@      1@     @m@      0@     �z@      @      �?      @@      @@     q@     @m@      "@      U@      ?@      @      @      @      @      S@      @     �d@       @              ,@      *@     �T@     �Q@       @     �A@      �?                                      �?                                      �?              @      @               @      >@      @      @      @      @     �R@      @     �d@       @              *@      *@     �S@     �P@       @      ;@      >@      @      @      @      @     @P@      @      a@      �?              @      *@     @Q@     �P@      �?      9@                                              $@              ?@      �?              @              "@              �?       @      B@      *@      @      @      (@     �c@      *@     Pp@       @      �?      2@      3@     �g@     �d@      @     �H@      >@      $@      @      �?      @     �[@      $@     �b@              �?      &@      2@     �]@      ]@      @      :@      2@      @      @      �?       @     �T@      @      `@              �?      @      .@      V@     �X@      @      2@      (@      @      �?              @      ;@      @      6@                      @      @      >@      2@       @       @      @      @       @      @      @      H@      @     �[@       @              @      �?      R@      H@              7@      @      @       @       @      @      C@      @      R@       @              @      �?      M@      F@              7@                              @              $@             �C@                      @              ,@      @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ/y`hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @��U���?�	           ��@       	                    @Ъc��?�           ��@                           �?�dF��?#           &�@                          �0@D���X�?9           ��@������������������������       ���.��?/             S@������������������������       �K+�}4�?
           H�@                            �?�HDR���?�           x�@������������������������       ���o+>�?@           ��@������������������������       ��u�{��?�            �p@
                          �;@ԗ�gۙ�?�           ��@                           !@+�:�G��?x           (�@������������������������       �c��F��?q           Ȃ@������������������������       ��q�q�?             (@                          �=@�K!�H��?2            �T@������������������������       �n�����?             >@������������������������       ���B�<�?            �J@                           �?�Λw3�?�           ��@                           @"�֖�K�?4           0~@                          �;@(�Tw��?�            �s@������������������������       �`:
:�?�            pq@������������������������       �<Cb�ΐ�?            �@@                          �:@�|rC(Q�?k            `e@������������������������       ��������?X            �a@������������������������       �*#|����?             ?@                          �=@�W�2/�?�           ؄@                          �0@��n��?v           ��@������������������������       �x9/���?             <@������������������������       �1���nG�?g           �@                          �@@� Ce���?             N@������������������������       �})Z6K�?            �G@������������������������       ��	j*D�?             *@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `j@      >@     �@@      8@     @^@     ��@      7@     �@      7@      $@      R@      O@     ؆@     �@      2@     �p@     @d@      6@      9@      2@      X@     �~@      3@     x�@      4@      @      P@     �I@     �~@     �w@      .@     @j@     �`@      1@      6@      0@     �S@     �w@      (@     �@      &@       @      J@     �B@     Pw@     �n@       @     `e@     @Q@       @      ,@      @     �A@      c@      @     �g@      $@              9@      1@     �e@     �[@      �?      S@       @      �?      �?       @      @      .@      �?      @      @               @       @      .@      .@              @     �P@      �?      *@      @      =@      a@      @     �f@      @              7@      .@     �c@     �W@      �?      R@      P@      .@       @      "@      F@     �l@      @     �s@      �?       @      ;@      4@     �h@      a@      @     �W@     �E@      *@      @      "@      ?@     �g@      @     �p@      �?              *@      &@      d@     @Y@      @     �N@      5@       @      @              *@     �C@      @      J@               @      ,@      "@     �C@      B@      �?      A@      =@      @      @       @      1@     @\@      @     �f@      "@       @      (@      ,@      ^@     �`@      @     �C@      ;@      @      @       @      1@     �X@      @     �b@      "@       @      (@      *@      X@     �_@      @     �C@      9@      @      @       @      1@      W@      @     �b@      "@       @      (@      *@      X@     @_@      @      C@       @                                      @                                                               @              �?       @                                      ,@              A@                              �?      8@       @                                                              $@              ,@                                      @       @                       @                                      @              4@                              �?      4@      @                     �H@       @       @      @      9@     �h@      @     @y@      @      @       @      &@     �m@     @_@      @      K@     �@@      @      @      @      *@      V@      @     �a@      �?       @      @      @     @V@      N@             �@@      3@      �?      @      @       @      P@             @U@      �?              @      �?     �O@      F@              0@      1@      �?      @      @      @     �O@             �R@                      @      �?      J@      D@              *@       @                              �?      �?              $@      �?                              &@      @              @      ,@      @      �?              @      8@      @      L@               @              @      :@      0@              1@      "@      �?      �?              @      8@      @     �B@               @              @      7@      .@              1@      @       @                      �?                      3@                                      @      �?                      0@      @      @      @      (@     �[@      �?     pp@       @      @      @      @     �b@     @P@      @      5@      0@      @      @      @       @     �V@      �?     �n@       @              @      @     �`@     @P@      @      5@                                               @              4@                                      @       @              �?      0@      @      @      @       @     @V@      �?     `l@       @              @      @      `@     �O@      @      4@                                      @      3@              0@              @                      1@                                                              @      3@              (@              @                       @                                                                                      @                                      "@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJU��WhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �:@x�\���?�	           ��@       	                    �?�C d��?0           �@                            @P�	�U�?�           t�@                           �?A��g���?�           <�@������������������������       ���[�y�?V            `a@������������������������       �Z�3
��?W            �@                           @#�\D��?�            �x@������������������������       �>�cp>�?�            �t@������������������������       ��)񎴠�?0            �Q@
                          �0@Z�D��'�?�           ��@                            @0�F����??            �W@������������������������       �2��k�?1             S@������������������������       �0\�Uo��?             3@                           @pәJ
!�?E           0�@������������������������       �7�}����?�           ��@������������������������       ��9X�m�?^           X�@                           �?g�[[e�?p           �@                           �??��̭��?�            �m@                           �?�Ls?���?5            �U@������������������������       ��w@	��?            �I@������������������������       � )O��?             B@                           @S^?����?c            �b@������������������������       ���%l��?R             `@������������������������       ���J��?             6@                          �=@��,\�?�            0u@                          �;@��x���?u            �e@������������������������       ��H���?2            �R@������������������������       �8gDio��?C             Y@                           @���|��?c            �d@������������������������       �""""""�?H             ^@������������������������       ���ˠ�?             F@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @h@      A@     �D@      ?@     �Z@     h�@      A@     l�@      $@      @     �Q@     �P@     �@     8�@      =@     �r@      f@      <@     �A@      <@     �V@     ؀@      =@     p�@      "@      @     �O@      O@     8�@     }@      :@     �o@     �V@      *@      @@      *@     �I@     �o@      .@     �u@      @      @      <@      >@     �p@     @j@      1@      ^@     �P@      "@      7@      *@      D@     �h@      &@      l@      @      @      4@      =@     �f@     `c@      1@     �Y@      @       @      @              @      .@      �?      E@      @              @      �?      >@      *@              *@     �O@      @      4@      *@     �A@     �f@      $@     �f@      @      @      ,@      <@     �b@     �a@      1@     �V@      7@      @      "@              &@      L@      @      ^@                       @      �?     �V@     �K@              1@      5@      @      "@               @      G@      �?     @V@                       @      �?     @S@      I@              .@       @      �?                      @      $@      @      ?@                                      *@      @               @     �U@      .@      @      .@      D@     �q@      ,@     ��@       @             �A@      @@     �u@     �o@      "@     �`@      �?                       @              7@              5@                      �?       @      5@      *@              &@      �?                       @              5@              &@                      �?       @      1@      &@              $@                                               @              $@                                      @       @              �?     �U@      .@      @      *@      D@     pp@      ,@     �@       @              A@      >@     0t@     @n@      "@     @^@      L@      $@      �?      $@      6@      h@      @     0w@       @              5@      2@      m@     @d@      @     �R@      >@      @       @      @      2@     �Q@      "@     �e@                      *@      (@     �V@      T@       @      G@      1@      @      @      @      .@     �T@      @     �i@      �?               @      @     �]@      K@      @     �H@      &@      @      @      @      $@      >@      �?     �Q@      �?              @       @     �B@      =@              =@       @              �?      @      @      "@              >@      �?              @       @      3@      @              @                      �?      @      @      @              *@      �?              @       @      (@      �?              @       @                                      @              1@                                      @      @              @      "@      @      @              @      5@      �?      D@                      �?              2@      9@              7@       @      @      @               @      2@      �?      C@                      �?              ,@      1@              6@      �?      �?      �?              �?      @               @                                      @       @              �?      @      �?                      @      J@      @     �`@                      @      @     @T@      9@      @      4@      @      �?                       @      9@              S@                      @       @      ?@      4@       @      "@       @      �?                       @       @              9@                               @      5@      "@              @       @                                      1@             �I@                      @              $@      &@       @      @       @                              @      ;@      @     �M@                      �?      �?      I@      @      �?      &@       @                              @      6@      @      G@                      �?              <@       @      �?      &@                                              @              *@                              �?      6@      @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ*� hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �1@P]�����?�	           ��@                           �?�[�l	O�?�           p�@                           @Y:]�$�?�            �t@                           @�R��?�            �s@������������������������       ��M��S�?�            �k@������������������������       ��x���?<             W@������������������������       ��F����?             1@                           �?ǻ���?�            0t@	       
                     �?5_�g���?             F@������������������������       ���ճC��?             6@������������������������       ��!pc��?             6@                            �?��߈���?�            pq@������������������������       � ���N�?i             e@������������������������       ��{�S��?G            �[@                            @8�i�F�?+           v�@                            �?�2�L��?�           ̡@                           �?�+��yT�?K           ��@������������������������       ��9��?�           �@������������������������       �䲣����?�           �@                           @C�9s;��?_           �@������������������������       ���Gb��?�            @p@������������������������       �y�2ѫ6�?�            �s@                          �2@mԩDo��?�           ��@                           �?dj`��?a            @c@������������������������       �ԭ�a�2�?,             R@������������������������       �s��;��?5            �T@                          �=@qm�����?            ؉@������������������������       ���Rv#��?�           ��@������������������������       ��l'V3�?7            �R@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      ;@      F@      ?@     �[@     ��@      B@     <�@      :@       @      T@      K@     @�@     p@      6@     �p@     �I@      @      ,@      �?      4@     �\@      "@     �b@      �?       @      5@      0@     �V@      ]@      @      E@      8@      @      *@      �?      2@     �J@       @     �M@      �?       @      &@      *@      C@     �L@      �?      <@      8@      @      (@      �?      &@     �J@       @      M@      �?       @      &@      *@      C@     �I@      �?      :@      3@      @      $@      �?       @      ?@      @     �@@                      $@      &@     �@@      B@      �?      5@      @               @              @      6@      @      9@      �?       @      �?       @      @      .@              @                      �?              @                      �?                                              @               @      ;@              �?               @     �N@      �?     �V@                      $@      @     �J@     �M@       @      ,@      "@                               @      @              @                                      ,@       @       @       @      @                                      @              @                                      $@                       @      @                               @      @              @                                      @       @       @              2@              �?                      K@      �?      U@                      $@      @     �C@     �L@              (@      (@                                      <@      �?     �M@                      @              8@      =@              &@      @              �?                      :@              9@                      @      @      .@      <@              �?     @e@      7@      >@      >@     �V@     0�@      ;@     Џ@      9@      @     �M@      C@     h�@     0x@      3@     �l@      _@      *@      2@      ;@     �R@     �v@      6@     0�@      ,@      @     �J@      B@     Px@      r@      2@     �g@     �S@      (@      .@      5@      I@     0r@      1@     @�@       @              @@      3@     �r@     @i@      *@     �^@      :@       @      @      (@      6@      Y@      @      h@      �?              5@       @      \@     �X@      �?      P@      J@      @      &@      "@      <@     �g@      *@     �t@      @              &@      &@     `g@      Z@      (@      M@      G@      �?      @      @      8@     �Q@      @     �_@      @      @      5@      1@     �V@     �U@      @     �P@      0@      �?       @       @      "@      >@             �O@      @       @      @      �?     �G@     �D@             �B@      >@              �?      @      .@      D@      @     �O@      @      @      .@      0@     �E@     �F@      @      >@      G@      $@      (@      @      1@     �c@      @     @w@      &@              @       @      i@     �X@      �?      D@      @               @      @      �?      6@              K@                      �?              G@      1@              @      @               @      �?      �?      @              6@                                      =@      @              �?      �?                       @              .@              @@                      �?              1@      &@              @      E@      $@      $@              0@     �`@      @     �s@      &@              @       @     @c@     �T@      �?      B@     �A@      $@      $@              (@     �^@      @      r@      @              @       @     �`@     �T@              B@      @                              @      (@              <@      @                              3@              �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��fhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@J�Ӂ��?�	           ��@       	                    �?(ϵҴ�?h           ު@                          �8@�J��Y�?�            �@                           @��ο^�?F           Ȕ@������������������������       �o��O*R�?n           ��@������������������������       �Fĝr�P�?�           ��@                           @��$���?�            �j@������������������������       ���J^��?y            �h@������������������������       �     ��?	             0@
                            @څ�{M�?�           ��@                          �0@�DLCa|�?L           L�@������������������������       ��@��Ƅ�?2            �U@������������������������       ��ʳ#gf�?           ��@                          �9@,�j��?T           ��@������������������������       �ڔl�W��?1           �}@������������������������       �n�Y���?#            �L@                          �>@V�.���?)           �}@                           @��7Z�?�            t@                           @|�l�]V�?�             q@������������������������       �MB_���?�            �k@������������������������       ���As��?             �I@                           �?f�Sc��?            �H@������������������������       �B{	�%��?             2@������������������������       �tH�����?             ?@                          �?@�/O��W�?a             c@                           �?DzA��d�?            �G@������������������������       �~IO���?            �B@������������������������       �R���Q�?             $@                            �?XA�H��?E            �Z@������������������������       ���]�&�?&            �L@������������������������       ��/@f�~�?            �H@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      >@      F@      7@     @W@     (�@      8@     ��@      4@      "@     @P@     �O@     ��@     ��@      2@      q@     �f@      9@     �E@      5@     �V@     �@      7@     X�@      &@      @     �N@     �L@      �@     �@      &@     �n@     �V@      2@      >@      &@     �K@     �q@      1@      u@      "@      @      >@      A@     `q@      k@      @     �_@     @T@      ,@      >@      @     �I@     `m@      *@     �r@      @      @      =@      @@      m@     �e@      @      [@     �C@      @      0@       @      >@      W@       @     �`@       @      �?       @      (@     �V@     @W@              E@      E@      $@      ,@      @      5@     �a@      @      e@      @      @      5@      4@     �a@     �T@      @     �P@      "@      @              @      @     �F@      @     �@@      @              �?       @     �F@     �D@              3@      "@      @              @      @     �E@      @      :@      @              �?       @     �F@      D@              *@                                               @              @                                              �?              @     @W@      @      *@      $@     �A@     Pt@      @     ؀@       @              ?@      7@     �x@     r@      @     �]@     �S@      @      @      @      ?@     �n@      @     �v@       @              =@      1@     �n@      k@      @      Y@      @                      �?              ;@              @                      @      �?      ,@      5@              @     @R@      @      @      @      ?@     �k@      @     �v@       @              :@      0@     �l@     �h@      @     @W@      ,@              @      @      @     �S@             �e@                       @      @     @c@      R@      �?      3@      ,@              @      @      @     �Q@             �c@                       @      @     �_@     �P@      �?      2@                                               @              .@                                      ;@      @              �?      7@      @      �?       @      @      R@      �?     @h@      "@       @      @      @      U@     �A@      @      :@      *@      @      �?       @      �?      H@             `b@       @              @      �?     �J@      8@       @      2@      *@      @      �?       @      �?     �E@              \@       @              @      �?      H@      8@       @      .@      $@      @      �?              �?     �B@              X@       @              @      �?      =@      5@       @      *@      @                       @              @              0@                                      3@      @               @                                              @             �A@                      �?              @                      @                                              @              @                      �?              @                      @                                              �?              <@                                       @                              $@                               @      8@      �?     �G@      @       @              @      ?@      &@      @       @                                      �?      (@      �?      &@                               @      @      @      @      @                                              "@      �?       @                               @      @      @      @      @                                      �?      @              @                                       @                      �?      $@                              �?      (@              B@      @       @              @      8@       @       @      �?      @                                      @              5@       @                      �?      0@       @                      @                              �?      @              .@      @       @               @       @               @      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�je-hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx                             �?#���2Z�?�	           ��@       	                    @�4�E}�?E           �@                          �<@�E�����?�           ��@                            @�5��*��?Q           ��@������������������������       �0R�j�?�           ��@������������������������       ������?�            �s@                           �?fP*L��?8             V@������������������������       ���P���?            �A@������������������������       �����#8�?$            �J@
                            @թ�B�?�           0�@                           @�ۗ�s�?q           ��@������������������������       �|�X�W�?           p|@������������������������       ��V���?R            @a@                          �2@�!p4l�?K            @]@������������������������       ��i�̄�?            �D@������������������������       �D�n�3�?/             S@                           !@�eN���?W           �@                          �;@^���?M           �@                           @k�B���?�           ��@������������������������       �.�����?�           ,�@������������������������       �lF�Ǟ��?�           �@                           �?��/�@�?�            �p@������������������������       �c��gS~�?             =@������������������������       ���Iu(��?�            �m@������������������������       �
ףp=
�?
             4@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `j@      6@      H@      8@     @Y@     ��@      >@     ��@      5@      @      Q@     �P@     �@     �@      .@     `l@     �Z@      .@      C@      (@     �P@     �s@      4@     �z@       @       @      7@      @@     @r@     @m@      "@     @]@     �N@      "@      8@       @      E@      g@      *@     `q@      @      �?      1@      &@     `d@     �`@      @      N@     �G@       @      6@       @     �C@     �f@      *@     �m@      @      �?      *@      $@      c@      `@      @      L@     �D@      @      0@       @      ;@      ]@      &@     @a@      @              *@      @     @V@     �U@      @     �D@      @      @      @              (@      P@       @     @Y@              �?              @      P@      E@              .@      ,@      �?       @              @      @             �C@                      @      �?      $@      @      �?      @                                       @      @              2@                      �?      �?      @                      @      ,@      �?       @              �?       @              5@                      @              @      @      �?      �?     �F@      @      ,@      @      9@     �`@      @      c@      @      �?      @      5@      `@     @Y@      @     �L@     �E@      @      (@       @      3@     �\@      @     �[@      @      �?      @      5@     �Z@     @V@      @     �J@      B@      �?       @       @      ,@     @V@      @     �S@      @              @      3@     �W@      N@      �?     �C@      @      @      @              @      9@      �?      @@              �?               @      &@      =@       @      ,@       @               @       @      @      3@      �?     �E@                      @              7@      (@              @       @                       @              @      �?      &@                       @              .@      @                                       @              @      ,@              @@                      �?               @      "@              @     @Z@      @      $@      (@      A@     @w@      $@     H�@      *@       @     �F@     �A@     �{@     �p@      @     �[@     @Z@      @      $@      (@      A@     �v@      $@     (�@      *@       @     �F@     �A@     �{@     �p@      @     �[@     @Y@      @      $@      &@      @@      s@      $@     ��@       @      �?     �C@     �A@     px@     �o@      @     �X@      J@      @       @      @      3@     `e@      @     �v@       @      �?      9@      4@     pp@     �d@       @     �J@     �H@       @       @      @      *@     �`@      @     @m@                      ,@      .@      `@     �V@      @      G@      @      �?              �?       @     �K@             �\@      @      �?      @              K@      &@      �?      &@                                      �?      @              @                                       @      @              @      @      �?              �?      �?     �H@             @[@      @      �?      @              G@       @      �?      @                                              &@              @                                              @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��phG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�<�A�k�?�	           ��@       	                     @D�P�G?�?I           H�@                           @qk�r]��?           h�@                           @ЕrTC�?�           h�@������������������������       �p��$&{�?2           �}@������������������������       �B�0�~$�?q             f@                           �?�9�5��?m           h�@������������������������       �h��9��?�             j@������������������������       ��t_Ic��?�            �w@
                          �<@�	l���?9           �@                           �?��%-+�?           }@������������������������       �]�6��?�            �n@������������������������       �쬙1A�?�            �k@                          �>@p�����?            �C@������������������������       �窷uJ��?             3@������������������������       �p=
ףp�?             4@                          �;@�*x6��?o           �@                            @�7p%���?�           �@                            �?��_pVn�?f           T�@������������������������       �    \��?�            �@������������������������       ����Ȕ�?�            Pu@                           @*�����?c           `�@������������������������       ����'W�?�            �u@������������������������       ��\y^��?�            `j@                           @[{v��s�?�            �n@                          �=@�h��9�?�             j@������������������������       �&ޏ���?6             V@������������������������       �DDDDDD�?W             ^@                            �?K&:~��?             C@������������������������       ��8��8��?
             (@������������������������       �~e�.y0�?             :@�t�b�{     h�h4h7K ��h9��R�(KKKK��h��B�       �h@     �A@      A@      ;@     �Z@     p�@      =@     ȑ@      2@      ,@      S@      K@     �@     (�@      (@     �p@      [@      6@      :@       @     �P@     @q@      4@     �z@      *@      $@     �C@      ;@     �r@     `o@      @     @b@     �S@      *@      4@      @      I@     �h@      1@     pp@      (@       @      A@      6@     �k@     �e@      @     �]@      D@      &@      "@      @      6@     �^@      &@     �`@      �?              3@      @     �_@     �U@      �?     �N@     �@@      "@       @      @      1@      T@      @     �Y@      �?              2@      �?     @T@      O@      �?     �J@      @       @      �?       @      @     �E@      @      ?@                      �?       @      G@      8@               @     �C@       @      &@       @      <@     �R@      @      `@      &@       @      .@      3@     �W@     @V@      @     �L@      1@              @       @      @      1@       @     �C@      @      @      @       @      D@     �B@      @      5@      6@       @      @              6@     �L@      @     �V@      @      @      &@      &@      K@      J@       @      B@      =@      "@      @      �?      0@     �S@      @     `d@      �?       @      @      @      T@      S@      �?      <@      3@      "@      @      �?      ,@     @S@      @     `b@      �?       @      @      @     �S@      R@              :@      .@      @      @              @     �@@      �?     �U@      �?       @      @       @      B@      C@              .@      @      @      �?      �?      &@      F@       @      N@                       @      @      E@      A@              &@      $@                               @       @              0@                                       @      @      �?       @      @                               @       @              @                                      �?      @                      @                                                      $@                                      �?      �?      �?       @     �V@      *@       @      3@     �D@     �u@      "@     @�@      @      @     �B@      ;@      }@     �p@      @     @^@     �T@      $@       @      3@     �B@     s@       @     ؂@      @      @     �@@      9@      z@      o@      @     �[@     @Q@      @      @      .@      <@     �m@      @     0w@      @      @      ?@      2@     @q@      h@      @     �W@     �E@      @      @      ,@      0@     �g@      @      s@      �?              (@      ,@     `j@     �a@      @     �L@      :@              @      �?      (@     �H@      @     @P@       @      @      3@      @     @P@     �I@             �B@      ,@      @      �?      @      "@     �P@      �?      m@      �?               @      @     �a@      L@      �?      1@      @       @      �?      @      @      @@             `d@      �?               @      @     �U@      :@              (@       @      �?                       @      A@      �?     @Q@                              @      L@      >@      �?      @      @      @                      @     �D@      �?     @[@      �?      �?      @       @      G@      1@              $@      @      @                      @      A@      �?     @U@      �?      �?      @      �?     �D@      0@              $@      @      �?                      �?      &@              E@                       @              "@      ,@              @       @       @                      @      7@      �?     �E@      �?      �?       @      �?      @@       @              @                                              @              8@                              �?      @      �?                                                              �?              @                              �?       @      �?                                                              @              1@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ@ �=hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@�Ć 1k�?�	           ��@       	                     @~�-���?}           b�@                            �?�������?            ޣ@                           @���A���?�           ̝@������������������������       ���o?�?           Ȋ@������������������������       ��2���?�           h�@                           �?�� ����?�           ��@������������������������       �ɖd2 ��?             �I@������������������������       ��7٥��?h           H�@
                          �2@N��:d�?]           �@                           @������?�            0q@������������������������       ��
�?�            �m@������������������������       �O��E��?             B@                           �?��S�m�?�           x�@������������������������       ���(��?�            �r@������������������������       �G�a�?�            `x@                           @��,x��?           �y@                           @��[�v��?�            �v@                          �=@�X8�?�            0r@������������������������       �]�>�=�?U            �_@������������������������       �?B�� �?l            �d@                           @l(�����?.             S@������������������������       ���}�+�?             C@������������������������       ��k(����?             C@                           �?�/�K.��?            �D@������������������������       �      �?              @                           @�B��j��?            �@@������������������������       �      �?             0@������������������������       �@�0�!��?             1@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      7@     �E@      2@     �]@      �@      =@     ��@      4@       @     �O@     @P@     �@      �@      (@      o@     @e@      4@     �D@      2@      \@     ��@      =@     ��@      .@      @      N@      M@     Ȅ@     `�@      "@     �l@     @a@      ,@      >@      2@     �V@     �{@      6@     ��@      &@      @     �I@      F@     �|@      x@      "@     @h@     �X@      @      6@      0@     �L@     �u@      0@     �@      @      @      >@     �@@     0w@     pp@      @      _@      H@      �?      3@      @      ;@     �c@      @     �n@      @              0@      @     �f@      U@      @     �I@     �I@      @      @      "@      >@     �g@      (@     @p@      @      @      ,@      :@     �g@     `f@      @     @R@     �C@      "@       @       @     �@@     �W@      @     �^@      @      @      5@      &@     @V@     @^@       @     �Q@       @      �?      �?      �?              @              @      @              @               @      @       @      (@     �B@       @      @      �?     �@@     �V@      @     �]@      �?      @      1@      &@     @T@     �\@              M@      @@      @      &@              6@     @c@      @      t@      @      �?      "@      ,@     �i@     �a@             �B@      @               @              &@      D@      �?      U@                       @      @      T@     �B@              @      @               @              &@      B@              P@                              @      S@     �@@              @      �?                                      @      �?      4@                       @              @      @                      :@      @      "@              &@     �\@      @     �m@      @      �?      @      "@     @_@     �Y@              >@      0@      @      @               @      J@      @     �T@      @      �?      @      �?     �J@     �F@              .@      $@      �?      @              @      O@       @      c@      �?              �?       @      R@      M@              .@      5@      @       @              @     �R@             �e@      @      �?      @      @      Q@      8@      @      2@      5@      @       @              @     �Q@             �a@      @      �?      @      @     �O@      7@      @      2@      (@      @       @              @      L@             �Z@       @      �?      @      @      I@      6@      @      2@      @      @       @              �?      =@              B@                      @      @      5@      *@      �?      $@       @                              @      ;@             �Q@       @      �?              @      =@      "@       @       @      "@                                      .@             �A@      @                              *@      �?                      "@                                       @              7@      �?                              @                                                                      *@              (@       @                              $@      �?                                                              @              ?@                                      @      �?                                                              @               @                                       @                                                                                      =@                                      @      �?                                                                              .@                                              �?                                                                              ,@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJⳬ7hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @0l����?�	           ��@       	                    @���u'��?�           ��@                           @,�c0C��?.           �@                          �0@'�N!	�?�           ��@������������������������       ���T����?>             Y@������������������������       �.:��9��?�           h�@                          �>@��{�<�?L            �@������������������������       ��H4Ea.�?E           `@������������������������       �N��)x9�?             ,@
                          �7@Ę�s��?�            �@                           �?�3����?)           �}@������������������������       ��tF����?            �i@������������������������       ����M��?�            �p@                           �?�U�w�R�?�            �m@������������������������       �W?�`uV�?7            �W@������������������������       �|ZE��?U            �a@                           �?��d�?�           �@                          �;@w9��?�           p�@                           @2��eA�?k           x�@������������������������       �O�Z~�?Q           H�@������������������������       � ٞ u�?             C@                          �?@;�9c�?B            �W@������������������������       �`,�Œ_�?-             N@������������������������       ��NV�#�?            �A@                          �?@5�U�H��?#           P}@                          �0@w���E�?           �|@������������������������       ��h$��W�?	             .@������������������������       ���p�y�?           �{@������������������������       �.y0��k�?             *@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      ?@      G@      A@     �Z@     @�@      <@     ��@      1@      @     �O@     �D@     8�@     @      2@     �q@     @d@      9@     �B@      =@     �T@     @@      :@     ��@      (@      @      J@     �@@      @     @v@      0@     �l@     @`@      2@      <@      :@     @P@     �w@      (@     x�@       @      �?      B@      7@     0w@      m@      $@     �f@     �W@      2@      2@      4@      G@     �q@       @     w@      @             �@@      3@     Pq@     @g@       @     `b@      @      �?              @      @      =@               @                      �?      @      4@      &@              *@     �V@      1@      2@      0@      D@      p@       @     �v@      @              @@      0@     p@     �e@       @     �`@      B@              $@      @      3@     �W@      @     �c@      @      �?      @      @     �W@      G@       @      A@      >@              $@      @      3@     �W@      @     �c@      @      �?      @      @     @V@      G@       @      A@      @                                      �?               @                                      @                              @@      @      "@      @      2@     �]@      ,@      e@      @      @      0@      $@     @_@      _@      @      I@      ?@      @      "@              $@      U@      (@     �W@      @      @      *@      "@     �Q@     �T@      @      B@      7@      @      @               @     �D@      @      A@      �?      @      @      @      C@      8@      @      ,@       @      @      @               @     �E@      @     �N@      @              $@      @      @@     �M@       @      6@      �?                      @       @      A@       @     �R@                      @      �?     �K@     �D@              ,@                                      @      @             �B@                       @      �?      *@      6@              @      �?                      @      �?      ;@       @     �B@                      �?              E@      3@               @      F@      @      "@      @      7@     �f@       @     Px@      @              &@       @     pq@     �a@       @     �I@      =@      @      @       @      ,@     �Z@       @     `o@      @              @      @     @a@     @T@       @     �A@      4@      @      @       @      (@     @V@       @     �i@      @              @      @      `@     @S@             �@@      4@      @      @       @      &@     �U@       @     �f@      @              @      @     �^@     �Q@             �@@                                      �?      @              6@                                      @      @                      "@                               @      1@             �G@       @                              $@      @       @       @      @                              �?      *@             �@@                                       @      @       @              @                              �?      @              ,@       @                               @                       @      .@      @      @      @      "@     �R@             @a@                      @       @     �a@      N@              0@      .@      @      @      @      "@     @R@             �_@                      @       @     �a@      N@              0@                                              @               @                                              @                      .@      @      @      @      "@     @Q@             �]@                      @       @     �a@     �L@              0@                                              �?              &@                                      �?                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�W`hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?H�����?�	           ��@       	                     @�m.��@�?O           ��@                            �?�.�8���?           �@                           @Қc,���?           �y@������������������������       ��G��v�?�            @t@������������������������       �������?7             U@                          �4@�"oҶ��?           h�@������������������������       ��|'���?           �z@������������������������       �r�q{�?�             x@
                          �:@v����`�?4            ~@                           @�0��p�?�            `x@������������������������       ���p�a�?�            �v@������������������������       ��q��/��?             7@                           �?�Ԍ��	�?8            �V@������������������������       ���]�`��?             *@������������������������       ��Q<��8�?-            @S@                          �<@�����%�?|           H�@                            @�X�JF�?�           L�@                           �?������?�           �@������������������������       �u� ���??           �@������������������������       �,�b-���?N           (�@                           @H>�Ħ��?p           `�@������������������������       �[{+n���?           @{@������������������������       ���kN�?_             c@                            @"����3�?             j@                          �@@=��e@��?Y            �b@������������������������       ������?L            @`@������������������������       ���Q���?             4@                           @(�#|���?&            �M@������������������������       ������?             E@������������������������       �ҳ�wY;�?	             1@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@     �D@      E@      :@     �Y@     ��@     �A@     ��@      *@      @     �T@      Q@     ؆@     ��@      :@     �o@     �X@      7@      =@      *@     �P@     �r@      8@     z@      $@      @     �A@      B@     pq@     �l@      *@     �^@     �Q@      ,@      6@      *@      I@     �j@      0@     �q@       @      @      <@      A@      g@     �d@      $@     @Z@      4@      @      @      @      ,@      S@      @     �[@       @              @      .@     @R@      I@      @      6@      $@      @      @      @      "@     �K@      @     @X@       @              @      (@      K@      G@      �?      0@      $@                              @      5@              ,@                              @      3@      @       @      @     �I@      &@      3@      "@      B@      a@      &@     �e@      @      @      5@      3@      \@     �\@      @     �T@      =@      @      *@       @      4@     �R@      @     �V@      @      @      ,@      ,@      F@     @Q@      @      ?@      6@      @      @      @      0@     �O@      @     @T@      @      �?      @      @      Q@     �F@              J@      ;@      "@      @              0@     @V@       @     �`@       @              @       @     �W@     @P@      @      1@      1@      @      @              .@     @S@       @     �X@                      @      �?     �S@     �M@              1@      1@      @      @              *@     �Q@       @     @X@                      @      �?      S@      J@              .@                                       @      @               @                                      @      @               @      $@      @      �?              �?      (@             �A@       @                      �?      .@      @      @              @              �?                       @               @                                       @       @                      @      @                      �?      $@             �@@       @                      �?      *@      @      @              ]@      2@      *@      *@     �B@     �v@      &@     x�@      @       @      H@      @@     @|@     �r@      *@     ``@     @Z@      0@      *@      *@     �A@     �s@      $@     (�@       @       @     �G@      >@     0y@     pr@      *@     �^@     �U@      &@      $@      &@      ;@      n@       @     �v@      �?       @     �E@      8@     �p@     @j@      (@     @Y@      F@      �?      @      @      @     �W@      @     �`@                      $@      1@     �[@     �K@       @      ;@      E@      $@      @      @      5@     `b@      @     �l@      �?       @     �@@      @     `c@     `c@      $@     �R@      3@      @      @       @       @     �R@       @     `k@      �?              @      @      a@     @U@      �?      5@      .@      @      @       @      @      M@       @     �b@      �?              �?      @     @[@      O@      �?      1@      @      �?                      @      1@              Q@                      @      �?      <@      7@              @      &@       @                       @      I@      �?     �R@      �?              �?       @     �H@      @              "@      $@       @                              :@      �?      J@      �?              �?       @     �D@      @              @      $@       @                              2@      �?      H@      �?              �?       @     �B@      @              @                                               @              @                                      @      @              �?      �?                               @      8@              6@                                       @                       @      �?                               @      (@              3@                                      @                       @                                              (@              @                                       @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJt�"!hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @/�s
��?�	           ��@       	                     �?2�6M��?�           ��@                           @/:�٠�?F           .�@                          �<@������?j           ��@������������������������       ��cog���?7            �@������������������������       ������?3             U@                          �0@]	S|�?�           |�@������������������������       ��Ӟ�@�?1            �Q@������������������������       �0*���o�?�           d�@
                           �?��\��?�           ȅ@                           @,G7�?�            pt@������������������������       �%���4�?�            �r@������������������������       �����3��?             :@                          �;@�p��{��?�             w@������������������������       �*�	Hk��?�             u@������������������������       �     @�?             @@                           �?�@Z"�Z�?�           �@                           @V�O�;�?�           x�@                           @��9�?�           8�@������������������������       � ��Nm�?U            �@������������������������       ��3�Y��?E            �X@                          �5@�(\����?             D@������������������������       ����|���?             &@������������������������       ���`���?             =@                           @��OSFJ�?           �|@                          �1@,�'��?�            Ps@������������������������       �     ��?#             P@������������������������       �r��a �?�            �n@                           @C��g��?`            �b@������������������������       �?=j��?)            �Q@������������������������       ��$�^�4�?7            �S@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `j@      >@     �E@      A@      Y@     0�@      :@     h�@      0@      &@     �T@      M@     h�@     ��@      .@     q@     �b@      1@     �B@      =@     �U@     ~@      5@     (�@      .@      @     �Q@      J@     p~@     �x@      *@     �l@     @X@      *@      7@      9@     �K@     �v@      0@     ��@      $@             �B@      >@     px@     �q@       @     @d@     �K@      @      .@      (@      =@     @g@      @     �n@      @              1@      $@      g@     �X@       @      U@     �I@       @      &@      (@      ;@     �e@      @     @l@      @              ,@       @     �e@     �W@       @     �P@      @       @      @               @      (@      �?      5@                      @       @      (@      @              1@      E@      "@       @      *@      :@     �e@      &@     �s@      @              4@      4@     �i@      g@      @     �S@      @                                      @              *@                      �?      �?      3@      *@              "@     �A@      "@       @      *@      :@     �d@      &@     �r@      @              3@      3@     �g@     �e@      @     @Q@     �J@      @      ,@      @      ?@     @^@      @      ]@      @      @     �@@      6@      X@     �\@      @     �P@      7@      @      $@      @      3@      P@       @     �G@      @      @       @      (@     �F@     �H@      @      ?@      7@      @      "@      @      3@      O@       @     �A@      @      @       @      (@     �E@     �D@      @      >@                      �?                       @              (@                                       @       @              �?      >@      �?      @      �?      (@     �L@      @     @Q@       @       @      9@      $@     �I@     @P@       @      B@      <@      �?      @      �?      (@      K@      @      N@       @       @      9@      "@     �C@      P@              A@       @                                      @              "@                              �?      (@      �?       @       @     �N@      *@      @      @      ,@     �h@      @     Pw@      �?      @      *@      @     `p@     `a@       @      F@     �D@      �?      @      �?      $@     �\@       @      n@      �?      @      @       @     �`@     �V@       @     �@@     �D@      �?      @      �?      $@      Z@       @     �l@      �?      @      @       @      _@     @T@       @     �@@      ?@      �?      @      �?      @     �T@       @     �h@      �?       @      @       @      [@     �Q@              >@      $@                              @      6@              ?@               @                      0@      $@       @      @                                              &@              $@                                      $@      "@                                                                              @                                      @                                                                      &@              @                                      @      "@                      4@      (@              @      @     �T@      @     �`@                       @      @      `@     �H@              &@      0@      $@                       @     �I@       @     �S@                      @      @     �Y@      @@              @      @      @                              &@              1@                              @      "@      "@              @      "@      @                       @      D@       @      O@                      @      �?     @W@      7@              @      @       @              @       @      ?@      �?      K@                      @              :@      1@              @      @                      @       @      *@              5@                       @              &@      *@              �?               @                              2@      �?     �@@                       @              .@      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ<�^hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@��Uis��?�	           ��@       	                    �?-��A��?           �@                            �?�(\ �u�?T           ��@                          �5@�=����?m             f@������������������������       ������??            @[@������������������������       ��� =[�?.             Q@                          �0@m�� 6�?�            0v@������������������������       �b���i��?             &@������������������������       �b�ټ�?�            �u@
                           @A0��?+           �@                          �:@z;�3��?I           Ȕ@������������������������       �X�M���?+           ��@������������������������       �<pƵH�?             J@                           @�AH����?�           �@������������������������       ��Qval��?C           ��@������������������������       ��c���?�            @p@                           @�$���>�?           |@                           �?�.!���?�             y@                           @6������?0            �T@������������������������       �N�(�l\�?#            �L@������������������������       ��q�����?             9@                           @���Q �?�             t@������������������������       �����Q��?�            Pq@������������������������       �ҽ��?            �E@                            �?�Z�&�?            �G@������������������������       �     ��?	             0@                           �?�����?             ?@������������������������       ��$I�$I�?             @������������������������       �      �?             8@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      B@      <@      :@     �[@     ��@      @@     ��@      1@      @      W@     �P@     �@     ��@      5@      o@      g@      ?@      <@      9@     �X@     �@      ;@     ��@      ,@      @      T@     �N@     ��@     �@      2@      l@      B@      �?      @       @      0@     �P@      @      c@      �?              0@       @     @X@     @W@      @      B@      3@      �?                      @      >@      @     �G@                      @             �@@      7@              "@      1@      �?                              4@      �?      6@                      @              8@      *@              @       @                              @      $@       @      9@                      �?              "@      $@              @      1@              @       @      $@      B@      �?     �Z@      �?              $@       @      P@     �Q@      @      ;@       @               @              �?                                              �?                      @                      .@              @       @      "@      B@      �?     �Z@      �?              "@       @      P@     @P@      @      ;@     �b@      >@      7@      7@     �T@      �@      7@     ��@      *@      @      P@     �M@     ��@     �y@      ,@     �g@     @V@      $@      ,@      .@      D@     p@      $@     @u@      "@      �?      :@      0@     �p@     `c@      @     �R@     �U@      $@      ,@      *@      B@     �o@      $@     �t@      "@      �?      :@      0@     �n@     `b@      @     �R@      @                       @      @      @              @                                      6@       @              �?      N@      4@      "@       @     �E@     �q@      *@     �z@      @      @      C@     �E@     �p@     p@      @     �\@      H@      1@       @       @      ;@     @o@      $@     �u@      @      @      ?@      B@     �l@     �l@      @     @V@      (@      @      �?              0@     �B@      @     �T@              �?      @      @      B@      <@      �?      9@      4@      @              �?      &@      T@      @     �d@      @              (@      @     @S@     �B@      @      7@      4@      @              �?      &@     �R@      @     �a@      @              &@      @      O@     �B@      @      7@      @      @                              (@              5@                      �?      @      &@      1@              @      @      @                              (@              "@                      �?      @      &@      @              @                                                              (@                                              *@                      .@       @              �?      &@      O@      @      ^@      @              $@      �?     �I@      4@      @      0@      (@       @              �?      &@     �G@      @     �[@      @              $@      �?      D@      .@      @      0@      @                                      .@              "@                                      &@      @                                                              @              9@                      �?              .@                                                                                       @                      �?              @                                                                      @              1@                                       @                                                                       @              @                                      �?                                                                      @              *@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJF�;hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @<���=q�?�	           ��@       	                     �?����4��?            �@                           @J|�\���?�           ��@                           @��<��?�           ��@������������������������       �^�G�0��?�           �@������������������������       �(������?             9@                           @P$+�_T�?�            �p@������������������������       ����zAp�?l            �e@������������������������       �I�O���?;             W@
                          �;@�f��m�?^           ,�@                           @Ԓ��ir�?�           x�@������������������������       ��p�˂�?�           ��@������������������������       �9��YN�?p           @�@                           �?�� �?��?j            �e@������������������������       ���~UZ��?+            @Q@������������������������       �C�����??             Z@                           �?�ه�7��?�           `�@                           �?��� ��?�            �@                           @�m��?r            �f@������������������������       �=�]���?X            �a@������������������������       �3�R�f�?             C@                          �6@�u�m�q�?&            }@������������������������       ��b����?�            `n@������������������������       ���]���?�            �k@                           @c򗛀{�?"           @}@                          �1@��H���?�            �l@������������������������       ���ͽ1��?            �B@������������������������       �l`2^v9�?v             h@                          �4@e��>��?�            �m@������������������������       ��q�q�?Q            �`@������������������������       ����s�?C            �Z@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@      :@      G@      <@     @\@     P�@      @@     ��@      1@      @     @Q@      R@     ��@     0�@      4@     �j@     `e@      6@      A@      :@      W@     �~@      <@     @�@      (@       @     �M@     �L@     @     �x@      1@      g@      M@      "@       @      $@      6@      h@      $@     @u@       @              0@      .@     �f@      b@      @     �F@     �H@      �?      @      @      3@     �c@      @     �p@       @              $@      ,@     `a@     @V@      @      >@     �H@      �?      @      @      0@     `c@      @     `o@       @              $@      *@      a@     �U@      @      =@                                      @      @              *@                              �?       @       @              �?      "@       @      @      @      @     �A@      @      S@                      @      �?      F@      L@      �?      .@      @      @      �?      @              =@      @      K@                      @              4@      F@      �?      @      @       @      @      �?      @      @      �?      6@                      @      �?      8@      (@              $@     @\@      *@      :@      0@     �Q@     �r@      2@     @w@      $@       @     �E@      E@     �s@      o@      &@     `a@     @W@      @      8@      ,@     @Q@     pq@      2@     `t@      $@       @      B@     �C@      q@     @m@      "@     �`@     �E@      @       @      $@      0@      Y@      @     �Y@      @              3@      .@     �^@     �W@      �?      L@      I@      @      0@      @     �J@     `f@      ,@      l@      @       @      1@      8@      c@     �a@       @      S@      4@      @       @       @      �?      7@              G@                      @      @      D@      ,@       @      @      ,@      @       @              �?       @              &@                      @              0@      &@              @      @       @               @              5@             �A@                       @      @      8@      @       @      @     �D@      @      (@       @      5@     `g@      @     �y@      @      �?      $@      .@     �m@     @_@      @      ?@      :@      �?      "@      �?      *@     @Y@      �?     @o@      @      �?      @      *@     �\@     �T@      @      3@      @              @              @      =@             �M@                      �?       @      E@      =@              @      @              @              @      3@              I@                      �?       @     �B@      .@              @                                              $@              "@                                      @      ,@                      6@      �?      @      �?      "@      R@      �?     �g@      @      �?       @      &@     @R@      K@      @      *@      @               @      �?      @      G@      �?      Y@       @      �?      �?      @     �@@      C@              @      0@      �?      @              @      :@             �V@      @              �?       @      D@      0@      @      @      .@      @      @      �?       @     �U@      @     �d@                      @       @     �^@      E@              (@       @       @      �?              @      D@       @     �R@                              �?     �R@      3@              @      @                                       @              $@                                      @      @              @      @       @      �?              @      @@       @     @P@                              �?     @Q@      *@              �?      @      �?       @      �?      @      G@      �?     @V@                      @      �?     �G@      7@               @      @                      �?      @      =@      �?      J@                      @              2@      (@              @       @      �?       @               @      1@             �B@                              �?      =@      &@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJA��&hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�#Nօ��?�	           ��@       	                     @~'�'`T�?G           ��@                          �1@���(��?            �@                           @���[�?�            �m@������������������������       �%����$�?k             c@������������������������       �E~����?4            �U@                           �?�q/x�_�?z           D�@������������������������       ��L��d�?�            @p@������������������������       ���R�e�?�           h�@
                          �:@V��[�Z�?.           �~@                          �7@�fCMji�?           �y@������������������������       �B� ����?�            Pt@������������������������       �/'��?3            �U@                          �=@d[�Ƃg�?+            �S@������������������������       ���!O|��?            �I@������������������������       ��P���?             ;@                            @��&���?C           ��@                           @���K:|�?�           8�@                            �?�pP�q�?�           ��@������������������������       �s^|���?�            �p@������������������������       �vrWQ�?�            y@                          �7@9�`1\V�?(           x�@������������������������       �Șu�U��?�           p�@������������������������       �2��)�?�            p@                           @�M@�A�?o           ��@                           @1�?��?           �|@������������������������       �5)U[�?�            @v@������������������������       ���u���?B             Y@                           @dp��w�?P            @a@������������������������       �i#[�G��?1             U@������������������������       �ȟa����?             K@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        j@      B@      A@      1@     �[@     h�@     �D@     X�@      .@      @     �T@     �Q@     ��@     ��@      .@     `p@     �]@      1@      <@       @     �R@     `r@      <@     0z@       @      @      F@     �C@     0r@     Pp@      @     @`@     �W@      0@      4@       @      O@     `i@      9@     0r@       @      @      @@      =@     @g@     �g@      @     �Z@      2@      @      @              (@     �D@      $@      ?@      @      �?      @       @      9@     �H@       @      :@      ,@      @       @              $@      ;@      @      2@      �?      �?       @      @      5@      7@      �?      5@      @               @               @      ,@      @      *@      @              @      @      @      :@      �?      @     @S@      *@      0@       @      I@     @d@      .@     @p@      @      @      ;@      5@      d@     �a@       @      T@      1@      @      @      �?      3@      I@             �Q@                      @      @      ?@      9@              <@      N@      @      *@      @      ?@      \@      .@     �g@      @      @      5@      1@     @`@     @]@       @      J@      7@      �?       @              *@     �V@      @      `@              �?      (@      $@     @Z@     �Q@              8@      2@      �?      @              (@     �S@      @     @Y@              �?      (@      @      V@     @P@              4@      ,@      �?      @              &@     �J@      @     @U@              �?       @      @     @P@      K@              3@      @                              �?      :@              0@                      @              7@      &@              �?      @              @              �?      (@              ;@                              @      1@      @              @      �?              @                       @              7@                                      (@       @              �?      @                              �?      @              @                              @      @      @              @     �V@      3@      @      "@      B@     pt@      *@     ��@      @       @      C@      @@     �z@     �r@      &@     �`@     �Q@      0@      @      "@      @@     Pp@      (@     �z@      @      �?      B@      :@     �r@     �k@      &@      ]@      >@      (@      �?      @      ,@      ]@      @     �e@       @              3@      (@      d@     �Q@       @      G@      *@      @              @      @     �N@      @     �U@                                      O@      8@      �?      @      1@       @      �?      @      "@     �K@       @     �U@       @              3@      (@     �X@      G@      �?      D@      D@      @       @       @      2@      b@      @      p@      @      �?      1@      ,@     �a@      c@      "@     �Q@      A@      @       @       @      *@      \@      @     `d@      �?              &@      (@     �V@     �\@      @      I@      @                              @     �@@             @W@       @      �?      @       @      I@     �B@       @      4@      5@      @      @              @     �P@      �?     `p@       @      �?       @      @      `@     �S@              0@      0@      @      @              @      I@      �?     �f@       @      �?       @      @     �Y@     @Q@              .@      *@       @      @              @      ?@      �?     �c@       @      �?       @      @      T@     �E@              (@      @      �?                              3@              9@                              �?      6@      :@              @      @                                      0@              T@                                      :@      $@              �?      �?                                       @             �J@                                      0@      @                      @                                       @              ;@                                      $@      @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��ZhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @
GaZu�?�	           ��@       	                    �?$��7��?�           R�@                            �?*w�d(P�?           ��@                          �=@x�|���?f           X�@������������������������       ������?H           ��@������������������������       �����?            �J@                          �4@������?�            Pq@������������������������       �����G��?b             d@������������������������       �(�����?M             ]@
                           @$���^u�?�           $�@                           �?"�Nc�?�           ��@������������������������       �e��9D��?�            @p@������������������������       ��5bi�B�?B           (�@                          �;@m��1GI�?            z@������������������������       ��*$�X��?�            �w@������������������������       �$�ɜoB�?             A@                           @&ޏ���?�           ��@                           �?�EW�R��?�            �@                           @���K��?5           �|@������������������������       �t[�T]0�?�            �v@������������������������       ��q�q��?@             X@                           �?Ԋ���?|           ȁ@������������������������       ��4����?D            �Y@������������������������       � ZRH���?8            }@                           !@��8��8�?             8@������������������������       �T�r
^N�?             ,@������������������������       ���Q��?             $@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      <@      C@      &@      _@     `�@      F@     ��@      0@      "@      S@      Q@     ��@     �@      3@      n@     �c@      3@      <@      "@     �X@     �}@     �@@      �@      (@      @     �P@     �M@     Ѐ@      y@      0@      i@     �R@      "@      2@      @      L@     �k@      2@     �q@      @      @      6@      B@     `j@     �e@      @      Z@      N@      @      .@       @     �F@     �g@      (@     �l@       @       @      2@      6@     �e@     @_@      @     �Q@     �M@      @      .@       @     �B@     `g@      (@     �i@       @       @      2@      6@      e@      \@      @     @Q@      �?                               @      @              7@                                      @      *@              �?      ,@      @      @       @      &@     �@@      @     �L@      �?      �?      @      ,@     �C@      I@      @      A@      @      @               @      @      6@      @      7@              �?      @      $@      2@     �@@      @      :@      &@      �?      @              @      &@      �?      A@      �?                      @      5@      1@               @     �T@      $@      $@      @      E@     @o@      .@     p|@      "@      @     �F@      7@     pt@      l@      "@     @X@     �Q@      @      @       @      :@     �g@      *@     �s@      @      @      <@      0@     �p@     `f@      @     �K@      3@      @      @               @      =@             �N@                      @      �?     �O@      F@      �?      5@     �I@      @      @       @      2@      d@      *@     p@      @      @      5@      .@     `i@     �`@      @      A@      *@      @      @      @      0@     �N@       @      a@       @              1@      @     �N@      G@       @      E@      *@      @      @       @      0@      K@       @     @^@       @              1@      @      J@      G@       @      E@                              �?              @              0@                              �?      "@                             �C@      "@      $@       @      :@     `f@      &@     x@      @       @      "@      "@     �k@     �Z@      @     �C@     �C@      "@      $@       @      :@     �e@      &@     �w@      @       @      "@      "@     �j@     @Z@      @      C@      :@      @      @      �?      0@      R@      @     @c@      �?       @       @      @     �U@     �K@      @      0@      3@      @      @      �?      ,@     @P@      @      \@      �?              @      �?     @Q@     �F@      @      ,@      @       @                       @      @      �?      E@               @      �?       @      2@      $@               @      *@       @      @      �?      $@     @Y@      @      l@      @              �?      @     �_@      I@              6@      @               @              @      &@      @     �B@                                      1@      0@              @      @       @      �?      �?      @     �V@      @     �g@      @              �?      @     @[@      A@              1@                                              @              @                                      "@       @              �?                                               @               @                                      "@      �?                                                              @              @                                              �?              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ1�i)hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @�׭;q�?�	           ��@       	                    �? hIU��?�           �@                           �?��u5�p�?           ��@                          �8@�����?_            @c@������������������������       ����*���?L            �^@������������������������       �     ��?             @@                          �1@O���s�?�           H�@������������������������       ���m���?�            @j@������������������������       �����;�?1            �@
                          �;@_˾uU�?�           h�@                           @8X�)��?f           |�@������������������������       �Z'&!��?U           ��@������������������������       �<Cb�ΐ�?            �@@                           @���~y�?u            `g@������������������������       �@��,*�?M            �]@������������������������       ��������?(             Q@                           �?�k���?�           �@                           �?�k	2B�?(           0|@                           @��s����?6            �R@������������������������       �,�wɃ�?'             J@������������������������       �ֳC��2�?             6@                           @p]K�E�?�            �w@������������������������       ��	��w�?            �g@������������������������       ��t�'�?s            `g@                          @@@R����?�            �@                           @���G���?�           (�@������������������������       ��¶�*�?*           �|@������������������������       ��4�gV�?g            `c@������������������������       ���B�f�?             ;@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `i@      4@      H@      8@     �[@     p�@      :@     ��@      1@      @     @R@     �Q@     ��@     (�@      1@      o@     �d@      ,@      ?@      3@     �U@     �}@      6@     І@      .@      @      Q@     �L@     �@     �x@      .@      j@     �U@      @      9@       @     �K@     @k@      @      q@      $@      @      7@      =@     �i@     `g@       @      ]@      "@              @               @      6@              B@      �?               @       @     �B@      ,@              ,@      "@              @              @      .@              @@      �?              @       @      8@      ,@              ,@                                      @      @              @                      @              *@                             @S@      @      6@       @     �G@     �h@      @     �m@      "@      @      .@      ;@      e@     �e@       @     �Y@      *@              @      �?      *@     �B@      @      9@      �?      �?      �?      &@      ?@     �E@      @      3@      P@      @      .@      @      A@     �c@       @     �j@       @      @      ,@      0@     @a@     @`@      @     �T@     @T@       @      @      &@      ?@     �o@      1@     �|@      @             �F@      <@     Ps@     `j@      @     @W@     �S@      @      @      $@      ?@      k@      .@     �w@      @              E@      :@     �p@     �h@      @     @U@      R@      @      @      $@      >@      j@      .@     �w@      @              E@      :@     0p@     `h@      @      U@      @                              �?       @              �?                                      &@      @              �?       @      @              �?              C@       @     �R@                      @       @     �C@      (@      @       @       @      @              �?             �@@       @     �@@                      �?      �?      ;@      @      @       @                                              @             �D@                       @      �?      (@      @                      B@      @      1@      @      8@     �f@      @     �x@       @      �?      @      *@     @n@     �]@       @      D@      8@       @      (@       @      2@     �R@       @     ``@      �?      �?      @      @     �W@      M@      �?      4@      @               @              @      (@              .@                      �?              ,@      0@              @      @               @              @      $@              @                      �?              "@      (@              @      @                                       @               @                                      @      @                      2@       @      $@       @      .@     �O@       @      ]@      �?      �?      @      @      T@      E@      �?      .@      @      �?      "@       @      @      5@      �?      O@      �?              @      �?      H@      8@              @      &@      �?      �?               @      E@      �?      K@              �?              @      @@      2@      �?      (@      (@      @      @      @      @     �Z@       @     `p@      �?              �?      @     �b@     �N@      �?      4@      (@      @      @      @      @     �Z@       @     �o@      �?              �?      @     �`@     �N@      �?      4@      &@       @      @      @       @      M@       @     `i@      �?              �?      @      Z@      G@              ,@      �?       @                      �?      H@              I@                              �?      >@      .@      �?      @                                      @      �?              "@                                      ,@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��LhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?��Al�?�	           ��@       	                   �1@��	�J�?R           �@                           @Ћ�Կ��?�            �s@                           @$�Y��v�?h            �c@������������������������       � ^�/��?Q            @_@������������������������       �F��'s��?             A@                          �0@{J��b,�?d            @c@������������������������       ��2�o�U�?%            �K@������������������������       ��u=WTK�??            �X@
                           @�$�4��?�           �@                           �?Dk{7B��?�           �@������������������������       ��Ęfb��?L           �@������������������������       �$Z���z�?i           P�@                            �?     ��?�             t@������������������������       �������?v            �f@������������������������       �)-��21�?[             a@                            @�O����?k           �@                            �?�^���<�?�           ��@                           @0	��@��?�           Ȓ@������������������������       �(.�JC��?�           (�@������������������������       ��8�i�?C           h�@                          �>@�}�%�W�?�            pw@������������������������       �V'�p�u�?�            �v@������������������������       ��θ�?             *@                          �2@�PBP%�?�            �@                           @��|D\�?f            `d@������������������������       �)�a��?I            @\@������������������������       ���=yX��?             I@                           @�F407��?$           |@������������������������       �����u�?           py@������������������������       �&�to@��?             E@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        f@     �A@      C@      9@     �Z@     X�@      =@     T�@      7@      "@     �Q@      M@     �@     �@      1@     �o@      T@      5@      >@       @     �Q@     ps@      0@     �x@      *@      @     �@@      =@     pu@     �k@      @     �a@      0@      @      .@              4@     �H@       @     �G@      @       @       @      @     �P@      C@       @      <@      @      @      @              @      A@      @      6@       @               @      @      A@      2@              1@      @      @      @              @      7@       @      ,@                       @      @     �@@      .@              1@      @              �?              �?      &@      @       @       @                              �?      @                      "@      �?       @              .@      .@      @      9@      �?       @      @      @      @@      4@       @      &@       @      �?      @               @       @      @      $@      �?              �?              ,@      @              @      @              @              @      *@              .@               @      @      @      2@      ,@       @      @      P@      1@      .@       @     �I@     `p@       @     �u@      $@      @      9@      6@     Pq@     �f@      @     @\@      M@      .@      *@       @      F@     �g@       @     �q@       @      �?      6@      3@     �k@     �`@      @     �Q@      ?@       @      @      @      3@      U@       @      _@      �?              (@      &@      W@     �S@             �C@      ;@      *@       @      @      9@     �Z@              d@      @      �?      $@       @      `@     �K@      @      ?@      @       @       @              @     �Q@      @     �P@       @       @      @      @     �L@      I@             �E@      @      �?                      @      C@      @      6@                      @       @      B@      <@             �C@      @      �?       @               @     �@@              F@       @       @              �?      5@      6@              @      X@      ,@       @      1@      B@     @w@      *@     @�@      $@      @     �B@      =@     �z@     r@      (@     �\@      R@      "@      @      *@      =@     �p@      *@     @}@      @      @     �A@      :@     �r@      l@      &@     �W@     �I@      @      @      &@      3@     �j@      "@     0x@      @              1@      1@     `m@      c@       @     @P@      A@      @      @       @      $@     �`@      @      j@      @               @      @      _@     �T@      @     �F@      1@      @              "@      "@      T@      @     `f@      �?              "@      $@     �[@     �Q@      @      4@      5@       @      @       @      $@     �L@      @     @T@              @      2@      "@     �N@     �Q@      @      >@      5@       @      @       @      $@     �L@      @     �Q@              @      2@      "@      M@     �Q@      @      >@                                                              $@                                      @                              8@      @      �?      @      @     @Y@             �n@      @      �?       @      @     @`@     @P@      �?      3@      "@              �?      @       @      9@             �I@                      �?             �J@      ,@              @      @              �?      @       @      .@              <@                                      D@      ,@              @      @                                      $@              7@                      �?              *@                              .@      @              �?      @      S@              h@      @      �?      �?      @     @S@     �I@      �?      .@      *@      @              �?      @     �O@             `f@      �?      �?      �?      @     �R@      H@      �?      ,@       @       @                              *@              ,@      @                              @      @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�tb>hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@��yX_�?�	           ��@       	                   �0@�N�ފ�?�           ��@                           �?��H.��?�             i@                           �?�ks����?            �F@������������������������       ���8��8�?             8@������������������������       �VUUUUU�?             5@                            �?ֵ�����?j            `c@������������������������       �:|z3�?             E@������������������������       �'7a��t�?O            @\@
                           @ڔ�̙x�?           d�@                            @h[�A�?�           d�@������������������������       ����%��?�           ��@������������������������       �5��1C�?           �{@                            @��󿦙�?V           d�@������������������������       ��c�q�?           ��@������������������������       ���xb��?=           P@                           @	m� �b�?"           �|@                           �?�:�S���?            z@                            @�s>1���?m            �e@������������������������       �I�N�V��?G            @]@������������������������       �YM�#:�?&             M@                            @��F[���?�            `n@������������������������       �k��5���?d            �d@������������������������       �̹�m���?2             S@                           �?���zm��?            �F@������������������������       �>;n,��?	             &@                          �=@����p�?             A@������������������������       �d��b��?             5@������������������������       ��n_Y�K�?             *@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      >@     �E@      :@     �U@      �@      @@     Б@      5@       @     �R@      M@     (�@     �@      7@      o@     �e@      <@      E@      9@     @T@     h�@      ?@     ��@      .@      @     �O@      J@     ��@     P~@      5@     �k@      @      �?              @      @     �A@      �?      B@      �?              @      @     �@@     �F@      �?      6@                                       @      &@              �?                                      (@      $@              "@                                       @       @                                                      @      $@              @                                              "@              �?                                      @                      @      @      �?              @      @      8@      �?     �A@      �?              @      @      5@     �A@      �?      *@                              �?       @      @              .@                       @              @      (@                      @      �?               @      �?      4@      �?      4@      �?              @      @      .@      7@      �?      *@      e@      ;@      E@      6@      S@     P�@      >@     ��@      ,@      @      M@      G@     ��@     �{@      4@      i@     @U@       @      =@      *@      @@     �m@      @     �{@      @      @      4@      6@     @t@     �d@      $@     @Y@     �P@      @      3@      $@      <@     @f@      @     r@      @      @      &@      4@     `j@     �]@      $@     �S@      3@       @      $@      @      @      M@             �b@                      "@       @     @\@     �G@              6@      U@      3@      *@      "@      F@     �q@      9@     �}@      &@      @      C@      8@     u@      q@      $@      Y@     @P@      (@      "@       @      ?@     @j@      6@     �r@      "@      @     �@@      4@     �j@     �k@      "@     �U@      3@      @      @      �?      *@      S@      @      f@       @      �?      @      @     �^@     �J@      �?      ,@      5@       @      �?      �?      @     �T@      �?     �g@      @      �?      (@      @     �S@      =@       @      9@      5@       @      �?      �?      @     �S@      �?     @d@      @      �?      $@      @     �Q@      =@       @      8@      .@      �?      �?               @      8@             �O@       @              @      @      :@      0@      �?      ,@      @      �?      �?              �?      1@              E@                      @              1@      ,@              *@      &@                              �?      @              5@       @                      @      "@       @      �?      �?      @      �?              �?      @      K@      �?     �X@      @      �?      @      �?     �F@      *@      �?      $@      @      �?              �?      �?      C@      �?      L@       @              @      �?      B@      (@      �?      "@      �?                               @      0@             �E@       @      �?                      "@      �?              �?                                              @              ;@                       @       @       @                      �?                                                              @                                      @                      �?                                              @              6@                       @       @      @                                                                      @              *@                       @              �?                                                                                      "@                               @       @                        �t�bub��      hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�iHhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?�~�̙�?�	           ��@       	                     @M #�+�?Y           t�@                            �?��`>���?0           8�@                          �2@��		A�?m           ��@������������������������       ��<����?�            �r@������������������������       ���t���?�           P�@                           @�.�|J�?�            �s@������������������������       ����#'�?�            �q@������������������������       ���S����?             ;@
                           @J�{t���?)           �|@                           �?J��3#�?�            `v@������������������������       �����?�            �p@������������������������       ��0����?;            @V@                          �;@\���'�?H            @Z@������������������������       �������??            �V@������������������������       �      �?	             ,@                           �?}�W���?c           ؠ@                          @@@�tϻ���?w           Ђ@                          �<@d��|��?p           P�@������������������������       �g�?;���?^           h�@������������������������       �΃�\�?             =@������������������������       �     @�?             0@                          �6@��)z+�?�           H�@                            @�K�R
��?c           @�@������������������������       �&�����?�           `�@������������������������       �8����R�?�            �o@                           @S@�����?�           P�@������������������������       ���X.L�?�            Pv@������������������������       �^��zg�?�            Pp@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        g@      =@     �B@      =@     �\@     H�@     �J@     L�@      8@      &@     �W@      L@     ��@     �~@      ?@     �n@     @V@      5@      9@      $@     �Q@     Ps@      9@     �{@      1@      @      I@      <@     �r@     �l@      "@      `@     @Q@      2@      4@       @      J@      l@      2@     �q@      *@      @      D@      9@      k@      f@      "@     �\@      M@      ,@      1@      @      >@      f@      *@     `m@      @       @      ;@      ,@     `d@     �_@       @     @U@      4@              @      �?      &@     �F@      @      J@      �?       @      @      @     �F@      N@      @      ;@      C@      ,@      $@      @      3@     �`@      @     �f@      @              4@      @     �]@     �P@       @      M@      &@      @      @      @      6@      H@      @     �I@       @      @      *@      &@     �J@     �H@      �?      =@      &@      @      �?      @      6@     �G@      @      E@      @      @      *@      &@     �H@      E@      �?      <@                       @                      �?              "@      @                              @      @              �?      4@      @      @       @      3@      U@      @     @c@      @      �?      $@      @     �T@      K@              .@      3@       @      @              0@     @P@      @      \@      @      �?      @      @      N@     �G@              *@      ,@              @              "@      F@      @      W@      @      �?      @       @     �F@      B@              "@      @       @                      @      5@      @      4@                              �?      .@      &@              @      �?      �?               @      @      3@      �?      E@                      @              6@      @               @      �?      �?               @       @      3@      �?     �@@                      @              2@      @               @                                      �?                      "@                                      @                             �W@       @      (@      3@     �E@     @w@      <@     ؄@      @      @     �F@      <@     �z@     `p@      6@      ]@      >@      �?      @      @      0@     �\@       @     �d@      �?              $@      *@     �b@      P@      @      7@      >@      �?      @      @      (@     �\@       @     �c@                      $@      *@     �b@      P@      @      7@      =@              @      @      (@     @Y@       @      c@                      $@      (@     �a@      O@      @      6@      �?      �?                              *@              @                              �?      @       @              �?                                      @                      $@      �?                              �?                             @P@      @       @      .@      ;@      p@      :@     @@      @      @     �A@      .@     `q@     �h@      2@     @W@     �G@      @      @      ,@      0@     @c@      (@     �p@      @      @      8@       @      c@     `a@      &@     @Q@     �@@      @      @      (@      &@     �Y@      @     �f@      �?      @      8@      @      \@     �\@      &@      M@      ,@      �?      @       @      @      J@      @     @V@       @                       @      D@      9@              &@      2@       @      �?      �?      &@      Z@      ,@     �l@      @      �?      &@      @     �_@     �M@      @      8@      (@       @      �?              @     �K@      (@     �b@      �?              @      @     �P@      5@       @      5@      @                      �?      @     �H@       @     @T@       @      �?      @      @     �M@      C@      @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ
�nhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @"=i݆��?�	           ��@       	                    �?W�;���?�           ��@                          �1@�[���?           H�@                          �0@    �3�?�             p@������������������������       �     @�?>             X@������������������������       ������<�?c             d@                           �?!�5KE�?p           ��@������������������������       �$i��6�?K            @]@������������������������       ���wOf�?%           �@
                           !@�	�� ��?�           ��@                            �? �����?�           |�@������������������������       � �Ke��?�           Ē@������������������������       �*D;���?�            �v@������������������������       �p=
ףp�?             $@                          �2@�YZ�&�?�           8�@                           @�,��n*�?�             q@                           �?¯	���?s            �e@������������������������       �ʵ�:"�?            �E@������������������������       ��=z�x�?U            �`@                          �0@��(�^�?>            �X@������������������������       �0\�Uo��?
             3@������������������������       ��Q��k�?4             T@                          �6@��?�K�?           ��@                           �?7�"��?�            �x@������������������������       �4�f�̞�?+            �Q@������������������������       �ʚ0D�?�            0t@                           @4v2�� �?            {@������������������������       ��NC���?h            `e@������������������������       �p�G��?�            pp@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @j@      C@      D@      4@     @[@     8�@      F@      �@      *@      @     �U@      P@     X�@     �@      ;@     �p@     �d@      7@      ?@      ,@     �T@     0}@     �@@     ��@      "@      @      S@     �M@     �@     @x@      7@     �l@     @T@      (@      8@      "@      F@      k@      0@     �p@      @       @      A@      :@      h@     `e@      (@     �^@      2@       @      @              $@      C@       @      ?@      �?      �?      @      $@      B@      E@      @      D@      @       @       @              @      &@      @      (@      �?                      �?      1@      9@       @      &@      .@              @              @      ;@      @      3@              �?      @      "@      3@      1@      @      =@     �O@      $@      2@      "@      A@     @f@       @     @m@      @      �?      ;@      0@     �c@      `@      @     �T@      @      @      �?              @      2@             �E@      �?              @      �?      8@      @              @     �M@      @      1@      "@      ?@      d@       @     �g@      @      �?      4@      .@     �`@     �^@      @     �S@      U@      &@      @      @      C@     `o@      1@     �z@      @       @      E@     �@@     t@      k@      &@     @Z@      U@      &@      @      @      C@     �n@      1@     �z@      @       @      E@     �@@     �s@      k@      &@     @Z@      M@      $@      �?      @      5@      h@      0@      w@      @              9@      (@     0p@      c@      @     �R@      :@      �?      @      �?      1@     �I@      �?      O@               @      1@      5@      N@     �O@      @      ?@                                              @                                                       @      �?                     �F@      .@      "@      @      ;@     �f@      &@     �x@      @       @      $@      @      m@     @]@      @     �D@       @                      @      "@      G@       @     �T@                      @      @     �S@      9@              &@      @                       @      "@      A@              G@                      �?      @      F@      5@              $@      �?                              @      "@              *@                      �?      �?      @      @              @      @                       @      @      9@             �@@                              @      C@      2@              @      @                      @              (@       @     �B@                       @              A@      @              �?                                              @       @      $@                                      �?       @                      @                      @               @              ;@                       @             �@@       @              �?     �B@      .@      "@      �?      2@     �`@      "@     `s@      @       @      @      �?     `c@      W@      @      >@      3@      @      @      �?      "@      M@       @      d@      �?              @             �I@      I@              7@      "@              �?                      0@      �?      5@                                       @      &@              $@      $@      @      @      �?      "@      E@      @     �a@      �?              @             �H@     �C@              *@      2@      &@      @              "@      S@      �?     �b@      @       @      @      �?      Z@      E@      @      @      @              @              @      3@              N@               @      @      �?     �E@      9@              @      &@      &@      �?              @     �L@      �?     @V@      @                             �N@      1@      @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ3��IhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @4��k�?�	           ��@       	                    @�IN,��?�           ��@                            �?ևn���?8           ��@                           �?���{���?<           ��@������������������������       ����y_��?�            0y@������������������������       �#�k�*��?E           �@                           �?�A>�S_�?�           ܘ@������������������������       ���@ mx�?           �{@������������������������       ��c�/D�?�           ��@
                           �?@e���?�            �o@                           �?\��"e��?4            �V@������������������������       ��"�O�|�?	             1@������������������������       ��i�%ʐ�?+            @R@                           @�]�ڕ��?e            �d@������������������������       �8h����?K            �^@������������������������       �҉�&S��?            �D@                           �?��ȴ�?�           �@                          �:@T{'fyP�??           P�@                           @�;s�f`�?           @{@������������������������       ����~jV�?�            �y@������������������������       �������?             <@                           @s�k����?0            �U@������������������������       ��u�f�?&             Q@������������������������       �B{	�%��?
             2@                           @/���?�           ��@                          �;@W��Y��?-           �|@������������������������       ����!��?           0y@������������������������       ��xp�dk�?"            �K@                          �2@9��8���?l            �e@������������������������       ��c�Α�?             =@������������������������       ���a���?\             b@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      A@     �C@      *@     @[@     Ȅ@      ;@     l�@      *@       @     �P@      O@     ��@     ��@      ,@     �o@     @c@      8@      A@      "@      V@     �~@      6@     @�@      $@      @      N@      I@      @      x@      &@     �i@      b@      6@      =@      "@      T@     �|@      5@     ��@      "@      @     �H@     �G@     �|@     �u@      &@     @g@     �E@      "@      @      @      2@      g@      @     �q@      @              "@      &@     `e@      ]@      �?     �I@      3@      @      @               @     �Q@      @      a@                      @      @     �P@     �I@              A@      8@      @      @      @      $@     @\@       @     @b@      @              @       @     @Z@     @P@      �?      1@     @Y@      *@      7@      @      O@      q@      0@     `u@      @      @      D@      B@      r@     @m@      $@     �`@      =@      @      @      �?      *@     �N@      �?     �U@       @              &@      $@      S@     �S@      @      K@      R@      @      0@      @     �H@     �j@      .@     �o@      @      @      =@      :@     �j@     �c@      @     @T@      $@       @      @               @      @@      �?     �U@      �?              &@      @     �C@      A@              5@      @              @              @      @      �?      <@                               @      (@      5@              $@                                              �?              ,@                                       @                              @              @              @      @      �?      ,@                               @      $@      5@              $@      @       @       @              @      9@             �M@      �?              &@      �?      ;@      *@              &@      �?               @               @      6@             �H@      �?              &@      �?      3@      "@              @      @       @                      @      @              $@                                       @      @              @     �I@      $@      @      @      5@     �e@      @     0y@      @       @      @      (@      p@     �b@      @     �G@      >@       @      @              3@     �U@      @     �a@      �?      �?      @      @      \@     @S@      �?      :@      7@      @       @              1@      T@      @     �Z@      �?      �?      @      @     @X@     @Q@              6@      6@      @       @              0@     �R@      @      Z@      �?      �?      @      @     @W@     �L@              5@      �?                              �?      @              @                                      @      (@              �?      @       @      �?               @      @              B@                              @      .@       @      �?      @      @       @      �?               @      @              6@                              @      .@      @      �?       @                                                              ,@                                               @               @      5@       @       @      @       @     @V@             @p@       @      �?      @      @     @b@     �Q@       @      5@      1@      �?       @      @      �?      K@             �h@      �?      �?       @      @     �\@      F@              *@      .@      �?       @      @              J@             �c@      �?               @      @     @[@     �E@              (@       @                              �?       @             �D@              �?                      @      �?              �?      @      �?                      �?     �A@             �N@      �?               @      �?      ?@      ;@       @       @      �?                              �?      @               @                       @              $@      @              @      @      �?                              >@             �M@      �?                      �?      5@      6@       @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�ȩhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@��<ٕ�?�	           ��@       	                    @[�T3���?k            �@                            @c8l3��?�           �@                           @�|8��K�?t           ,�@������������������������       �2:��b
�?�           x�@������������������������       ��0�Z�q�?�           h�@                           �?�_��B�?           (�@������������������������       ��%Fs�?�            pw@������������������������       �t4l�\�?/           �~@
                           @�d�`T��?�            �@                          �0@b�5�,1�?m           (�@������������������������       ��� ���?            �G@������������������������       �j[��Y�?R           ��@                            @�Ԕ�M�?{            `g@������������������������       ���8�6L�?j             d@������������������������       �؉�؉��?             :@                           �?&����?           �{@                          �@@D�<���?q            @f@                           @���+��?f            `c@������������������������       ��8��c�?L            �\@������������������������       �@+�*h�?            �D@������������������������       ���;5r�?             7@                           �?�����?�            pp@                            @�q�q�?             H@������������������������       ���4Vk��?            �B@������������������������       �t�E]t�?             &@                           @u) 3�?�            �j@������������������������       �n^���?t            `f@������������������������       �b�2�tk�?             B@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        h@     �B@     �I@      ?@     �[@     x�@     �A@     ��@      *@      @     �R@     @S@     x�@     �@      2@      r@     �d@      >@      F@      >@     �Y@     8�@     �A@     ��@      &@      @      Q@      S@      �@     �}@      ,@     �p@     �`@      9@      @@      8@     �N@     P{@      <@     p�@      $@      @     �M@      P@     �@     0w@      $@     �f@     @Y@      0@      8@      6@      I@     �q@      4@     `z@      $@      @      H@      K@     �t@     0p@      $@     `b@      Q@      ,@      1@      ,@     �C@     �e@      @     �q@      @       @      6@      <@      l@     �_@      @      V@     �@@       @      @       @      &@     �\@      ,@      a@      @      �?      :@      :@     �Z@     �`@      @     �M@     �@@      "@       @       @      &@     �b@       @     �r@              �?      &@      $@     �f@      \@             �A@      8@      @      @               @     �Q@      @     �Z@              �?      @      @      O@     �J@              5@      "@      @       @       @      @     �S@      �?     �g@                      @      @     @^@     �M@              ,@      @@      @      (@      @     �D@     �\@      @      n@      �?      �?      "@      (@     ``@     �Y@      @     �T@      ;@      @      $@      @      <@     @X@       @     �h@      �?              @       @     �X@     @Q@      �?     �L@                                      �?      *@              $@                      �?              �?      $@              &@      ;@      @      $@      @      ;@      U@       @     �g@      �?              @       @     �X@     �M@      �?      G@      @       @       @              *@      1@      @     �E@              �?       @      @      @@     �@@      @      9@      @               @              *@      .@       @      @@              �?      �?      @      =@      ?@      @      7@               @                               @      @      &@                      �?              @       @               @      :@      @      @      �?       @      R@             @e@       @              @      �?     �R@      C@      @      8@      6@      @      @              @      *@              P@                       @              <@      2@      �?      *@      3@      @      @              @      *@              K@                       @              ;@      "@      �?      *@      ,@      @      @              @      (@              ?@                       @              5@      @      �?      $@      @                                      �?              7@                                      @      @              @      @                                                      $@                                      �?      "@                      @      @              �?       @     �M@             �Z@       @              @      �?     �G@      4@      @      &@      �?       @                      �?       @              ,@                                      "@      &@               @      �?       @                              @              @                                      "@      $@               @                                      �?       @              @                                              �?                      @      �?              �?      �?     �I@              W@       @              @      �?      C@      "@      @      "@      @      �?                      �?      D@              T@      �?              @      �?      ;@      "@      @      "@                              �?              &@              (@      �?                              &@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��VhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?綊���?�	           ��@       	                   �<@dr�<_D�?G           ��@                           @%&�D�?            Ș@                           �?�a�]���?Z           X�@������������������������       �����,�?>            ~@������������������������       ��%|��`�?           �|@                          �0@�j�y���?�           8�@������������������������       �r�&�I�?             �I@������������������������       �f��)���?�           ��@
                           �?<�A+K&�?G            �\@                           @����y��?            �G@������������������������       �������?            �A@������������������������       ��8��8��?             (@                          @@@r�G-6z�?,            �P@������������������������       �c}h���?%             L@������������������������       �������?             &@                            @��{0��?{           J�@                            �?��8�Pn�?�           $�@                           @@P����?           d�@������������������������       �#�S����?L           ؀@������������������������       �Mj�h��?�           ��@                           @-s�[��?�             w@������������������������       �y��@:�?�            �l@������������������������       �wtz��t�?Y            `a@                           @g�V�U�?�           ��@                           �?��j���?Y           ��@������������������������       �0 pBX��?]            `b@������������������������       �zx���?�            @x@                           @,�.���?*            @Q@������������������������       ��0\K5��?            �B@������������������������       �     p�?             @@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        g@     �B@      D@      8@     �]@     ��@      ;@     ��@      1@      @      R@      P@     ��@     ��@      4@     �q@     �Y@      6@      ?@      $@     �P@     �s@      *@     Px@      "@      @      <@     �A@     `r@      l@      ,@     �a@     �U@      6@      =@      $@      N@     s@      *@     �u@      "@      @      8@      @@     �q@     �j@      (@     �`@      J@      *@      0@      @      =@     �h@      $@     �k@      @      �?       @      $@     �e@     �_@      @     @P@      @@      "@      ,@       @      *@     @U@      @      ]@      @      �?      @      @     @T@     @Q@       @      C@      4@      @       @       @      0@     �[@      @     �Z@       @              @      @     �V@      M@      @      ;@     �A@      "@      *@      @      ?@     @[@      @     �_@       @      @      0@      6@     �[@     @U@      @     �Q@      @      @                      @       @      �?      "@      �?      �?                      (@      @              "@      @@      @      *@      @      ;@     �Z@       @     �]@      �?      @      0@      6@     �X@     �S@      @     �N@      .@               @              @      *@              D@                      @      @      (@      (@       @      @      �?                              �?       @              1@                      @      @      &@      �?               @                                      �?       @              .@                      @      @      @                      �?      �?                                                       @                                      @      �?              �?      ,@               @              @      @              7@                      �?              �?      &@       @      @      &@               @              @      @              7@                      �?              �?      @       @       @      @                                      �?                                                              @              �?     �T@      .@      "@      ,@      J@     @w@      ,@     ��@       @              F@      =@     �z@      s@      @     �a@     @P@      (@       @      $@     �E@     pp@      (@      }@      @             �D@      8@     �r@     `l@      @     @`@     �G@      &@       @      @      9@      j@      (@     �x@      @              6@      3@      n@      e@      @     �S@      :@      @      �?      @      "@     �W@       @     �c@       @              @      &@     @^@      O@       @     �B@      5@      @      �?      @      0@     �\@      $@     `m@      �?              1@       @      ^@     �Z@       @     �D@      2@      �?      @      @      2@     �K@             �Q@      @              3@      @     �L@      M@       @      J@      (@      �?      @       @      ,@     �E@              H@                      @      @      E@      @@      �?      6@      @              @      �?      @      (@              7@      @              ,@      �?      .@      :@      �?      >@      2@      @      �?      @      "@     @[@       @     `l@       @              @      @     �`@     @S@              (@      0@      @      �?      @      "@     �V@       @     `h@       @              @      @      ^@     �R@              &@      @                      �?              &@             �M@                                     �C@      ?@              @      *@      @      �?      @      "@      T@       @      a@       @              @      @     @T@     �E@               @       @                                      2@              @@                              �?      (@      @              �?       @                                      �?              6@                              �?      "@      �?              �?                                              1@              $@                                      @       @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���;hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx         
                    �?�T=6�?�	           ��@       	                    @��gxM�?6           Ț@                            @
�ߴLL�?/           ��@                            �?v�Y���?            ��@������������������������       � ��{���?�            �w@������������������������       ��lA�_��?	           Љ@                          �9@�3ݏ�?/           �~@������������������������       �������?�            �x@������������������������       ��֥ɴ�??            �W@������������������������       �����W�?             *@                          �;@�-񮣮�?u           .�@                          �9@�J�M��?�           Ğ@                            @������?]           ̛@������������������������       �ء��
��?           ȓ@������������������������       �*n��O��?@           �@                           @t�(!�b�?w            �g@������������������������       �[�x����?Q            @`@������������������������       �	���ĳ�?&             N@                            @	�0�?�            �l@                           @�:�����?q            `d@������������������������       ��tz���?[            @`@������������������������       ��9K�Nq�?            �@@                           �?�@��TM�?0            �P@������������������������       �L䯦s#�?%            �J@������������������������       �N��)x9�?             ,@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@     �B@      F@     �C@     @Z@     h�@      ;@      �@      8@      *@     �Q@     �M@     ��@      �@      0@     0p@     �\@      2@      @@      4@     �Q@     �r@       @     �y@      1@      @      B@      @@     q@     �l@      "@     ``@     �\@      2@      @@      4@     �Q@     �r@       @     �y@      1@      @      B@      @@     q@     �l@      "@      `@     �U@      $@      9@      2@     �M@     �i@      @     �p@      0@      @      =@      =@      e@      e@      "@     �Z@      >@      @       @      @      0@      P@      @      [@                      @      &@     �M@     �G@       @      9@      L@      @      7@      (@     �E@     �a@      @      d@      0@      @      7@      2@     @[@     @^@      @     @T@      =@       @      @       @      &@     �V@       @      b@      �?      �?      @      @     @Z@      N@              6@      6@      @      @       @      $@      U@       @     @[@              �?      @       @      V@      E@              4@      @      @       @              �?      @              B@      �?                      �?      1@      2@               @                                      �?      @              �?                                               @              @     @Z@      3@      (@      3@      A@     �s@      3@     H�@      @      "@      A@      ;@     �z@     �q@      @      `@     �Y@      1@      (@      3@      @@     pq@      0@      �@      @      @      ?@      9@     �w@     q@      @     �^@     @V@      .@      (@      2@      :@     Pp@      .@     X�@      @       @      ;@      9@      t@     �o@      @     �\@     @T@      (@      $@      &@      6@     �f@      (@      w@      @       @      6@      4@     `j@     @i@      @     @Y@       @      @       @      @      @     �S@      @     `k@      �?              @      @     �[@     �J@              ,@      *@       @              �?      @      2@      �?     �L@              @      @             �L@      2@               @       @       @                      @      $@      �?     �C@                       @             �H@      "@              @      @                      �?       @       @              2@              @       @               @      "@               @      @       @                       @     �C@      @     @Y@       @       @      @       @     �I@      *@       @      @       @       @                      �?      7@      @     @P@       @              @       @      E@      (@       @      @       @       @                      �?      2@      @      E@       @              @       @      C@      &@       @      @                                              @              7@                                      @      �?                      �?                              �?      0@              B@               @                      "@      �?              �?      �?                              �?      (@              ?@               @                      @      �?              �?                                              @              @                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJy�zhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @Ip44r��?�	           ��@       	                    �?@��ʇ#�?�           ��@                           �??5�F��?           L�@                           �?D܅��u�?�            �t@������������������������       ����5�?g            �b@������������������������       ��Ⱥ� �?o            �f@                           @B\�=�p�?<           0�@������������������������       ���7�\�?t            `g@������������������������       ���� ]�?�           X�@
                            �?(�� 	��?�           ��@                            �?��K=�?�           Ē@������������������������       ��'kk/��?�           ��@������������������������       ��O�:�E�?s           ؂@                          �1@�Bd
&$�?�            �w@������������������������       ���1��!�?%            �P@������������������������       ���xS��?�            ps@                           �?��6�EL�?�           ,�@                          �:@�w��AJ�?0           ~@                           @0�z �k�?           �y@������������������������       �##$��?�            �p@������������������������       ��!n��x�?X            `a@                          �=@�Gw��?/            @R@������������������������       ��q�q�?             H@������������������������       �Zd;�O��?             9@                           @��_��M�?�           P�@                           �?��֗�l�?(           `}@������������������������       ��Bj�N�?�            @s@������������������������       ���V���?j            @d@                          �;@x�Ӵ��?`            �b@������������������������       ��(\����?P             ^@������������������������       ����S�r�?             <@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      B@     �@@      ;@     �]@     H�@      D@     ��@      3@      @      S@     �R@     ��@     �@      :@     @p@     @f@      4@      7@      7@     �V@      ~@      :@     ��@      $@      @     �Q@      Q@     ��@     �w@      9@     `k@     �S@      (@      0@      "@      K@      m@      *@     �o@      @      @      <@      @@     @i@      f@      $@      \@      (@      @      @       @      1@      M@       @     �R@      �?              *@      @     �G@      E@      �?     �G@      @      @      �?       @      @      3@      �?      C@      �?              "@      @      ?@      1@              *@      @       @      @              $@     �C@      �?      B@                      @      @      0@      9@      �?      A@     �P@      @      $@      @     �B@     �e@      &@     �f@      @      @      .@      :@     `c@     �`@      "@     @P@      4@      �?       @      @      @      ;@      @      B@      �?               @       @      <@      D@              *@      G@      @       @      @      ?@     `b@      @      b@       @      @      *@      8@     �_@     �W@      "@      J@      Y@       @      @      ,@     �B@      o@      *@     z@      @      �?      E@      B@     pt@      i@      .@     �Z@     @Q@      @       @      $@      :@     �h@      "@     �u@      @              .@      6@     �p@     �b@       @     �P@      ?@      @      �?       @      *@     �U@      @      f@      @              @      @      c@      R@      @      9@      C@      �?      �?       @      *@      \@       @     �e@      �?              &@      .@     �[@     @S@      @     �D@      ?@       @      @      @      &@     �H@      @     �P@      �?      �?      ;@      ,@     �O@      J@      @     �D@      @              �?      @              3@              @                      @      @      �?      (@      @      @      8@       @      @              &@      >@      @     �N@      �?      �?      5@      $@      O@      D@      @      B@      E@      0@      $@      @      <@      e@      ,@     x@      "@      �?      @      @     �l@      a@      �?     �D@      8@      $@      @      �?      4@     �T@      "@     �a@      @      �?      @       @     �V@     �Q@              1@      4@      @      @      �?      2@     @S@      "@      \@       @      �?      @       @     @S@     �M@              0@      2@      @      @              "@      N@      @     �M@       @      �?       @       @     �F@     �D@              ,@       @      �?              �?      "@      1@       @     �J@                       @              @@      2@               @      @      @       @               @      @              =@      �?                              *@      &@              �?      �?      @       @                      @              3@                                      @      $@              �?      @                               @      �?              $@      �?                              @      �?                      2@      @      @      @       @     �U@      @     �n@      @               @      @     `a@     �P@      �?      8@      *@      �?      @      @      @      M@      @     �i@      @               @       @      [@      C@              4@      $@      �?      @      @      @     �A@      @     �`@      @               @      �?     �M@      <@              4@      @              �?               @      7@             @R@                              �?     �H@      $@                      @      @                      �?      <@             �C@       @                      @      ?@      =@      �?      @      @      @                      �?      2@              >@                              @      8@      =@      �?      @                                              $@              "@       @                              @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJh�s
hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?47��u�?�	           ��@       	                     @��F�?[           d�@                           @�T�Y�?           L�@                          �1@4��!�o�?�           ܑ@������������������������       �\���4�?�            @o@������������������������       ���Vg��?H           �@                           @��g��?<             W@������������������������       �UUUUU��?             H@������������������������       �9����!�?             F@
                          �5@�[��$=�?<           0�@                           @�������?�            �p@������������������������       �[!���8�?�            �j@������������������������       �	j*D>�?             J@                           @�"�X0�?�            �o@������������������������       �F��O��?s            `h@������������������������       �����h�?%            �M@                           @q� ��?<           �@                           �?�"����?           \�@                            @���4���?           �{@������������������������       ����D��?�             s@������������������������       �P���߶�?Q            �a@                           @t���_��?           `�@������������������������       ������]�?�           ��@������������������������       ��9�u���?           �{@                            @���?)           �}@                          �8@7o�d��?�            �x@������������������������       ��/��w�?�            �t@������������������������       ��������?*             Q@                           �?<��rD �?*            �R@������������������������       ��)O�?             2@������������������������       ���J���?"            �L@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      A@      C@      ,@     �W@     H�@      @@     P�@      9@      @     @U@      J@     ��@     �~@      6@     q@     �X@      7@      :@      @      K@     �r@      3@     �z@      *@       @     �F@      <@     �t@     �l@      "@     �a@      R@      $@      3@      @      E@     `i@      2@     �q@      $@      �?     �A@      ;@      l@     `e@      "@      [@     �Q@      $@      1@      @      D@     `h@      0@     �o@      $@      �?     �A@      :@     `i@      c@      "@     @Y@      0@      @      @      �?      ,@     �A@      "@      ?@      @              $@       @     �E@     �D@      �?      ?@      K@      @      *@      @      :@      d@      @     �k@      @      �?      9@      2@      d@     �[@       @     �Q@       @               @               @       @       @      ;@                              �?      6@      3@              @       @              �?              �?      @       @      &@                                      2@      @              @                      �?              �?      @              0@                              �?      @      *@              @      :@      *@      @      �?      (@     �X@      �?     �b@      @      �?      $@      �?     @Z@      N@              @@      $@      @      @      �?      $@      B@             @U@              �?      $@      �?     �L@      <@              1@      @      @      @      �?      "@      @@              N@                       @              I@      7@              0@      @      �?                      �?      @              9@              �?       @      �?      @      @              �?      0@       @      @               @      O@      �?     �O@      @                              H@      @@              .@      0@      @      @              �?      L@      �?     �E@      @                             �A@      :@               @              @      �?              �?      @              4@                                      *@      @              @      Y@      &@      (@      "@     �D@     �u@      *@     8�@      (@      @      D@      8@     �|@     `p@      *@     �`@     �S@       @      @      @      <@     �q@      (@     �@      "@      @      :@      1@     �w@      j@      @      X@      C@      @      @      �?      @      O@             @]@                      @       @     �]@     �N@      @      :@      C@      @      @      �?      @      H@             @Q@                      @       @     @P@      F@      @      2@                                              ,@              H@                                      K@      1@               @     �D@      @       @      @      8@      l@      (@     �x@      "@      @      3@      .@     `p@     `b@      @     �Q@     �A@      @      �?      �?      .@      c@      @     @p@      @       @      &@      @     �f@      Q@       @     �G@      @      �?      �?      @      "@     �Q@      @      a@      @      @       @       @     @T@     �S@       @      7@      5@      @      @       @      *@      O@      �?     �d@      @              ,@      @     @S@      K@      @     �B@      4@       @      @       @      *@     �K@      �?     @^@      �?              ,@      @      P@      J@      @      B@      4@       @      @       @      "@     �E@      �?     �V@                      ,@      @      H@      I@      @     �@@                                      @      (@              >@      �?                              0@       @              @      �?      �?                              @             �F@       @                      @      *@       @              �?                                                              ,@                              @      �?                              �?      �?                              @              ?@       @                              (@       @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�0�.hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?e࢝��?�	           ��@       	                   �;@Sτ�
�?X           ��@                           @�����?�           �@                            �?4��n��?�           X�@������������������������       ���I��?�            �q@������������������������       ������?�           ȇ@                            @�Dm~ab�?@           P~@������������������������       ������?�            �u@������������������������       ���cZ��?S            �`@
                          �=@�����?w            �g@                            �?H�z�G�?E             Y@������������������������       ��A`��"�?#             I@������������������������       ����1��?"             I@                            �?�������?2            @V@������������������������       �bX9���?             I@������������������������       �~T��@o�?            �C@                          �;@W�����?P           "�@                            @o�z��-�?�           P�@                            �?�rJY��?X           ��@������������������������       ���_�?�           p�@������������������������       �S�w���?�            �t@                           @�$)���?X           X�@������������������������       ��MK,�?           Pz@������������������������       ���}D(�?U            �`@                          �@@�1��/��?�            �o@                          @@@��sd��?�             m@������������������������       ����E��?�             k@������������������������       �����2�?	             .@                          �A@�Ń����?             5@������������������������       ��θ�?	             *@������������������������       �      �?              @�t�bh�h4h7K ��h9��R�(KKKK��h��B�        j@     �@@      D@     �A@     @\@     ��@      ;@     �@      7@      @     @U@      O@     0�@     �@      1@     �p@      V@      3@      ;@      0@     @P@     �r@      1@     �{@      ,@      @     �A@      B@     �q@      m@      @     @`@     �R@      .@      :@      0@      L@     �q@      1@     �w@      (@      @      =@     �@@     Pp@      j@      @     �\@      K@      @      3@      (@     �G@     �h@       @     �p@      @       @      4@      2@     �f@     �_@      @     �R@      0@               @       @      &@     �M@      @     @U@                      @       @      E@      :@       @      0@      C@      @      1@      @      B@     `a@      @     @g@      @       @      .@      $@     @a@     @Y@       @     �M@      5@      &@      @      @      "@     �T@      "@     @Z@      @      �?      "@      .@     @T@     �T@      @      D@      2@      @      @      @      @      O@      "@      Q@      @              "@      (@      I@     �N@      @     �A@      @       @      �?               @      5@             �B@      �?      �?              @      ?@      5@              @      *@      @      �?              "@      3@             @Q@       @              @      @      8@      8@              .@      @      @      �?                       @              C@                      @              1@      "@              (@      @      @      �?                      @              *@                      @               @       @              @      �?                                      �?              9@                                      "@      @              @       @                              "@      &@              ?@       @                      @      @      .@              @      �?                              @      @              6@                                       @      *@              �?      @                              @      @              "@       @                      @      @       @               @     @^@      ,@      *@      3@      H@     `t@      $@     (�@      "@      �?      I@      :@     �z@     @q@      $@      a@     �\@      ,@      *@      .@      F@     @q@      "@     ؂@      @      �?      F@      7@     pw@     �p@      $@     �_@     �X@      *@      "@      *@      B@      i@       @     �w@      @      �?     �C@      5@     @n@     `j@      "@     @Y@      R@      $@       @      $@      6@      c@       @     �t@      @              4@      $@     �h@      b@      @      N@      :@      @      @      @      ,@      H@             �E@      @      �?      3@      &@     �F@     �P@       @     �D@      1@      �?      @       @       @     �R@      �?     `l@                      @       @     �`@     �J@      �?      :@      ,@              @       @      @     �G@      �?      g@                      @       @     �Y@     �A@              3@      @      �?                       @      <@              E@                       @              >@      2@      �?      @      @                      @      @      I@      �?     �Z@       @              @      @      I@      (@              "@      @                      @      @     �E@      �?      Y@       @              @       @     �F@      &@               @      @                      @      �?     �E@      �?      W@      �?              @       @      E@      &@               @                                      @                       @      �?                              @                                                                      @              @                              �?      @      �?              �?                                              @              @                              �?      @                                                                      @               @                                      �?      �?              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx         
                   �0@������?�	           ��@       	                    @��uʛ$�?w            �f@                           �?<�����?o            �e@                            @�Cp��?1            @S@������������������������       �     T�?)             P@������������������������       ��θ�?             *@                           �?UUUUU��?>             X@������������������������       ��q����?            �J@������������������������       ��C�_�;�?            �E@������������������������       �R���Q�?             $@                            @�����u�?,	           $�@                           @!�<<��?�           ��@                          �1@zEDla��?�           (�@������������������������       �B2���?U            �`@������������������������       �B�Z2��?�           �@                            �?]j�-���?�           �@������������������������       �S�F���?<           �~@������������������������       ���.X�$�?L           ��@                           �?���_U�?�           �@                          �;@��x��?�           @�@������������������������       ��^\�$��?Z           ��@������������������������       �dY�a��?8            @T@                           �?pߒ�q�?           �{@������������������������       �Z�^�q�?Q            �`@������������������������       ��%���?�            Ps@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        m@      >@      F@      <@     �[@     Ȅ@      ?@     0�@      0@      &@     @Q@     �N@     ȇ@     �~@      6@     �m@      "@       @       @      @      @     �C@      @      6@      �?       @      @      @      F@      =@      �?      $@      "@       @       @      @      @     �C@      @      5@      �?       @      @      @     �D@      ;@      �?      "@               @       @      @      @      .@       @      $@      �?              @      �?      5@      *@              �?               @       @      @      @      .@       @      @      �?              �?      �?      3@      "@              �?                                                              @                       @               @      @                      "@                      �?              8@      �?      &@               @              @      4@      ,@      �?       @      @                                      $@      �?       @               @              @      ,@      @      �?      @       @                      �?              ,@              "@                                      @       @              @                                      @                      �?                                      @       @              �?     �k@      <@      E@      8@     @Z@     ��@      <@     ؐ@      .@      "@     �P@     �K@     h�@      }@      5@     �l@      e@      3@      ?@      4@     �V@     @{@      5@     0�@      ,@      @      M@      H@     �~@     0t@      ,@     �g@     @U@      ,@      5@      ,@     �C@     �i@      @     �s@      @       @      ;@      7@     @p@     �\@       @     �U@      4@              @               @      >@              1@                      �?      @      ;@      2@      �?      &@     @P@      ,@      1@      ,@     �B@     �e@      @     �r@      @       @      :@      3@      m@      X@      @      S@      U@      @      $@      @     �I@      m@      2@     px@       @      @      ?@      9@      m@      j@      @      Z@      :@       @       @      @      *@      M@      @     �c@      @              @      @     �Z@     @U@      @      *@      M@      @       @      @      C@     �e@      (@      m@      @      @      <@      2@     @_@      _@      @     �V@      K@      "@      &@      @      .@     �g@      @      w@      �?      @       @      @      l@     �a@      @      C@     �F@      @      "@      �?      "@     �W@      @     �j@      �?      @       @      @      ^@     �W@      @      >@      C@      @      "@      �?      @     �U@      @     �e@               @       @      @     �[@     �U@      @      ;@      @                               @       @              D@      �?       @                      "@      @       @      @      "@      @       @      @      @     �W@      @      c@                      @      �?     @Z@     �G@               @      @                              �?      ?@       @      @@                      @             �@@      5@              @      @      @       @      @      @      P@      �?     @^@                      @      �?      R@      :@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJn]	hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?�?gV��?}	           ��@       	                    �?k�s+6�?J           ��@                          �0@�x����?o           ��@                           �?�p=
ף�?             4@������������������������       ��s�n_�?	             *@������������������������       ��$I�$I�?             @                          �>@u6B7�?`           ��@������������������������       �C��.�?L           ��@������������������������       �     `�?             @@
                          �?@qUh4�?�           T�@                          �1@DCǺ&@�?�           �@������������������������       �QM�ı��?�             m@������������������������       �d*a����??           Ќ@������������������������       �B+K&:~�?             3@                            @CI�ܠ�?3           Ƞ@                          �4@g�����?�           x�@                          �0@jPEQ1�?�           ��@������������������������       ��c���+�?/            �S@������������������������       ��^&MI��?~           H�@                          �;@4�T���?           8�@������������������������       �w�#�A�?�           ��@������������������������       ��<y����?p            �f@                           @�!����?p           0�@                           @Nݹ��A�?           |@������������������������       ��"L���?�            �u@������������������������       �r�Kv׏�?=            �X@                           @o�2���?T            �`@������������������������       �t�M�.�?G            �[@������������������������       ��Z�Y��?             7@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      >@     �@@      =@     �W@     ؃@     �@@     Ȑ@      7@       @     �U@     �O@     ��@     8�@      3@     Pq@     �Z@      1@      6@      .@      M@      r@      2@     Py@      .@      @     �F@      >@     pu@     @o@       @      a@     �B@      "@      &@      @      6@     @X@      @     @c@      @      �?      4@       @     @X@     �T@       @      C@                                       @                      �?                       @      @      @       @              �?                                       @                      �?                       @      @      �?      @                                                                                                                       @      @              �?     �B@      "@      &@      @      4@     @X@      @      c@      @      �?      2@      @     �W@     �R@       @     �B@     �A@      "@      &@      @      4@      W@      @      a@      @      �?      2@      @     �V@     @R@      �?      B@       @                                      @              1@                                      @       @      �?      �?     �Q@       @      &@      "@      B@      h@      .@     `o@      &@      @      9@      6@     �n@     �d@      @     �X@      Q@       @      &@      "@      B@      h@      .@     �m@      &@      @      9@      6@     @n@     �d@      @     �X@      (@      �?      @       @      $@     �B@      @      =@      @       @      "@      @      E@     �A@       @      A@      L@      @      @      @      :@     �c@      (@      j@       @      @      0@      .@      i@     �`@      @      P@       @                                                      *@                                      @                             �\@      *@      &@      ,@     �B@     �u@      .@     �@       @       @     �D@     �@@     �z@     �p@      &@     �a@     @Y@      *@      @      $@      ?@      p@      &@     {@      @       @     �A@      7@     �q@     �l@      $@     @]@     �H@       @      @      @      "@      _@       @      d@      �?              3@      .@     �]@      [@      "@     �O@      @                       @              .@              "@                      �?      @      0@      &@              *@     �E@       @      @       @      "@     @[@       @      c@      �?              2@      $@     �Y@     @X@      "@      I@      J@      &@       @      @      6@     �`@      @      q@      @       @      0@       @     �d@     @^@      �?      K@     �G@       @       @      @      6@      W@      @     �j@       @       @      0@      @     @_@     @[@             �D@      @      @               @              D@              N@      �?                       @     �D@      (@      �?      *@      ,@              @      @      @     @V@      @     �m@      @              @      $@     `a@      D@      �?      8@      &@              @      @      @      K@      @     �h@      @              @       @      [@      :@              2@      @              @      @      @      D@      @     `b@      �?              @       @     �V@      3@              1@      @                              �?      ,@             �I@      @                              2@      @              �?      @                               @     �A@              C@                      �?       @      ?@      ,@      �?      @      @                               @      >@              9@                               @      =@      *@      �?      @                                              @              *@                      �?               @      �?              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��p(hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?��*&�r�?�	           ��@       	                   �=@l���V4�?Z           ��@                            �?���/�?-           ��@                           @i���K�?           `z@������������������������       �ƨ\�x��?�            Pt@������������������������       ��~	c���?A            @X@                          �1@�D�a5h�?'           ��@������������������������       �    ���?�             p@������������������������       ����d3:�?�           ��@
                          �?@��P�M��?-            �N@                            �?�������?            �@@������������������������       �d�����?             3@������������������������       ��>4և��?             ,@                            �?/����?             <@������������������������       �     @�?             0@������������������������       �      �?
             (@                           @��ڳ�?P           Р@                            @�R��۴�?$           `�@                            �?��6w@�?�           Б@������������������������       �������?7           ��@������������������������       ��6�!z��?�             l@                           �?[�Lb	P�?W            �@������������������������       ��qǞ�?�             x@������������������������       ��]��\��?e            �d@                            �?����x[�?,            }@                           @S;�@b�?F            �[@������������������������       �/�5���?            �D@������������������������       ��j����?-            @Q@                           @dw���?�             v@������������������������       �n��<�)�?k            �d@������������������������       ������?{            �g@�t�b�     h�h4h7K ��h9��R�(KKKK��h��B�       �i@      C@      A@      B@      ]@     �@      <@     ��@      3@      $@      Q@     �N@     �@     �}@      3@      n@     @Z@      9@      9@      7@     �R@     �s@      1@     �z@      ,@      @      ?@      >@     �s@     �i@      (@     �`@     �W@      9@      9@      7@     @P@     Ps@      1@     �y@      *@      @      ?@      <@     `s@     @i@      &@     �`@      0@      @      @      @      *@      U@      @     �_@       @              @      $@      R@      G@      @      8@      &@       @      �?      @      &@     @P@      @     @Z@       @              @      "@      N@      <@      �?      *@      @      �?       @               @      3@      �?      6@                      �?      �?      (@      2@       @      &@     �S@      6@      6@      0@      J@      l@      (@     �q@      &@      @      8@      2@     �m@     �c@       @     @[@      1@       @      @              3@     �F@      @     �B@      �?              @      @     �I@      @@       @      =@      O@      4@      2@      0@     �@@     �f@      @     �n@      $@      @      2@      ,@     `g@      _@      @      T@      $@                              "@      @              4@      �?                       @      "@      @      �?      �?      @                              "@      �?              "@                               @      @      �?      �?      �?                                      @                       @                                      @                      �?      @                               @      �?              �?                               @       @      �?      �?              @                                       @              &@      �?                              @      @                                                               @              @                                      @      @                      @                                                      @      �?                              �?                             �X@      *@      "@      *@      E@     Pv@      &@     ��@      @      @     �B@      ?@     0|@     �p@      @     �Z@      U@      &@      @       @      9@     �q@      "@     @�@       @      @      =@      0@     �w@     `l@      @     @S@      P@       @      @      @      6@     �h@      "@      t@       @      @      9@      (@     �m@     �d@      @     �M@     �H@      @       @      @      .@     �c@      @     �q@       @              .@      "@     `h@     �_@       @     �D@      .@       @      @              @     �B@      @     �C@              @      $@      @     �E@     �B@      @      2@      4@      @      �?       @      @     @U@              i@               @      @      @     �a@     �O@      �?      2@      1@       @               @       @     �O@              b@               @      @      @     �S@      G@      �?      2@      @      �?      �?              �?      6@             �K@                      �?             �O@      1@                      .@       @       @      @      1@      S@       @     �e@      @               @      .@     �Q@     �E@      �?      >@      @       @              @      @      ,@             �I@                              �?      1@      &@      �?       @      @       @               @              �?              2@                                       @      @              �?                               @      @      *@             �@@                              �?      "@      @      �?      �?      &@               @      �?      ,@      O@       @     �^@      @               @      ,@      K@      @@              <@      @              �?              @      =@       @      P@                      @       @      *@      0@              .@      @              �?      �?      @     �@@             �M@      @              @      @     �D@      0@              *@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��UhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�^�?�	           ��@       	                     @0���?<           ��@                          �0@�=��Yg�?           ,�@                           �?"�$�F�?7            �W@������������������������       �v0f��#�?             K@������������������������       �\F���?            �D@                            �?��>�J�?�           ��@������������������������       �'�� ���?           p�@������������������������       �-�S��?�            �q@
                           @h��(�+�?7            @                           @���8���?           �{@������������������������       ��#�Q�?            z@������������������������       ����QI�?             9@                           @[��b���?%            �K@������������������������       ���QN�?             ?@������������������������       �9��8���?             8@                            @��M�4��?_           �@                           �?�%�h�&�?�           ��@                           @��,�?	           �y@������������������������       �^&�I�o�?�            `t@������������������������       ����By�?:            @V@                            �?2��B��?�           �@������������������������       ��Ͼ�WO�?'           Ћ@������������������������       ��!B3#��?�            �p@                           @�K��@�?�           P�@                           @�^�⳿�?b           ��@������������������������       �Ծ�����?
           p{@������������������������       ��qK��?X            �`@                           @p�u=q��?             G@������������������������       �6�d�M6�?            �@@������������������������       ��5��?             *@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      ?@      A@      <@     @[@     ��@      ?@     P�@      &@      &@     �U@     �Q@     �@     �@      6@     `n@     @Y@      .@      7@      ,@     �P@     `r@      ,@     @{@      @       @      G@      D@     �q@      o@      @      _@      S@      "@      2@      $@     �G@      j@      $@     �q@      @      @      B@     �B@     `h@     �f@      @     @Y@      @      �?      �?              &@       @      @      (@               @       @       @      .@      :@               @              �?      �?              &@      @      @      @                              �?       @      0@                      @                                      �?              @               @       @      �?      @      $@               @     @R@       @      1@      $@      B@      i@      @     �p@      @      @      A@     �A@     �f@     �c@      @     @W@     �M@      @      ,@      "@      :@     @d@      @     `k@      �?      �?      :@      2@      b@     �W@      @     �N@      ,@      @      @      �?      $@     �C@       @     �I@       @       @       @      1@     �A@     �O@       @      @@      9@      @      @      @      3@     @U@      @     @c@      �?      @      $@      @     �V@     @P@              7@      8@      @      @              (@     @S@       @      b@      �?      @      @      @     �T@     �L@              4@      8@      @      @              (@     �R@       @     �_@      �?      @      @      @     �S@     �L@              3@                                               @              2@                      �?              @                      �?      �?      �?              @      @       @       @      "@                      @              "@       @              @      �?                      @      @      �?              @                       @              @      @              @              �?                      @      @       @      @                      �?              @      �?                      V@      0@      &@      ,@     �E@     �t@      1@      �@      @      @     �D@      ?@     @|@     `p@      0@     �]@     �P@      $@      "@      (@      ?@     �l@      1@     @~@      @      �?      D@      ;@      t@     �i@      .@      X@      4@       @       @      @      *@     �P@      @     �[@      �?              @      $@     @Y@      M@       @      .@      3@       @       @      @       @     �K@      @     �S@                      @      @     �S@     �I@       @      (@      �?                              @      (@             �@@      �?                      @      7@      @              @      G@       @      @      "@      2@     @d@      ,@     Pw@      @      �?     �@@      1@     �k@     �b@      *@     @T@      >@      @       @      @      &@      `@      "@     �s@      @              1@      *@     �f@      Z@      $@      I@      0@       @      @       @      @     �@@      @     �K@      �?      �?      0@      @      D@      F@      @      ?@      6@      @       @       @      (@     �Y@             �o@       @       @      �?      @     @`@      L@      �?      7@      2@      @       @       @      (@      U@              n@      �?       @      �?      @      _@      K@      �?      4@      &@      @       @       @      $@      L@             `i@      �?       @              �?      X@     �A@              1@      @      @                       @      <@              C@                      �?      @      <@      3@      �?      @      @                                      3@              &@      �?                              @       @              @      @                                      $@              "@      �?                              @       @               @                                              "@               @                                      �?                      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJt�EhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?)��H.��?�	           ��@       	                    �?���i���?�           �@                           �?ܷ�k�?�?�           8�@                          �2@��@N�h�?8            �V@������������������������       ��!�>���?            �A@������������������������       �D'0���?$            �K@                          �<@�qH��?f           h�@������������������������       ��!L���?R           X�@������������������������       ��)�8��?             A@
                            @]�n����?U           ��@                          �2@�ir:(��?�            px@������������������������       �F�{0X��?T            �a@������������������������       ��5��l�?�            `o@                           @A���!�?b            �a@������������������������       �>��\<%�?V            �_@������������������������       �����>�?             ,@                          �<@L��Un~�?�           �@                           @b[���?=           2�@                            @Ϟ��<��?�           ��@������������������������       ��=μ�?M           H�@������������������������       �d%�=�?�           ��@                           �?�$�~�?n           ��@������������������������       ���f��?             C@������������������������       ��'�����?T           `�@                          �@@�s��LR�?�            �n@                           �?��[q{��?�            @k@������������������������       �T�r
^N�?             <@������������������������       ����>`��?r            �g@                            �?��S����?             ;@������������������������       �ݾ�z�<�?
             *@������������������������       ���X��?             ,@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@     �A@     �I@      =@     �X@     �@     �@@     ̐@      (@      @      U@      L@     �@     ��@      5@     �p@     �T@      @      1@      (@      ?@     @h@      @     r@      @              9@      4@     �p@     `d@       @     @V@      G@      @      (@      @      6@     �_@      @      `@      @              7@      (@     `a@      Z@       @     �F@      @      �?      �?              @      &@              6@                      @      @      "@      0@              &@      �?              �?                      @              ,@                              @       @      @               @      @      �?                      @       @               @                      @              @      $@              "@      E@      @      &@      @      3@      ]@      @     �Z@      @              1@      @     @`@      V@       @      A@     �D@      @      &@      @      2@      ]@      @     @W@      @              (@      @     �^@     �U@       @      =@      �?                              �?                      ,@                      @              @      �?              @     �B@              @      @      "@     �P@       @      d@       @               @       @     ``@     �M@              F@      B@              @      @      "@      M@       @      X@       @              �?      @     �V@     �H@              ?@      2@              @       @      �?      =@              <@                              @      A@      $@              $@      2@               @      @       @      =@       @      Q@       @              �?       @      L@     �C@              5@      �?                      �?              "@              P@                      �?      �?     �D@      $@              *@                              �?               @              L@                      �?             �C@      $@              (@      �?                                      �?               @                              �?       @                      �?      _@      ?@      A@      1@      Q@     �}@      ;@     ��@      @      @     �M@      B@     0}@     �v@      3@     �f@     @\@      >@      A@      1@      P@     P{@      :@     �@      @      @     �K@      A@     �z@     v@      3@     `d@     �W@      9@      8@      &@     �C@     �v@      5@     �~@      @      @      C@      <@     �t@     Pr@      *@     �Z@     �Q@      6@      *@      $@      >@     �n@      2@     �r@      @      @     �@@      3@     �i@     �j@      &@     �X@      8@      @      &@      �?      "@     @^@      @     @h@      �?      �?      @      "@     @_@      T@       @       @      2@      @      $@      @      9@     �Q@      @     @f@               @      1@      @     @X@      N@      @     �L@                              @              *@      �?      .@                      �?      �?      @                              2@      @      $@      @      9@     �L@      @     `d@               @      0@      @     @W@      N@      @     �L@      &@      �?                      @      C@      �?     @\@       @      �?      @       @      C@      *@              1@       @      �?                      @      B@      �?     @Z@       @      �?      @              >@      "@              1@       @                              �?      @              "@                      �?                      @              @      @      �?                      @      ?@      �?      X@       @      �?      @              >@      @              &@      @                                       @               @                               @       @      @                                                               @              �?                               @      @      @                      @                                                      @                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��QFhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B(                             !@��Q�(}�?�	           ��@       	                    @�H�d#|�?�	           `�@                           �?�M��o�?c           Л@                           �?���R���?!           4�@������������������������       �^�q�"c�?<           �@������������������������       ��l�����?�           ��@                           @٥a�d�?B           p~@������������������������       ���wu^�?           �z@������������������������       ��w����?+             O@
                            @pt�b�}�?9           x�@                          �7@�>ȇ��?�           �@������������������������       ����2�?�           p�@������������������������       �*�bR8��?           �z@                           �?5h�"��?j           ��@������������������������       �1f߻��?�            �q@������������������������       ����[���?�             r@                           @Dio����?             9@������������������������       �      �?             0@������������������������       ���E���?             "@�t�bh�h4h7K ��h9��R�(KKKK��h��B�	       @j@     �@@      :@      5@      \@     �@      <@     T�@      *@      @      T@     �R@     p�@     p@      .@      p@      j@     �@@      :@      5@      \@     ��@      ;@     H�@      *@      @      T@     �R@     `�@     P@      .@     p@      Y@      ,@      (@      (@      P@     �r@       @     �@      @      @     �B@      C@     w@      h@      @      \@     �T@      @      @       @     �G@     @l@      @     �u@      @       @      >@     �A@      o@      d@      @      U@      :@      �?      @      �?      3@     @U@             `c@                      4@      (@     �S@     �Q@      �?      B@      L@      @      @      @      <@     �a@      @     �g@      @       @      $@      7@     `e@     @V@      @      H@      2@      $@      @      @      1@     �R@      @     @d@              �?      @      @      ^@     �@@      �?      <@      2@      $@      @      �?      .@     �P@      @      b@              �?      @      @      Y@      7@      �?      <@                      �?      @       @      "@              1@                                      4@      $@                      [@      3@      ,@      "@      H@     `v@      3@     ��@       @      @     �E@     �B@     �w@     @s@      $@      b@      V@      &@      (@      "@      C@     �n@      1@     y@      @       @     �B@      ?@     q@     �l@       @     �`@     �S@      &@      (@       @      ;@      e@      (@     Pp@      @       @      ;@      ;@     �i@     @f@      @     �V@      $@                      �?      &@      S@      @     �a@       @              $@      @     @Q@      J@       @      E@      4@       @       @              $@     @\@       @     �h@       @       @      @      @     �Z@     �S@       @      *@      .@      @       @               @     �F@       @     @W@       @       @      @      @     �D@      H@       @       @      @      @                       @      Q@             @Z@                       @      �?     @P@      >@              @       @                                      ,@      �?      @                                       @       @              �?       @                                      "@      �?      @                                              �?                                                              @                                                       @      �?              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��(EhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?�!����?�	           ��@                          �1@�wc��U�?9           �@                           @1�BZx��?�            �r@                           @�ͧ$���?�            �q@������������������������       ��qH-��?�             m@������������������������       �k�����?            �J@������������������������       ���2Tv�?	             .@                           @�/z�?z           T�@	       
                     @���?8           ԓ@������������������������       �a�I�!J�?7           �@������������������������       �
�ӽZ�?           �w@                           �?�����Z�?B             X@������������������������       ��K8��?              J@������������������������       �.�袋.�?"             F@                          �;@�L߆t��?p           ��@                           @�_t��?�           �@                            @c���$�?�           Ș@������������������������       �6�@����?�           ��@������������������������       ��p:��{�?/           �|@                          �4@*ں��?�            �x@������������������������       � a~L;��?�            �j@������������������������       �!kOLI�?p            `f@                           @���d��?�            �p@                           @C��.q�?�            �l@������������������������       ���p/"�?m            �f@������������������������       ��q�q\�?!             H@                            �?�Rͦ$�?            �B@������������������������       �T�r
^N�?             ,@������������������������       �I�O���?             7@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      C@      B@      :@     @]@      �@      A@     (�@      5@      @     �Q@      R@     P�@     �@      1@      p@     �Z@      7@      >@      "@     �Q@     Pt@      .@     0w@      (@      @     �@@     �@@     `q@     @j@      @     `a@      0@       @      $@              ,@      N@      @      B@      �?      �?       @      ,@     �G@     �F@      �?     �C@      0@       @      @              $@      N@      @      A@      �?      �?       @      ,@     �G@     �D@      �?      C@      ,@       @      @              @     �I@      @      6@      �?      �?       @      ,@      D@      ?@      �?      A@       @              @              @      "@      �?      (@                                      @      $@              @                      @              @                       @                                              @              �?     �V@      5@      4@      "@     �L@     �p@       @     �t@      &@       @      9@      3@     �l@     �d@      @      Y@     �U@      5@      3@      "@     �L@     0p@      @     ps@      "@       @      9@      3@      i@     �b@      @     @V@      N@      *@      .@      "@     �D@     @h@      @     �h@      @      �?      3@      0@     ``@     @[@      @     �Q@      ;@       @      @              0@     @P@       @     @\@      @      �?      @      @     �Q@      D@              2@      @              �?                      @       @      8@       @                              >@      0@              &@      @                                      �?              ,@                                      6@      @               @      �?              �?                      @       @      $@       @                               @      (@              @     �\@      .@      @      1@      G@     �u@      3@     ��@      "@      �?      C@     �C@     @{@     �r@      $@     @]@     �Z@      ,@      @      0@      F@     pr@      3@      �@      @      �?     �A@      B@     �x@     pq@      @      [@     �W@      "@      @      ,@      >@     �m@      0@     �}@      @      �?      :@      ?@     pt@     �m@      @      S@      S@      @      @      &@      7@     �e@      .@     �r@      @      �?      9@      6@     �j@     �f@      @     @P@      2@      @      �?      @      @      O@      �?     `e@      �?              �?      "@      \@     �M@      �?      &@      *@      @      �?       @      ,@     �M@      @     �a@       @              "@      @     �P@      D@       @      @@       @       @               @      @      ;@      @     @V@       @              @       @      =@      5@      �?      0@      @      @      �?              @      @@             �I@                      @      @     �B@      3@      �?      0@       @      �?              �?       @      L@             �\@       @              @      @     �E@      6@      @      "@       @      �?              �?       @     �I@              V@       @              @      �?      D@      6@      @      "@       @      �?              �?       @      A@             �S@       @              @      �?      ;@      ,@      @      "@                                              1@              $@                                      *@       @                                                              @              ;@                               @      @                                                                      �?              "@                               @       @                                                                      @              2@                                      �?                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�1�ohG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�}�)�|�?�	           ��@       	                    @e��	z�?C           ؚ@                          �=@@�<b���?�           ��@                          �0@~E�Kz��?p           ��@������������������������       � 9�����?             F@������������������������       ��B� ���?S           ��@                          �?@:����?+            �Q@������������������������       ���{�~�?             E@������������������������       ��ΑL�?             =@
                           �?C���@O�?�           ��@                           @"�t�q�?�            �o@������������������������       �a5�;�H�?Y            �`@������������������������       ���C�E��?M            @^@                          �1@j�ٷ2�?           @y@������������������������       ��iP7�?=            �Y@������������������������       ����;ƈ�?�            �r@                          �;@�ګ;��?b           &�@                          �0@N-V�i�?�           ��@                           @�E��Y�?<            �[@������������������������       �y'�L��?/             U@������������������������       �PS!����?             :@                            @V���?y           ��@������������������������       �N-�Gvb�?/           �@������������������������       ���>���?J           �@                          �=@�x
�2�?�            �r@                            @*��T8�?F            �^@������������������������       �&ޏ���?1             V@������������������������       ��aE'��?            �A@                           @ϡc��w�?g            �e@������������������������       �B�,V ��?0            �S@������������������������       ���ЇL��?7            �W@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      >@      F@      9@      Y@     ��@      ?@     @�@      1@      @     �O@      P@     ��@     ��@      3@      o@      U@      0@     �A@      0@     �N@      u@      ,@     `y@      (@      @      <@      ;@     pq@     0p@      $@      `@      L@      &@      ?@      @      C@     @l@       @      p@      @       @      &@      $@      e@     �b@      @     �R@      I@      &@      ?@      @      @@     �j@       @      l@      @       @      &@      $@     �d@     �a@       @     �R@                       @              @      $@      �?      �?                               @      $@      (@              @      I@      &@      =@      @      =@     �i@      @     �k@      @       @      &@       @     `c@      `@       @     �Q@      @                              @      (@              @@                                      @      "@      �?      �?      @                              @       @              5@                                      @      @      �?      �?      @                                      $@              &@                                              @                      <@      @      @      $@      7@     �[@      @     �b@      @      @      1@      1@     �[@     @[@      @      K@      "@       @       @      @      "@     �G@              F@      @              @      @     �H@      F@      @      5@      @       @                      @      ;@              2@      @              @      @      A@      ,@      @      "@      @               @      @       @      4@              :@                       @      �?      .@      >@              (@      3@      @       @      @      ,@     �O@      @     �Z@      �?      @      $@      (@     �N@     @P@       @     �@@       @               @              @      *@      @      1@              @      @      @      2@      1@              $@      1@      @              @      "@      I@      @     @V@      �?              @       @     �E@      H@       @      7@     �\@      ,@      "@      "@     �C@     @t@      1@     Ѕ@      @      �?     �A@     �B@      |@     �s@      "@      ^@     �Y@      &@      "@       @      B@     �p@      *@     �@       @      �?      ?@      A@     px@     �r@      @      [@      @                                      9@              4@                      �?      @      9@      2@              $@      @                                      7@              2@                      �?      @      2@      @              $@      �?                                       @               @                                      @      ,@                     �X@      &@      "@       @      B@     `n@      *@     p�@       @      �?      >@      <@     �v@     �q@      @     �X@      U@       @      @      @     �@@     �e@      &@      w@      �?      �?      =@      5@      o@     �j@      @      S@      ,@      @      @       @      @      Q@       @     �g@      �?              �?      @     �]@     �Q@       @      6@      &@      @              �?      @      L@      @      ^@      @              @      @     �L@      .@      @      (@      "@      �?              �?              6@             �L@                       @              .@      "@      @      @      "@      �?              �?              .@              A@                       @              ,@      @      @      @                                              @              7@                                      �?      @              �?       @       @                      @      A@      @     �O@      @               @      @      E@      @      �?       @       @       @                      @      4@      @      9@      @               @       @       @      �?      �?      @                                              ,@              C@                              �?      A@      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJU��{hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @ܕ����?�	           ��@       	                   �0@�XV��?�           �@                            �?�2�/��?r            �f@                           �?P1n��?%             M@������������������������       ���R[s�?            �A@������������������������       �T#G�h�?             7@                           @r��%3@�?M             _@������������������������       ��r8��?=            �W@������������������������       �CbΊx�?             =@
                            �?�m�T��?�           ��@                           �?�k��`�?�           4�@������������������������       ��3�1��?+            �@������������������������       �H�%����?�           $�@                           �?�^q��?�           ��@������������������������       ���])���?I            �\@������������������������       �������?X           `�@                           �?��d'8�?�            �@                          �6@?�0w�A�?2           0~@                          �0@� �?�            0q@������������������������       �������?             2@������������������������       �1��:���?�            p@                           �?n_Y�K�?�             j@������������������������       �V&k{L��?)            �R@������������������������       �>��t��?X            �`@                           �?���=-�?�           (�@                           @E
o*'��?�            �w@������������������������       ��x��.�?�             q@������������������������       ��WV��?@             Z@                           @��`�'�?�            `m@������������������������       ��t��*�?o             e@������������������������       ��e�i���?&            �P@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@      >@     �D@      8@     �X@     8�@      <@     d�@      7@       @     @V@      N@      �@     �@      7@     �q@     @b@      6@      <@      5@      S@     0}@      9@     ��@      3@       @     �T@      G@     �@      x@      4@      m@      @               @      �?      @      7@       @      9@      �?      �?       @      @     �B@      H@      �?      1@      �?                              �?       @       @      &@                      @              *@      1@               @                                      �?      @       @       @                                      @      *@              �?      �?                                      @              @                      @               @      @              �?      @               @      �?      @      .@              ,@      �?      �?      @      @      8@      ?@      �?      .@      @               @      �?      @      ,@              *@      �?      �?      @      @      2@      .@              .@       @                               @      �?              �?                                      @      0@      �?             �a@      6@      :@      4@     �Q@     �{@      7@     ��@      2@      @     �R@      E@     �}@      u@      3@     �j@     �Y@      0@      0@      .@      F@      u@      1@     X�@      (@      �?     �L@      1@     �w@     �n@      (@      a@      M@      @      &@      @      :@     �c@      @      n@      @      �?     �@@      &@     �b@     �X@      @      U@      F@      $@      @      $@      2@     �f@      &@     �u@      @              8@      @      m@      b@      @      J@      C@      @      $@      @      :@     �Z@      @      ]@      @      @      2@      9@     �V@     �W@      @     �S@      @      @      @      �?       @      5@              ,@      @              @       @      *@      *@      @      9@      A@      @      @      @      8@     @U@      @     �Y@      @      @      ,@      7@     @S@     @T@      @      K@     �K@       @      *@      @      7@     �f@      @     x@      @              @      ,@     �l@     @^@      @      H@     �C@      @      "@              .@     �S@      @     @b@      �?              @      @      V@     �P@       @      5@      (@      @      @              ,@     �D@      @     �W@                      @      @     �E@     �@@              1@      �?                              @               @      �?                      �?       @      @       @              @      &@      @      @              &@     �D@      �?     @W@                       @      @      D@      ?@              ,@      ;@       @      @              �?     �B@              J@      �?                      �?     �F@     �@@       @      @       @                                      (@              ,@                              �?      0@      4@              @      3@       @      @              �?      9@              C@      �?                              =@      *@       @      �?      0@       @      @      @       @     �Y@             �m@      @              @       @     �a@     �K@      �?      ;@      "@               @      @      @     �O@             `a@      �?              �?      @     �T@      E@      �?      8@      @               @      @      @      B@             �[@      �?              �?      @      O@      8@              5@      @                              �?      ;@              =@                              �?      5@      2@      �?      @      @       @       @              @     �C@              Y@       @               @      @     �M@      *@              @      @               @              @      8@             �S@                       @             �E@      &@                       @       @                              .@              6@       @                      @      0@       @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�6++hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�͓.���?�	           ��@       	                     �?Po*Z��?�           ��@                          �<@��۟��?/           t�@                          �0@����Z��?�           8�@������������������������       ��=�@4��?T            �`@������������������������       ��l0-F��?f           �@                           �?f)}8�I�?u            �e@������������������������       ������?/            �Q@������������������������       �v�f��?F            �Y@
                           @&N�)1�?�           ��@                          �9@��� ��?�            @r@������������������������       �;G���?�            �l@������������������������       �     @�?*             P@                           �?��(�1�?�            @w@������������������������       �	��	�?L            �^@������������������������       �* ��q�?�            @o@                           �?Sj�L�?�           ܑ@                          �3@׆�[	��?�           ��@                          �0@Lt�<��?�            �l@������������������������       �M�h���?             :@������������������������       �ID���/�?x            @i@                          �;@�#3����?)            }@������������������������       ��nΛ��?�            pw@������������������������       �!Θ�?:            @V@                           @�������?           0|@                           @��f���?y            `i@������������������������       ��ӭ�a�?V             b@������������������������       ���_#w��?#            �M@                           �?�/�n��?�             o@������������������������       �Y�5���?N            �`@������������������������       �����?Q            �\@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @j@      9@     �B@      @@     @V@     �@     �B@     ��@      6@       @     @U@     �Q@     ��@     �@      6@     �o@     `c@      0@      <@      <@     �Q@     @}@      ?@     ��@      2@      @      S@      J@     (�@     �w@      5@     �i@      \@      (@      2@      7@      B@     @w@      4@     �@      *@      �?     �J@      <@     �y@     `q@      *@     @a@     �Z@      (@      .@      7@      A@     �t@      4@     �@      &@      �?     �I@      <@     �w@     �p@      *@     @`@      @               @      �?      @      9@      @      6@      @              �?              ?@      8@              &@     �Y@      (@      *@      6@      ;@     Ps@      1@     �~@       @      �?      I@      <@     �u@      n@      *@     �]@      @              @               @      C@             �P@       @               @              @@      ,@               @      @              @               @      $@              ?@                       @              @      "@               @      �?                                      <@             �A@       @                              9@      @              @     �E@      @      $@      @      A@      X@      &@     �]@      @      @      7@      8@     @Z@     @Z@       @     �P@      .@      @      @      @      .@     �B@       @     �H@      @              (@      �?     �F@     �K@      @     �D@      *@              @      @      .@      :@             �A@      @              @      �?      E@     �F@      @      ?@       @      @                              &@       @      ,@                       @              @      $@      �?      $@      <@      �?      @       @      3@     �M@      "@     �Q@       @      @      &@      7@      N@      I@      @      :@      @      �?      @      �?      &@      "@       @      ,@       @      @       @       @      >@      *@              .@      5@              �?      �?       @      I@      @      L@              �?      "@      .@      >@     �B@      @      &@     �K@      "@      "@      @      3@     �i@      @     px@      @       @      "@      2@     �m@     �_@      �?     �G@     �E@      @       @      @      $@     �\@      @     @m@      @       @      @      *@     �_@     �U@      �?     �@@      ,@               @       @      @      @@      @      K@                      �?      @     �F@     �G@              0@                                      @                      @                      �?      @      �?       @              @      ,@               @       @      @      @@      @     �I@                              �?      F@     �C@              $@      =@      @      @       @      @     �T@       @     �f@      @       @      @       @     �T@      D@      �?      1@      5@      @      @       @       @      O@       @      a@       @       @      @      @      S@     �B@      �?      *@       @                               @      4@              F@      �?                      �?      @      @              @      (@      @      �?              "@     �V@             �c@      �?              @      @     �[@     �C@              ,@       @       @      �?              @      9@             �M@                      @      @     �Q@      5@              @      @       @                      @      0@             �F@                       @              M@      "@              @       @              �?               @      "@              ,@                      �?      @      (@      (@              @      @      @                      @     �P@             �X@      �?               @       @     �D@      2@               @      �?      @                      @      D@             �H@                      �?       @      4@      @              @      @      �?                              :@             �H@      �?              �?              5@      (@              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJw��QhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@y۾bp�?�	           ��@       	                    @(>���?�           Z�@                          �:@��z���?~           ��@                          �0@�����??           ��@������������������������       ��@��,�?i            `d@������������������������       ��G6C��?�           ��@                            �?�$�ny��??            �W@������������������������       ����c�H�?$            �H@������������������������       ���g��?             G@
                            @�Bi�qi�?           ��@                           �?��͏��?�           0�@������������������������       ��w��?�            �r@������������������������       �|'8�8�?�            �u@                           @��L���?�            @i@������������������������       ��Iy4�%�?o            `d@������������������������       �ۛ�xt�?            �C@                           @��*�>��?	           �y@                          �=@0=�W���?�            �v@                           @E��!�?n            �e@������������������������       ��5�O[�?[            �a@������������������������       ��B'U�?            �@@                          �?@�����?             g@������������������������       ���r��?I            �[@������������������������       �d�&����?6            �R@                          �?@�m��1�?             J@                            �?j��ۑ�?            �B@������������������������       �8�Z$���?             *@������������������������       �      �?             8@������������������������       �n�����?             .@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        k@      ;@      D@      ;@      \@     X�@      <@     ��@      2@      @     @U@      J@     ��@     �~@      8@      o@      i@      6@     �B@      9@     �Y@     P�@      :@     @�@      ,@      @     �R@      H@      �@     0}@      5@     �l@     `d@      *@      =@      7@     @U@     z@      3@     @�@      @      @      P@     �B@     �@     ps@      ,@     �f@     @d@      $@      <@      7@     �T@     0y@      3@     p�@      @      @      P@      B@     �@     �r@      ,@     �f@      @              �?       @      @      =@      @      ?@      �?      �?      @       @     �C@      0@              3@     �c@      $@      ;@      5@     @S@     `w@      ,@     x�@      @       @      M@      A@     P}@     �q@      ,@     @d@      �?      @      �?              @      ,@              :@                              �?     �@@      &@               @      �?                               @      @              0@                              �?      5@      @              �?              @      �?              �?      &@              $@                                      (@      @              �?     �B@      "@       @       @      1@      a@      @      l@      @      �?      &@      &@     �d@     �c@      @     �G@     �@@       @      @       @      .@     @Z@      @     �b@      @      �?      &@      "@     @_@     �_@      @     �D@      5@              @              @     @P@      @     �O@      @               @      @      H@     �I@      @      6@      (@       @               @      "@      D@      �?      V@      @      �?      "@      @     @S@     �R@      �?      3@      @      @      �?               @      @@      �?     @R@                               @      E@      >@       @      @      @      @      �?              �?      =@             �J@                               @      B@      :@       @      @              @                      �?      @      �?      4@                                      @      @              �?      1@      @      @       @      $@     @P@       @     @d@      @              $@      @      T@      ;@      @      2@      1@      @      @       @      $@     �N@       @     �_@      @              $@      @      Q@      ;@      @      2@      $@      @      @       @      �?      B@             �L@                      "@       @      9@      0@      �?      "@      "@      @      @       @      �?      6@             �G@                      "@       @      5@      (@      �?      "@      �?                                      ,@              $@                                      @      @                      @      �?                      "@      9@       @     �Q@      @              �?      �?     �E@      &@       @      "@       @      �?                      @      &@      �?      C@      �?              �?      �?      A@      @       @       @      @                               @      ,@      �?      @@      @                              "@      @              �?                                              @             �A@                              �?      (@                                                                       @              >@                                      @                                                                      �?               @                                      @                                                                      �?              6@                                      �?                                                                       @              @                              �?      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ(.jxhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�a	h[��?�	           ��@       	                    �?CS#��?�           �@                          �=@���y�?#           |�@                           �?��{�*��?           Ȓ@������������������������       �	�8�6��?[            @b@������������������������       �"�W��?�           ��@                          �@@I�7�&��?            �F@������������������������       �4�݃�R�?            �A@������������������������       �ffffff�?             $@
                          �:@.(0׽��?�           `�@                            �?�ln��?C           ��@������������������������       ��ٌ>�?e           x�@������������������������       �Y�=�"��?�            @u@                            �?1�R^|�?�            �n@������������������������       ���FG�?E            @W@������������������������       �$����%�?R             c@                           �?o�*O�?�           H�@                           @l&�&�P�?7           @                          �=@�� i���?�            px@������������������������       ����mr�?�            @w@������������������������       ��8	���?             3@                           �?J+�K��?@            �Z@������������������������       ��EC�?"             M@������������������������       ��q�q\�?             H@                          �;@�Ds�y=�?�           �@                          �9@�x���$�?]           P�@������������������������       �4K��G�?:           }@������������������������       ������?#            �L@                           @��C��?6            �U@������������������������       ���d���?0             S@������������������������       ���!pc�?             &@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      8@      A@      ?@     �[@     ��@      A@     Ԑ@      6@       @     �R@     �P@     p�@     ��@      0@     �q@     �a@      1@      7@      :@     �W@     �}@      9@     �@      3@      @     �P@      M@     P@      y@      ,@     �m@     @P@      @      4@      0@      L@     @m@      *@     �p@      (@      @      7@     �@@     `i@      e@      @     �^@     �O@      @      4@      0@      J@      m@      *@     �n@      (@      @      7@     �@@      i@     �c@      @     @^@       @       @      @       @      @      .@      �?      F@       @              @      @      :@       @              5@     �K@      @      .@      ,@     �G@      k@      (@      i@      $@      @      3@      >@     �e@     �b@      @      Y@       @                              @       @              6@                                       @      (@              �?      �?                              @       @              3@                                               @              �?      �?                                                      @                                       @      @                     �R@      $@      @      $@      C@     @n@      (@     0{@      @      �?     �E@      9@     �r@     @m@      $@     @]@     �Q@      @      @       @      A@     @j@      (@     �u@      @             �D@      2@     @m@     �j@      "@     �X@      G@      @       @      @      ,@     �c@      &@     �q@      @              8@      (@     @g@     �b@       @      O@      9@      �?      �?       @      4@     �I@      �?     �P@      �?              1@      @      H@     �O@      �?     �B@      @      @               @      @      @@              U@      �?      �?       @      @      P@      4@      �?      2@      �?                      �?       @      @              >@      �?              �?      @      ?@      (@              @      @      @              �?       @      9@              K@              �?      �?      @     �@@       @      �?      ,@      I@      @      &@      @      1@     �j@      "@     �w@      @       @      "@      "@      k@     @`@       @     �G@      @@      @       @      �?      "@     �W@      @     �a@       @              @      @     �T@     �R@      �?      ;@      :@      @      @      �?       @     @T@      @      Y@      �?              @      �?     �Q@      L@      �?      8@      4@      @      @      �?       @      T@      @      X@                      @      �?      P@      L@              8@      @                                      �?              @      �?                              @              �?              @      �?       @              �?      ,@      �?     �E@      �?              �?       @      *@      2@              @       @               @              �?      @              >@      �?                              @       @               @      @      �?                               @      �?      *@                      �?       @      @      $@              �?      2@       @      @      @       @     @]@       @      m@      �?       @       @      @     �`@      L@      �?      4@      2@       @      @      @      @      V@       @     `i@                       @      @     @^@     �I@      �?      1@      2@       @      @      @      @     �T@       @     �f@                       @      @      X@      H@      �?      .@                                      �?      @              5@                                      9@      @               @                                      @      =@              >@      �?       @                      *@      @              @                                      @      4@              =@               @                      *@      @              @                                              "@              �?      �?                                                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��KhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @I�,��`�?�	           ��@       	                     �?!̇�}��?           �@                           @l��ˆ�?D           ��@                           @��"N��?�           ��@������������������������       ��i߳-��?�           �@������������������������       ��2Tv��?             >@                            �?yv6Lm��?^           h�@������������������������       ��&bf�n�?�            �l@������������������������       ���ɲ�}�?�            �t@
                           �?�(9<R��?�           ؅@                           �?PS!����?I             Z@������������������������       �؍����?!            �F@������������������������       �J������?(            �M@                           @U8;X`��?w           ��@������������������������       ��qĀu��?N           ��@������������������������       ���<S%�?)            @P@                           �?ߧ��g�?�           ��@                           �?a�ʎ2�?�            �r@                           �?#G�h��?y             g@������������������������       �UUUUU��?             H@������������������������       �|�l�]�?Z             a@                          �1@���+���?S            �]@������������������������       �9��8���?             8@������������������������       �/M�EG��?A            �W@                           �?R����?�           ��@                          �6@P�%�W�?             �J@������������������������       �     ��?             0@������������������������       ��d��3��?            �B@                           �?���r$�?�           ��@������������������������       ����	��?�            �q@������������������������       �T�s�	�?           �{@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@     �B@     �G@      :@     �\@     (�@     �D@     ��@      .@      @      T@      N@     ��@     �@      :@     �l@     @c@      :@      A@      :@     @W@     �}@     �A@     ��@      $@      @     �Q@      K@     �}@     �x@      9@      h@     �[@      7@      9@      4@      O@     x@      <@     h�@      @      �?     �F@      >@     �u@     �q@      "@      `@     �U@      4@      6@      *@     �D@     @r@      7@     �z@      @             �B@      9@      p@      l@      @     @W@     �T@      2@      6@      *@      D@     @r@      2@     �z@      @             �B@      9@     p@      k@      @      V@      @       @                      �?              @      @                                      �?       @              @      8@      @      @      @      5@     @W@      @      h@      @      �?       @      @      W@     �L@      @     �A@       @       @              @      @      A@       @      X@                       @      @      C@      1@      @      &@      0@      �?      @      @      ,@     �M@      @     @X@      @      �?      @       @      K@      D@      �?      8@     �E@      @      "@      @      ?@     �W@      @      a@      @      @      9@      8@     �^@      \@      0@      P@      @      �?      �?       @       @      4@      �?      1@      �?              @      �?      *@      "@      @      1@       @                       @      @      @              @      �?              @               @      @       @      "@      �?      �?      �?              @      0@      �?      ,@                      �?      �?      @      @      @       @      D@       @       @      @      7@     �R@      @     �]@       @      @      4@      7@     �[@     �Y@      &@     �G@      D@       @      @      @      7@     @Q@      @     �W@      �?      @      1@      7@      X@      V@      &@     �F@                      �?                      @              8@      �?              @              ,@      .@               @      G@      &@      *@              5@     �d@      @      {@      @              $@      @     �k@     �[@      �?     �B@      .@       @       @              @      E@      @     �Y@                      @      �?     �R@      >@              4@      @               @               @      :@       @      Q@                       @             �E@      4@              0@                                              "@              .@                                      &@       @              @      @               @               @      1@       @     �J@                       @              @@      (@              &@      (@       @                      @      0@      �?      A@                       @      �?      @@      $@              @      @                                      @              (@                                      @       @                       @       @                      @      *@      �?      6@                       @      �?      =@       @              @      ?@      "@      &@              .@      _@      @     �t@      @              @      @     �b@      T@      �?      1@       @              @                      @              @@      �?                               @      @              �?       @              @                      @              @                                      �?      �?              �?                      @                       @              ;@      �?                              �?      @                      =@      "@      @              .@     �]@      @     �r@      @              @      @     @b@      S@      �?      0@      3@      @      @              $@     �G@       @      Y@      �?               @       @     �G@     �B@      �?      @      $@       @       @              @      R@      �?     �h@      @              @      @     �X@     �C@              "@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��OhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @��6P��?�	           ��@       	                     �?X���'��?�           ,�@                          �:@�ft<=��?�           ,�@                           @�����?           ��@������������������������       �3�x�$��?           X�@������������������������       �)\���(�?             4@                           @O�mL�?i            �e@������������������������       �R�I1-��?Z            �b@������������������������       �;n,�R�?             6@
                            �?�;	[u�?Y           ,�@                          �4@��P�1�?�           ��@������������������������       �Vo#��?S           ��@������������������������       ��vR)�?Z           x�@                           @u�)F+��?�           X�@������������������������       ��c�M���?�            �r@������������������������       ���ڣʳ�?�            �w@                           @�&����?�           ̐@                          �;@v��j��?n           ȍ@                           @7�O� �?$           ��@������������������������       ��8�Hs��?_           @�@������������������������       ���(�2Y�?�            �r@                           @J��3n�?J            @Z@������������������������       ���*��?(            �K@������������������������       ��HP��?"             I@                           �?a㟌�V�?N            �^@                           @
�%����?/             R@������������������������       ��b�=y�?              I@������������������������       ��!pc��?             6@                           �?��ڊ�e�?             I@������������������������       ��(\����?             $@������������������������       ��������?             D@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      :@      =@      0@      Z@     �@      4@     ��@      *@       @     �V@     �O@     P�@     (�@      6@     �p@     �c@      0@      7@      .@     �T@      ~@      1@     0�@      *@      @      S@     �L@     �@     �z@      4@     @l@      E@      @      �?      @      3@      h@      @      t@       @              .@      1@     @i@      b@      @     �K@     �D@      @      �?      @      (@     �e@       @      p@       @              ,@      0@     �c@     ``@      @     �B@     �A@      @      �?      @      &@     �d@       @     �o@       @              ,@      0@     �c@     ``@      @     �B@      @       @                      �?      @               @                                       @                              �?                              @      3@      @     �P@                      �?      �?     �E@      *@              2@      �?                              @      2@      @      J@                      �?      �?     �C@      $@              2@                                              �?              ,@                                      @      @                     @]@      &@      6@      "@      P@     �q@      (@     @x@      &@      @     �N@      D@     @s@     �q@      *@     `e@      Q@      @      .@      @     �@@     @h@      @     @p@      @       @     �@@      8@     @i@     `c@      @     �Y@      D@       @      @      �?      4@     �[@      @     ``@       @       @      3@      (@     �W@      U@      @      ;@      <@      @      "@      @      *@     �T@      @      `@      @              ,@      (@     �Z@     �Q@              S@     �H@      @      @       @      ?@     @W@      @      `@      @      @      <@      0@     �Z@      `@       @      Q@      0@      @      @      �?      .@     �B@              H@       @      @      (@      �?     �J@      O@      @      B@     �@@       @       @      �?      0@      L@      @      T@       @              0@      .@     �J@     �P@      @      @@     �G@      $@      @      �?      5@     �g@      @     �w@               @      ,@      @     �m@     �^@       @     �C@      F@      "@      @      �?      0@      d@       @     pu@               @      (@      @     �i@     �[@       @     �@@      B@      "@      @      �?      (@      a@       @     Pr@              �?      (@      @     �h@     �Z@      �?      >@      7@      @      @      �?      $@     �R@      �?     �h@                      $@      �?      b@     �N@              4@      *@      @                       @      O@      �?      X@              �?       @      @      J@      G@      �?      $@       @                              @      9@              I@              �?              �?       @      @      �?      @       @                              @      ,@              5@              �?              �?      @      @              @      @                                      &@              =@                                      @              �?              @      �?                      @      <@      �?      A@                       @              ?@      &@              @              �?                      @      3@      �?      ,@                       @              2@      "@              @                                      @      1@               @                      �?              *@      @                              �?                      �?       @      �?      @                      �?              @       @              @      @                                      "@              4@                                      *@       @              @       @                                      @               @                                      �?                       @      �?                                      @              2@                                      (@       @              �?�t�bub�     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�c%hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @2�
e��?�	           ��@       	                     �?0���?            �@                           @�������?�           �@                          �?@ɕ�+�?           8�@������������������������       ��p�(�I�?�           X�@������������������������       �T�r
^N�?             <@                          �2@$�.�@�?�            `k@������������������������       ���/��@�?-            @Q@������������������������       �������?_            �b@
                          �1@W�2��?s           8�@                           �?�@!����?�             t@������������������������       �V�R����?u            �e@������������������������       �e��}`\�?T            �b@                           �?h	�[�?�           0�@������������������������       ����]� �?�             j@������������������������       �^EW~S�?*           �@                           �?<vo���?�           �@                          �<@��Y��1�?.           �}@                          �5@]ۡ�u&�?           �z@������������������������       ��<�A��?�            pp@������������������������       ��<G` �?g             d@������������������������       ��):���?             I@                          �2@rE�h��?�           ��@                           @>`p��0�?Y             a@������������������������       ��/��C�?P            @_@������������������������       ��q�q�?	             (@                           @� �� r�?1           `}@������������������������       �N�]���?�             q@������������������������       �p�eW~C�?�            �h@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@     �A@      C@      =@      \@     ��@      @@     H�@      3@      @      W@     @R@     �@     ��@      2@     �p@     `b@      :@      A@      8@     �V@     `|@      ;@     `�@      0@      @     �R@     �O@      �@     @y@      0@     `k@     �@@      $@      @      $@      4@     �d@      0@     �s@      @              2@      1@      j@     �a@      "@      G@      ;@      $@      @      @      *@      a@      .@     �m@      @              0@      ,@      e@     @\@      @     �B@      ;@      $@      @      @      *@      a@      .@     @k@      @              0@      *@     �d@      [@      @      B@                                                              2@                              �?      @      @              �?      @                      @      @      ?@      �?     �T@      �?               @      @      D@      <@      @      "@      @                      �?       @      1@      �?      3@                      �?       @      @      $@              @      @                       @      @      ,@              P@      �?              �?      �?     �@@      2@      @      @     �\@      0@      ;@      ,@     �Q@     �q@      &@     �x@      (@      @     �L@      G@     0s@     pp@      @     �e@      6@      �?      @      �?      "@      K@      @      D@      @      �?      0@      (@     �J@      R@              >@      3@              @              "@      <@      @      1@      @      �?      @      @      >@      =@              6@      @      �?              �?              :@              7@                      &@      "@      7@     �E@               @      W@      .@      6@      *@      O@      m@       @     Pv@      "@      @     �D@      A@     �o@     �g@      @     �a@      (@       @      @       @      $@      7@             �G@      @              @      "@     �J@      4@      @      0@      T@      *@      2@      &@      J@     @j@       @     `s@      @      @     �B@      9@      i@     `e@      @     �_@      E@      "@      @      @      5@     �e@      @     `x@      @       @      1@      $@     �k@     @`@       @     �F@      8@      @       @      @      *@     �R@      @     �a@      @      �?      *@      @     �W@      P@              ;@      .@      @       @      @      (@     @R@      @     �^@      �?      �?      *@      @     �V@      L@              8@       @       @              @      &@      B@       @     �U@              �?      "@      @      J@      ?@              1@      @      �?       @              �?     �B@       @      B@      �?              @              C@      9@              @      "@                              �?      �?              4@       @                      �?      @       @              @      2@      @       @       @       @     @Y@      �?     �n@              �?      @      @     �_@     �P@       @      2@      @                      �?      @      7@              C@                              �?     �H@      (@              @      @                      �?      @      6@              >@                              �?     �G@      &@              @                                              �?               @                                       @      �?                      ,@      @       @      �?      @     �S@      �?      j@              �?      @      @     @S@      K@       @      (@      @      �?       @      �?      @     �A@             �`@              �?      @       @      E@      ?@               @      @      @                             �E@      �?      S@                               @     �A@      7@       @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��6hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B(                             !@�}��Ϝ�?�	           ��@       	                    @$��i��?�	           N�@                           �?[b\?�Y�?c           �@                           �?����q�?�           h�@������������������������       �ƽ�-��?}           ��@������������������������       ��������?k           (�@                           �?�9Ձ�!�?{           p�@������������������������       �W���g�?           p|@������������������������       ���l&���?^           8�@
                            @�rs���?:           |�@                           @n����3�?�           �@������������������������       ��� J�?p           ��@������������������������       �t���i�??            @W@                           @B���%%�?�            �l@������������������������       �G{����?:            �W@������������������������       ��Ҿ�6�?Q            �`@                           @�*�u��?             A@������������������������       ��˹�m��?	             3@������������������������       �؂-؂-�?             .@�t�bh�h4h7K ��h9��R�(KKKK��h��B�	       @l@      A@     �E@      8@     �Y@     ��@      :@     ��@      3@      @      S@      L@     ؇@     ��@      8@     �o@     @l@      A@     �E@      8@      Y@     @�@      7@     ��@      3@      @      S@      L@     ؇@     ��@      8@      o@     `b@      3@      :@      *@      N@     `{@      ,@      �@       @      @      I@      ?@     X�@     �u@      1@      a@     �U@      ,@      6@      &@      C@      o@       @     �{@      @      @      @@      4@     �s@     `i@      "@      X@     �C@      @      2@       @      5@     @[@      �?      e@      @       @      5@       @     �Y@      T@      @      F@      H@      "@      @      "@      1@     �a@      @     pq@      @      �?      &@      (@     �j@     �^@      @      J@      N@      @      @       @      6@     �g@      @     p@      �?      �?      2@      &@     �m@     �a@       @      D@      A@      @               @      *@     �W@      @     �\@      �?              @       @     @W@      O@      @      5@      :@       @      @              "@     �W@      �?     �a@              �?      &@      "@     @b@     @T@      @      3@     �S@      .@      1@      &@      D@     @j@      "@     @v@      &@      �?      :@      9@      j@      g@      @      \@      R@      &@      ,@      $@     �B@     �d@      @     q@      @      �?      5@      6@     �d@     @d@      @      [@     �Q@      &@      &@      $@      B@     �c@      @      n@      @      �?      2@      3@      c@     �a@      @     �Y@      �?              @              �?      "@      �?     �@@      �?              @      @      (@      4@              @      @      @      @      �?      @     �E@       @     �T@      @              @      @      F@      6@              @      �?       @                      �?      @              H@                      @              7@      @               @      @       @      @      �?       @      B@       @     �A@      @              �?      @      5@      .@               @                                       @      0@      @       @                                              @              @                                              &@               @                                              @              �?                                       @      @      @                                                      �?              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJx�EhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @KC2ylt�?�	           ��@       	                    �?=�	���?�           �@                          �1@lvk.p�?           ��@                           @Ktuc���?�            �o@������������������������       �d���1��?p            @g@������������������������       �o(T���?+            �P@                           @.
�&�?u           P�@������������������������       �%�׫��?m           ��@������������������������       �s
^N���?             ,@
                          �;@8��S�.�?�           0�@                            �?#�O�?Y           ��@������������������������       �k	
���?�           �@������������������������       ��r5�O��?�            �s@                           @�J{��?x            �i@������������������������       �w^�����?\            @d@������������������������       �`Ӹ����?            �F@                           @����O�?�           \�@                           �?6+�Ҽ/�?           �@                           @���F�{�?�            �w@������������������������       �0i?��Q�?�            �t@������������������������       �t�!~���?!            �E@                           �?1&[ץ��?           �|@������������������������       ��,V����?Z             a@������������������������       �R���)�?�             t@                           �?�S���?�            @q@                           @��P�??            �[@������������������������       �DzA��d�?6            �W@������������������������       ��������?	             1@                           �?���5�?d            �d@������������������������       ��q�q�?             8@������������������������       ��.Pe���?S            �a@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      C@     �B@      2@     �W@     ��@      C@     ��@      <@      "@     @V@      P@     ��@     �@      4@     �m@     �a@      <@      ;@      $@     �T@     p}@      @@     H�@      4@      @     �R@      H@     8�@     �w@      2@     �h@      R@      *@      3@      @     �H@     �l@      ,@     Pq@      *@      @     �@@      :@     �j@      d@      "@     @\@      &@      @      @              @      B@      "@      @@      @      @      @      $@      G@      H@       @     �@@      $@      @       @               @      2@       @      6@      �?              @      $@      E@     �A@       @      :@      �?              @              �?      2@      �?      $@       @      @      �?              @      *@              @     �N@      $@      (@      @      G@     @h@      @     �n@      $@      @      ;@      0@      e@      \@      @      T@     �N@      $@      (@      @     �E@     @h@      @     `n@      $@      @      ;@      0@     �d@      [@      @     �S@                                      @               @       @                                      �?      @               @      Q@      .@       @      @     �@@      n@      2@     @}@      @      �?      E@      6@     s@     �k@      "@      U@     �O@      ,@       @      @      @@     @j@      0@     @x@      @      �?     �A@      1@     Pp@     �j@      @     �Q@      F@      $@      @      @      2@     �e@      (@     �t@      @              5@      (@     �i@     @b@      �?     �F@      3@      @      @              ,@     �B@      @      N@      @      �?      ,@      @     �K@     �P@      @      :@      @      �?              �?      �?      ?@       @      T@      �?              @      @      F@      &@      @      *@      @      �?                      �?      1@       @     �P@      �?              @      @      <@      &@      @      *@                              �?              ,@              ,@                                      0@                             �H@      $@      $@       @      *@     �g@      @     �w@       @       @      ,@      0@     �m@     �_@       @      D@      D@      @      $@       @      (@     �]@      @     0r@      @              &@       @     �h@     �V@       @      A@      <@      @      @              $@     �Q@      �?     �W@       @               @      @     �U@      F@       @      3@      9@      @      @              "@     �N@      �?     @V@       @              @      @     �S@      A@       @      .@      @              �?              �?      "@              @                      �?               @      $@              @      (@      �?      @       @       @      H@      @     �h@      �?              @      @     �[@      G@              .@                               @              *@              J@                       @       @      B@      7@              @      (@      �?      @      @       @     �A@      @      b@      �?              �?      @     �R@      7@               @      "@      @                      �?     �Q@             �V@      @       @      @       @      D@     �B@              @      @      �?                              5@              A@       @       @      @      @      1@      1@               @      @      �?                              4@              8@       @       @              @      ,@      1@               @                                              �?              $@                      @              @                               @      @                      �?     �H@             �L@      @                      @      7@      4@              @      �?                              �?      @              @                                      @       @                      �?      @                             �E@              J@      @                      @      4@      (@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��4IhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B(                             !@6,|�.w�?�	           ��@       	                    @��qt�?�	           Z�@                            @ڴ��P�?C           @�@                          �0@,��¾��?           t�@������������������������       ���(W�?.             U@������������������������       ��u%@��?�           $�@                          �;@��ǎ�?0           �@������������������������       �l<�>�H�?�           ��@������������������������       ���f���?N            �`@
                            @}�f:��?E           4�@                          �;@��)a��?�           ̐@������������������������       �n�5�.�?�           8�@������������������������       �?�ƨ�?.             S@                          �0@$^�7a�?�            @k@������������������������       �Er���&�?             1@������������������������       ��Qje�A�?~             i@                            �?*x9/��?             <@������������������������       �����>4�?
             ,@������������������������       �������?             ,@�t�bh�h4h7K ��h9��R�(KKKK��h��B�	       �j@     �C@     �B@      9@     @X@     ��@      ?@     ��@      .@      $@     @W@      M@     H�@     `~@      1@      o@     �j@     �C@     �B@      9@     �W@     ��@      =@     ��@      .@      $@     @W@      M@     @�@     0~@      1@     �n@     `a@      9@      9@      ,@      L@     �{@      1@      �@      @      @      O@      ;@     8�@     `v@      @     `b@      W@      6@      ,@      (@     �C@     �r@      ,@     @z@       @       @     �L@      .@     0t@     p@      @     @^@                       @              @      .@       @      "@                              @      7@      2@              @      W@      6@      (@      (@      B@     �q@      (@     �y@       @       @     �L@      "@     �r@     �m@      @     �\@     �G@      @      &@       @      1@     `b@      @      t@      @      @      @      (@     �h@     @Y@      �?      :@      B@      @      &@       @      (@     �_@      @     p@      @      @      @      (@     �e@     @W@              9@      &@                              @      4@             �O@              �?                      7@       @      �?      �?     �R@      ,@      (@      &@     �C@     �j@      (@     x@      $@      @      ?@      ?@      l@     @_@      &@     @X@      R@      "@      "@       @     �@@     �f@      &@     �r@       @      @      =@      ?@     `f@     �Z@      &@     �U@      P@      "@      "@       @     �@@     �e@      &@     `p@       @      @      =@      =@      d@     �Y@      &@     @U@       @                                      @             �A@                               @      2@      @               @      @      @      @      @      @      >@      �?      V@       @               @              G@      3@              $@                                                      �?      @                                      "@      @                      @      @      @      @      @      >@              U@       @               @             �B@      0@              $@                                       @      &@       @      @                                      �?      @              @                                       @      @       @      �?                                      �?      �?                                                              @              @                                               @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�W
hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@���0M��?�	           ��@       	                     @W/����?�           X�@                          �0@d�%�"�?C           ��@                           @Ʒ?�?d            �b@������������������������       ��k�{�9�?[            �`@������������������������       �      �?	             0@                           @'�x6�?�           t�@������������������������       �t�u�%��?�           ��@������������������������       ��<�:�*�?9           P�@
                           �?c��6y�?b           ؎@                          �6@�h[�D#�?
           �z@������������������������       �����?�            s@������������������������       �l���?L            �]@                          �2@Sep����?X           ��@������������������������       ��qDQ`*�?l            �f@������������������������       �x~�q%�?�            �w@                           @��d��M�?           �y@                           @ǘb����?�            �v@                           @�B����?�            Pq@������������������������       �t��A��?K            @]@������������������������       �H�z�G�?k             d@                           @/��	�?<            �U@������������������������       ���=A��?             C@������������������������       �9��8�#�?              H@                           �?/�$���?"             I@������������������������       �X�<ݚ�?             "@                           �?��01m��?            �D@������������������������       �r`�����?             3@������������������������       �x?r����?             6@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        l@      ;@     �J@      4@     �W@     �@      A@     А@      1@      $@     �U@     �P@     Ї@     �@      6@     �p@     �i@      4@      I@      4@     �U@     ��@      @@     Ȍ@      &@       @      S@      O@     ؅@     �}@      2@     `n@     �d@      ,@     �C@      0@     �Q@     �y@      8@     Ђ@       @       @     �N@      K@     P}@     �v@      1@     �h@      (@              @              "@      >@      �?      .@              �?              @      ?@      @@              (@      (@              @              @      9@      �?      ,@              �?              @      >@      9@              (@                                       @      @              �?                                      �?      @                      c@      ,@      A@      0@      O@     �w@      7@     X�@       @      @     �N@     �I@     `{@     �t@      1@      g@     �U@      @      5@      $@      =@      d@      @     �q@       @      @      4@      8@      k@     �^@      @      Q@     @P@      $@      *@      @     �@@     `k@      0@      s@      @      @     �D@      ;@     �k@     �i@      $@      ]@     �E@      @      &@      @      .@     �c@       @     �s@      @              .@       @     �l@     �]@      �?     �G@      6@      @      @      �?      "@     @T@      @     @]@                      &@              W@      L@              1@      3@       @      �?      �?      "@      H@      @      W@                      "@              P@      C@              1@      @      @      @                     �@@      �?      9@                       @              <@      2@                      5@              @      @      @     �S@       @     @i@      @              @       @     @a@      O@      �?      >@      @              �?      @       @      4@              G@                      �?      @      M@      ?@              $@      1@              @              @      M@       @     �c@      @              @      @      T@      ?@      �?      4@      1@      @      @              "@     �R@       @     `c@      @       @      &@      @     �O@      @@      @      8@      1@      @      @              "@      P@       @     �_@      @       @      "@      @      K@      @@      @      8@      "@      @       @              @     �I@       @     �Y@      @       @      "@      �?     �@@      :@      @      3@      @      @       @              @      <@      �?     �A@      @       @      @      �?      &@      @      �?      @      @       @                              7@      �?     �P@                      @              6@      6@      @      (@       @              �?               @      *@              9@      @                       @      5@      @              @      @              �?                      @              2@                               @      @                       @      @                               @      "@              @      @                              .@      @              @                                              $@              <@                       @      �?      "@                                                                      @               @                                      �?                                                                      @              :@                       @      �?       @                                                                      @               @                       @      �?      @                                                                      �?              2@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ{uhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @Y�-E���?�	           ��@       	                    @�(G%��?�           �@                          �0@�c/��?;           �@                           @R�����?^             d@������������������������       �ҤI�&M�?+            @R@������������������������       ��mI���?3            �U@                           @(��Q��?�           ��@������������������������       ��U�����?           D�@������������������������       ��*.jI�?�           0�@
                           !@    �o�?�             p@                          �;@(�He���?�            `n@������������������������       ����ք��?�            �h@������������������������       �x��J�?             G@������������������������       ��s�n_�?	             *@                           �?���VL�?�           H�@                           @R�
�@_�?�           ��@                          �4@<��^�?�           ��@������������������������       �
 �����?�             n@������������������������       ���F��?           @z@������������������������       �{�G�z�?             $@                           @πKl�?#           0{@                          �2@lzW&���?�            �t@������������������������       ��Z�J��?H            �[@������������������������       �"�K"z��?�            �k@                          �5@b������?I            @Y@������������������������       ��ѳ�w�?$            �I@������������������������       ���3���?%             I@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        j@      9@      >@      8@     @]@     h�@      <@     p�@      7@       @     �U@     �R@     ��@     �@      8@     Pp@      d@      4@      6@      6@     @W@      {@      8@     �@      0@      @     @S@      P@     ��@     �v@      5@      k@     �c@      4@      4@      6@     �U@     Py@      0@     �@      *@      @      Q@     �N@     �~@     �t@      5@     �g@      @      �?      �?       @      "@      >@              ,@      @      @      @      (@      =@      ?@       @      &@       @                              @      $@              @                              (@      0@      4@       @      @       @      �?      �?       @      @      4@              $@      @      @      @              *@      &@              @     `c@      3@      3@      4@     �S@     pw@      0@     ��@      $@       @     �N@     �H@     �|@     �r@      3@     �f@     �Z@      .@      (@      (@      E@     �q@      (@     @|@      @      �?     �F@      >@     �t@      k@      .@     @Z@      H@      @      @       @      B@     @W@      @      f@      @      �?      0@      3@     �`@     @T@      @     �R@      �?               @              @      ;@       @     �W@      @              "@      @     �D@     �B@              9@      �?               @              @      8@      @     �W@      @              "@      @      D@     �A@              8@      �?               @              @      3@      @     �P@      @               @       @      >@      A@              7@                                              @              ;@                      �?      �?      $@      �?              �?                                       @      @      @                                              �?       @              �?      H@      @       @       @      8@     �g@      @     �w@      @       @      $@      &@     @l@     �a@      @     �F@     �B@       @      @       @      *@      \@      �?     �m@      @       @      @      "@      ]@      W@      @      >@     �B@       @      @       @      *@      [@      �?     `m@      @       @      @      "@      \@      W@      @      >@      1@              @       @      @      8@             @S@      @              @       @     �D@     �G@              .@      4@       @      @               @      U@      �?     �c@      �?       @              @     �Q@     �F@      @      .@                                              @               @                                      @                              &@      @       @              &@     @S@      @     �a@      �?              @       @     �[@     �I@              .@       @       @       @              &@     �J@       @     �]@                      @             @U@      B@              (@      �?                               @      6@              >@                                      D@      (@              @      @       @       @              "@      ?@       @      V@                      @             �F@      8@               @      @      �?                              8@      �?      8@      �?               @       @      9@      .@              @      @      �?                              @      �?      *@                       @       @      1@      @               @                                              3@              &@      �?                               @      $@              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ؜*BhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @N7�����?�	           ��@       	                   �:@�p�CQ=�?�           ҥ@                           �?� ���K�?�           �@                          �4@80ј)��?�           ��@������������������������       ���ѡ��?�           ��@������������������������       ���a��?!           P|@                          �0@_~$���?>           ܔ@������������������������       ��.�袋�?4             V@������������������������       ��ʇ ��?
           |�@
                            �?B>=܂y�?�            Pw@                           @�.�@���?f            �c@������������������������       �V�F�?�?U            @_@������������������������       ���paR�?             A@                           @ߛm�
��?�            �j@������������������������       �n۶m���?I             \@������������������������       �ݑF��d�??            �Y@                           �?�h3��3�?�           ��@                           @r����?>           �@                          �2@D	�c��?�            �u@������������������������       ��/�<n�?;            �V@������������������������       ��tx<��?�            @p@                          �6@PY�����?b            �c@������������������������       �(vb'vb�??             Z@������������������������       ��U}��`�?#            �K@                           @�����?�           �@                           @� i����?$           �|@������������������������       �r��/ �?           py@������������������������       �U���N@�?             I@                           @���u�?c            @c@������������������������       �Mb�R>�?Y            �a@������������������������       �������?
             *@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      B@      J@      3@      ^@     ؃@      =@     ��@      2@      @     @Y@      O@     `�@     ��@      2@     Pr@     `d@      ;@      E@      0@     �X@      |@      :@     `�@      ,@      @     �V@     �K@      ~@     �x@      0@     �m@      b@      5@      A@      0@     �T@      y@      7@     ��@      &@      @     �R@      I@     �y@     �v@      .@     �i@     �N@      *@      7@      @     �F@     `i@      "@      i@      "@       @      >@      ?@     �f@     @c@      "@     @[@     �H@      (@      3@       @      :@     �Y@      @     �\@      @       @      .@      4@     @V@     �Z@      @     �L@      (@      �?      @      @      3@      Y@      @     �U@      @              .@      &@     �V@      H@       @      J@     �T@       @      &@      $@      C@     �h@      ,@     �v@       @      �?      F@      3@      m@     �i@      @     �X@      "@                      �?              1@              ,@                      @      @      (@      .@              "@     �R@       @      &@      "@      C@     �f@      ,@     �u@       @      �?     �C@      *@     �k@      h@      @     @V@      3@      @       @              0@      G@      @      ^@      @      �?      0@      @      Q@      @@      �?      =@                                      "@      .@       @     @Q@       @              @      �?     �A@      $@              &@                                      "@      *@       @      K@       @              @      �?      4@       @              &@                                               @              .@                                      .@       @                      3@      @       @              @      ?@      �?     �I@      �?      �?      &@      @     �@@      6@      �?      2@      0@      @       @              @      ,@              ,@      �?              @      @      :@       @      �?      @      @                                      1@      �?     �B@              �?       @      �?      @      ,@              *@     �E@      "@      $@      @      5@     `g@      @     @x@      @              &@      @     �m@     `a@       @     �L@      ;@      @       @              *@     �V@      @      _@      @              "@      @      \@      S@      �?      A@      ,@      @      @               @     �Q@       @     �Q@       @              "@       @      U@      L@              9@                                      @      4@              *@                              �?      A@      $@              "@      ,@      @      @              @      I@       @     �L@       @              "@      �?      I@      G@              0@      *@      �?      @              @      5@      �?      K@       @                      �?      <@      4@      �?      "@      @                              @      (@              E@                              �?      4@      *@               @      "@      �?      @              �?      "@      �?      (@       @                               @      @      �?      �?      0@      @       @      @       @      X@             �p@                       @      @      _@     �O@      �?      7@      ,@      �?       @      @       @     �K@             �j@                       @      @      Y@      D@              0@      $@      �?       @      @       @      F@             �f@                       @      @      X@     �C@              .@      @                                      &@              =@                                      @      �?              �?       @      @                             �D@              J@                                      8@      7@      �?      @       @      �?                              B@              I@                                      6@      6@      �?      @              @                              @               @                                       @      �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJu	&hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@�U�:5��?�	           ��@       	                     @�x�3���?�           �@                           �?$=�G�??           ��@                            �?�7��~�?�           ��@������������������������       �nL�"�?           �@������������������������       ���);� �?�            `r@                           @JS+\��?�           ܕ@������������������������       ��!Ñ��?n           l�@������������������������       �����X�?             <@
                           �?�
�:~�?Y           h�@                           @���x��?           �z@������������������������       �U����)�?�            �q@������������������������       �h{�U�?R            �b@                           �?    �V�?Q            �@������������������������       �G��o>8�?L            �_@������������������������       ��-]
�?            x@                           @>�\��p�?            |@                            @�y �c�?�            `w@                          �@@Zos=��?�            `m@������������������������       �0���?�             k@������������������������       �J�w�"w�?             3@                          @@@8�E��?T            `a@������������������������       ������?C            @Z@������������������������       �}�@�m�?             A@                          �?@����k�?0             S@                           �?7��o�?)            @P@������������������������       ��
t�F��?             1@������������������������       ��q�q��?             H@������������������������       ���ˠ�?             &@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@     �B@     �D@      9@     �Z@     ��@      C@     |�@      8@      0@     �R@      P@     (�@     Ѐ@      3@      q@     �f@      =@      D@      8@     @Y@     x�@      B@     ȍ@      8@       @     �O@      N@     Ѓ@     @      &@     `n@      b@      5@      ?@      5@     �S@     �y@      7@     ؃@      1@      @      L@      I@     �{@     �v@      &@      j@     �N@      "@      ;@      "@      H@     `j@      ,@     �n@      0@       @      4@      :@     �e@     �b@      @     @Y@     �H@      @      1@      @     �@@      d@      *@     �i@      @              *@      2@     �`@     @X@      @     �P@      (@      @      $@      @      .@     �I@      �?      D@      "@       @      @       @      E@      K@       @     �A@     �T@      (@      @      (@      >@      i@      "@     @x@      �?      @      B@      8@     �p@     �j@      @     �Z@     �R@      $@      @      (@      =@      i@      "@      x@      �?      @      B@      8@     �p@     �i@      @      Z@       @       @                      �?      �?               @                                      @      @              @     �B@       @      "@      @      7@     `b@      *@     �s@      @      �?      @      $@     �g@     �`@             �A@      0@      @      @      �?      .@     @Q@       @     �\@      @      �?      @      @     �U@      R@              4@      *@      �?      @      �?      $@     �I@      @     @Q@                      @      �?     �Q@     �C@              (@      @      @      �?              @      2@      @     �F@      @      �?              @      0@     �@@               @      5@       @       @       @       @     �S@      @     �i@       @              @      @     �Y@      O@              .@      �?                                      ,@             �D@                       @      �?      C@      6@              @      4@       @       @       @       @      P@      @     `d@       @              �?      @      P@      D@               @      4@       @      �?      �?      @     �Q@       @     �d@               @      &@      @     �R@     �D@       @      =@      .@       @      �?              @      K@       @      b@               @      &@      @      J@     �A@       @      ;@      "@       @      �?              @      B@       @      U@                      &@      @      9@      7@      @      8@       @       @      �?              @      >@       @     @T@                      &@       @      8@      1@      @      7@      �?                                      @              @                              �?      �?      @              �?      @                               @      2@              N@               @              �?      ;@      (@       @      @      @                              �?      2@              E@                              �?      6@      (@       @      @       @                              �?                      2@               @                      @                              @                      �?              1@              6@                                      7@      @               @      @                      �?              *@              1@                                      6@      @               @      @                      �?              @              @                                       @      @                      �?                                      $@              (@                                      4@      @               @      �?                                      @              @                                      �?                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��FhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �:@_1�A`�?�	           ��@       	                    @��Z|��?           Щ@                            @��e���?           p�@                           �?��P���?K           D�@������������������������       �J;6C]x�?�           ؉@������������������������       ��FcsG>�?P           ��@                          �2@���D�?�           8�@������������������������       ��M���?�             o@������������������������       �l�����?;           �~@
                           !@n�6����?�           ��@                           @+x�v��?�           ��@������������������������       �BD�����?�           ��@������������������������       �%�jE�P�?B            �[@������������������������       �Iє�?
             1@                            @�4�*��?           �@                           @�������?�            �x@                           @@��f~�?�            �p@������������������������       ����C�y�?�            �k@������������������������       �4և����?            �H@                           �?ִi� �?K            �^@������������������������       ����A�?             G@������������������������       ��!>y��?/            @S@                           @�oGM���?�            �j@                           �?'&��|��?,            �P@������������������������       �����|��?             F@������������������������       �l �&��?             7@                          �?@O�[�?W            �b@������������������������       �N<+	��?F             ^@������������������������       ��Cc}h�?             <@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `f@      @@      E@      ;@     �Z@     ��@      B@     8�@      0@      @     �Q@      P@     H�@      �@      0@     pp@     `c@      6@      A@      :@     @X@     ��@      A@     H�@      *@      @     �N@     �L@     X�@     @      .@     �l@     @^@      *@      9@      8@     �T@     �y@      3@     ��@       @      @      F@     �B@      |@      u@      $@     �f@     @Y@      *@      0@      1@     @P@     �r@      &@     �|@      @      @      @@      @@     pr@     �m@      $@      b@      I@      @      ,@       @     �F@      c@      @     @f@      @       @      0@      1@     �a@     @Z@      @     @S@     �I@      @       @      "@      4@     �b@      @     �q@              �?      0@      .@     `c@     �`@      @     �P@      4@              "@      @      2@     �\@       @     @p@      �?              (@      @      c@     �X@              C@      "@              @      @      @     �B@             �Q@                       @       @      O@      C@              *@      &@              @       @      *@     @S@       @     �g@      �?              $@      @     �V@      N@              9@      A@      "@      "@       @      ,@      ^@      .@      k@      @      �?      1@      4@     `a@      d@      @      H@     �@@      "@      "@       @      &@     �\@      .@     �j@      @      �?      1@      4@     `a@     �c@      @     �G@      >@      @      "@       @      "@     �X@      (@     �f@      @      �?      .@      3@     @]@      b@      @      ?@      @       @                       @      .@      @      @@                       @      �?      6@      *@              0@      �?                              @      @               @                                              @              �?      8@      $@       @      �?      $@     �W@       @     �l@      @              $@      @     �_@     �I@      �?     �@@      0@      @      @      �?       @      L@       @      `@      �?              $@      @     �U@      D@      �?      ;@      .@      @      @      �?      @      D@      �?      R@      �?               @       @     �P@      ;@      �?      3@      $@      @      @      �?      @      @@      �?      L@                       @       @     �M@      .@      �?      3@      @                                       @              0@      �?                              @      (@                      �?                              �?      0@      �?     �L@                       @      @      5@      *@               @                                               @      �?      2@                                      @      @              @      �?                              �?       @             �C@                       @      @      0@      @              �?       @      @      @               @      C@              Y@       @                       @     �C@      &@              @      �?              @               @      @              <@                               @      2@      @              @      �?               @              �?      @              6@                               @      @      @              @                      �?              �?       @              @                                      (@      �?                      @      @                             �@@              R@       @                              5@      @              @      @      @                              ;@             �O@                                      ,@      @              @      @                                      @              "@       @                              @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��uRhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�;c��s�?�	           ��@       	                     �?\�,���?�           �@                          �0@���7���?:           �@                           @��&�'�?O             _@������������������������       �ƯsY�h�?G            �[@������������������������       �*x9/��?             ,@                           �?�;��)y�?�           ��@������������������������       �%�'�*��?�            @u@������������������������       �J��t���?           ��@
                           �?V��2��?�           �@                          �7@�xp�dk�?             �K@������������������������       �T]���b�?            �@@������������������������       ��袋.��?
             6@                           �?�mN����?w           0�@������������������������       �#1��o��?�            �p@������������������������       ��@2�?�            �s@                           �?T�:�{��?�           `�@                           @���h�'�?C           p@                           @�0��	��?�            �t@������������������������       �y�a=Z��?�            �q@������������������������       �dz���2�?            �E@                           @׈2>�?k            �e@������������������������       �C�꫊:�?^            `c@������������������������       �B{	�%��?             2@                          �;@�Ua�	��?�           �@                           @D������?N           �@������������������������       ��
[L�p�?�            `w@������������������������       � �N���?X            �`@                           @���o��?;            �Y@������������������������       ��Mozӛ�?5             W@������������������������       ���!pc�?             &@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@     �@@      C@      4@      \@     ��@      C@     ��@      ,@      *@      P@     @Q@     Ȇ@     P�@      =@      p@     @b@      9@     �@@      4@      W@     �{@      <@     0�@      $@      *@     �K@     �O@     �@     0x@      <@     �i@      ]@      0@      6@      1@     �O@     �v@      4@     Ђ@      @       @     �D@     �F@     @z@     �p@      3@     �a@      @              @      �?      @      ?@      @      "@      �?               @      @      8@      4@              ,@      @              @      �?      @      6@      @      "@      �?                      @      8@      1@              ,@                                              "@                                       @                      @                      \@      0@      3@      0@      M@     �t@      1@     ��@      @       @     �C@      C@     �x@      o@      3@     �_@      6@      �?              �?      1@      B@             �]@      �?              *@      �?     �P@     �C@       @      5@     �V@      .@      3@      .@     �D@     �r@      1@     �}@      @       @      :@     �B@     �t@      j@      1@     �Z@      >@      "@      &@      @      =@     �S@       @     �a@      @      &@      ,@      2@     @V@     �]@      "@      P@      �?       @      @                      @              @       @              @              ,@      @       @      $@               @      @                      �?              @       @              @              @      �?       @       @      �?                                      @              @                                       @      @               @      =@      @      @      @      =@     �R@       @     �`@       @      &@      &@      2@     �R@     �\@      @      K@      .@      @       @      �?      0@     �@@      @      N@       @      @      @      *@      @@     �G@       @      5@      ,@      @      @       @      *@     �D@       @     @R@              @      @      @     �E@      Q@      @     �@@      I@       @      @              4@      g@      $@     �y@      @              "@      @     �k@     �`@      �?     �I@      >@      @      @              ,@     �X@      "@     �b@       @              @       @     @T@     @R@      �?      9@      1@       @      @              &@     @Q@       @     �W@                      @              O@      G@              1@      .@       @      @              "@      K@       @      V@                      @             �L@     �B@              0@       @                               @      .@              @                       @              @      "@              �?      *@      @      �?              @      =@      @      L@       @              �?       @      3@      ;@      �?       @      *@      @      �?               @      6@      @      J@       @              �?       @      0@      8@      �?       @                                      �?      @              @                                      @      @                      4@       @      �?              @     �U@      �?     p@       @               @      @     `a@      O@              :@      4@       @      �?              @     @P@      �?     �h@      �?               @      @     �_@      M@              8@      1@              �?              �?      D@      �?     @c@      �?               @      @     �Y@      @@              3@      @       @                       @      9@             �F@                                      8@      :@              @                                      @      6@              M@      �?                              *@      @               @                                      @      0@              L@                                      &@      @               @                                              @               @      �?                               @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��4hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@�7����?�	           ��@       	                    @<���?�           .�@                           �?�3����?�           �@                          �3@��`s�+�?�           ��@������������������������       ��xQ�`#�?           �|@������������������������       �}�[<�?{           P�@                          �:@���P?��?�           h�@������������������������       �l��NY��?�           ��@������������������������       ��B�f��?"             K@
                            @#w��y��?           ,�@                           !@qFfOK�?G           h�@������������������������       ����j>�?=           ؍@������������������������       � )O��?
             2@                          �2@XV��7�?�            �s@������������������������       �ٗ���N�?,            @Q@������������������������       �zd�Qw�?�             o@                            @��=H���?            {@                           �?����p��?�             s@                            �?�t�����?g             d@������������������������       �j��`5�?/            �P@������������������������       �����?8            �W@                           @  ����?]            �a@������������������������       ���E���?/             R@������������������������       ��[��_�?.            �Q@                          �@@��z��7�?Z            @`@                           �? �Cc=�?O             \@������������������������       �1ogH���?            �@@������������������������       �L�jT���?:            �S@������������������������       ��)O�?             2@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @i@      D@     �A@      6@     �_@     ��@      C@     ��@      0@      $@     �R@      O@      �@     ��@      4@     @n@     �g@      B@      ;@      4@     �]@     ��@     �@@     ��@      $@      $@      Q@      M@     ��@     �~@      2@     `l@      \@      0@      4@      ,@     @U@     �u@      (@     H�@      "@      @     �D@      8@     P~@      q@      *@      b@      M@       @      $@      &@      K@     `f@      "@     �j@      @      @      4@      .@     `k@     �_@      @     @R@      =@      @      @      @      8@     �M@      @     �W@              @      *@      @      \@      P@      @      >@      =@      @      @       @      >@      ^@      @     �]@      @      �?      @       @     �Z@      O@      �?     �E@      K@       @      $@      @      ?@     �d@      @     @w@      @      �?      5@      "@     �p@     �b@       @      R@      J@      @      $@      @      9@     @d@      @     �v@      @      �?      5@      "@      n@      b@       @     �Q@       @       @                      @      @              "@                                      :@      @              �?      S@      4@      @      @     �@@      k@      5@     �t@      �?      @      ;@      A@      j@     `k@      @     �T@      P@      &@      @      @      <@     �d@      3@     �k@      �?       @      8@      =@      c@     �d@      @     �R@      O@      &@      @      @      <@     �c@      *@     �k@      �?       @      8@      =@     �b@     �d@      @     �R@       @                                      @      @                                              �?       @                      (@      "@      �?              @     �I@       @      \@              �?      @      @      L@     �J@      �?      @      @       @                      @      @              .@                      @      �?      0@      1@               @      "@      @      �?                      G@       @     @X@              �?              @      D@      B@      �?      @      ,@      @       @       @       @     @S@      @     �d@      @              @      @     �R@     �D@       @      .@      "@      @      @       @      @     �K@      @     �Y@      @              @      @     �L@      @@      �?      *@      @      @      @              @      A@      @      F@                      @       @      9@      1@      �?      $@       @                              @      $@       @      =@                      �?              @      @              @      @      @      @                      8@      @      .@                      @       @      2@      &@      �?      @      @                       @      �?      5@              M@      @               @      �?      @@      .@              @      �?                              �?      "@              >@                       @              (@      ,@              @      @                       @              (@              <@      @                      �?      4@      �?                      @              �?              @      6@             @P@       @                      �?      2@      "@      �?       @      @              �?              @      6@             �I@       @                      �?      .@      "@      �?       @                                       @      @              $@       @                      �?      @      @              �?      @              �?               @      .@             �D@                                      $@      @      �?      �?      �?                                                      ,@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�� hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B(                             !@|�mΔ�?�	           ��@       	                     @�{ğ,��?�	           `�@                            �?�~���?�           ȥ@                           �?    ���?            �@������������������������       �N��~)�?B           p�@������������������������       ��%p'�"�?�           ȑ@                           @��=����?�            �@������������������������       �Q�n#�?\            �@������������������������       ��d5��?r            �h@
                           �?�;����?�           0�@                           �?��g"���?�            �t@������������������������       �<������?�            `i@������������������������       �����?S            @`@                           �?����a��?�           ��@������������������������       �,i܁���?�            �s@������������������������       ���E���?%            |@                           �?{�G�z�?             9@������������������������       �      �?              @������������������������       �:���I�?
             1@�t�bh�h4h7K ��h9��R�(KKKK��h��B�	        i@     �@@      G@      :@     �[@     ��@     �D@     x�@      9@      @     �S@     �P@     ؆@     �}@      5@     �p@      i@     �@@      G@      :@     �[@     H�@      C@     l�@      9@      @     �S@     �P@     І@     �}@      5@     �p@     @c@      8@      @@      5@     �U@      }@     �@@      �@      3@      @      Q@     �L@     �@     �v@      1@     �l@     @[@      3@      6@      5@      H@     �u@      9@     �@      &@              H@      A@     �w@     �n@      "@     �b@     �F@       @      1@      &@      9@     �e@      @     �k@      "@              =@      2@     �b@     @Z@      @     @T@      P@      &@      @      $@      7@     �e@      2@     �u@       @              3@      0@      m@     �a@      @     @Q@     �F@      @      $@             �C@     @]@       @     ``@       @      @      4@      7@     �^@     �]@       @     �S@     �C@      @      "@              A@     �R@      @      X@      @      @      0@      4@     @X@      R@      @     �N@      @              �?              @      E@       @     �A@      @      �?      @      @      9@     �G@      @      1@      G@      "@      ,@      @      8@     �f@      @     �y@      @              &@      "@      l@     �Z@      @     �D@      &@       @       @       @       @     �M@       @     �\@                      @             @T@     �@@              2@      @               @       @      �?      B@      �?      U@                      @             �B@      3@              ,@      @       @                      �?      7@      �?      >@                      @              F@      ,@              @     �A@      @      (@      @      6@      _@      @     �r@      @              @      "@      b@     �R@      @      7@      5@       @       @      �?      ,@     �M@      @     �Y@       @              �?      @     �M@      ?@       @      "@      ,@      @      @       @       @     @P@             `h@      @              @      @     @U@     �E@       @      ,@      �?                                      ,@      @      @                                      �?      @                      �?                                      @      @                                                      �?                                                              &@              @                                      �?       @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJz�shG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @�v�
�a�?�	           ��@       	                   �;@��ۥ�e�?w           ��@                           �?�L��|�?           Ԙ@                            @��,Ų��?�            �@������������������������       ���"�5��?�            v@������������������������       �S�����?�            0p@                          �2@�0���?z           ��@������������������������       ���-��?�            u@������������������������       �33333]�?�            �@
                          @@@�g����?s             g@                           �?"L�S�?e            �c@������������������������       �G���H�?             5@������������������������       �[{�f��?W             a@                           �?�h�Cד�?             ;@������������������������       �:���I�?             1@������������������������       �ףp=
��?             $@                          �<@��c�RQ�?-           ��@                           �?�w����?�           p�@                           �?"�I&��?�           h�@������������������������       �@!z���?H            �\@������������������������       �Q����	�?�           ؅@                            @PX�hP�?�           ��@������������������������       ���yěq�?�           p�@������������������������       �U"�����?�            v@                           �?�Oy���?q            �g@                           @�Kc�&�?            �B@������������������������       ��G�z��?             4@������������������������       �������?	             1@                           �?CW����?]            @c@������������������������       ���{�~�?             E@������������������������       �*x9/��?A             \@�t�b��     h�h4h7K ��h9��R�(KKKK��h��B�       �h@      A@      D@      .@     �W@     h�@      ?@     8�@      0@      $@     �T@     �P@     p�@     ��@      3@     �p@     �V@      2@      8@      $@      H@     @n@      *@     h�@      @      @     �A@      A@     �w@      j@      @     �`@     �T@      (@      6@      $@     �C@     �k@      (@     |@      @       @      @@      =@     `u@      i@      @     �^@      6@      @      &@      @      (@      S@      �?      i@                      ,@      @      \@     �U@       @      M@      0@      @      @      @      "@     �F@             �Y@                      &@      @      M@     �I@       @     �D@      @              @              @      ?@      �?     �X@                      @       @      K@      B@              1@     �N@      "@      &@      @      ;@     `b@      &@      o@      @       @      2@      6@     �l@     �\@      @     @P@      ;@      @      @       @      (@      G@      @     �P@       @              @       @     �V@     �A@      @      ;@      A@      @      @       @      .@     @Y@       @     �f@      �?       @      *@      ,@     �a@     �S@              C@       @      @       @              "@      3@      �?      S@      @       @      @      @      A@       @              "@       @      @       @              @      2@      �?      N@      �?              @      @      ?@       @              "@      �?      @                              @              @                      �?      �?      @                              @      @       @              @      &@      �?     �L@      �?               @      @      :@       @              "@                                      @      �?              0@       @       @                      @                                                                      �?              &@       @                              @                                                              @                      @               @                                                     �Z@      0@      0@      @     �G@     �u@      2@     �@      $@      @      H@      @@     `w@     0t@      (@     @a@     �W@      0@      0@      @     �G@      t@      2@     0�@       @      @      E@      @@      u@     Ps@      (@     �`@      G@      $@      "@      �?      5@     `b@       @     �h@      @       @      4@      .@     @a@      ]@      @      R@      @      @              �?      @      0@       @      ;@       @              @              @@      @               @     �C@      @      "@              2@     ``@      @     @e@      @       @      ,@      .@     �Z@     @[@      @      P@     �H@      @      @      @      :@     �e@      $@     v@      �?      @      6@      1@      i@      h@       @      O@     �B@      @      @       @      4@      [@       @     `k@      �?      @      6@      &@     �`@      c@      @     �H@      (@      @      @       @      @     @P@       @     �`@                              @     @P@      D@       @      *@      &@                                      ;@             �V@       @              @              B@      ,@              @      @                                      @              *@                       @              @      @              �?      @                                      @               @                       @              �?                      �?                                              @              @                                       @      @                      @                                      4@             �S@       @              @             �@@       @              @      @                                       @              4@                                       @      @               @                                              2@              M@       @              @              9@      @              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��bkhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @2m��y�?�	           ��@       	                   �=@�GU3_��?�           ̥@                          �1@i��N �?�           ��@                           �?k�Y�H��?B            ~@������������������������       �����=&�?�            �n@������������������������       �t��A��?�            @m@                           !@��Q#y��?f           ��@������������������������       ��u��<��?\           ޠ@������������������������       �     ��?
             0@
                           �?΁�>�?V            �`@                          �?@ffffff�?             D@������������������������       ��W��H��?             1@������������������������       ���"8̺�?             7@                           @��nV�?:            �W@������������������������       ��z�G��?3             T@������������������������       �l�l��?             .@                           �?)P�e]��?�           ��@                          �:@辕lC�?A           �@                           @�BDY\�?           �z@������������������������       ��l�]��?�             q@������������������������       ���/����?a            �c@                           @f�Ya��?3            @T@������������������������       �      �?(             P@������������������������       ��"�O�|�?             1@                           @*�N�k��?�           (�@                           �?Y롯�[�?            �{@������������������������       ��J]`	�?(            �L@������������������������       �������?�            0x@                           @�o`�v�?l             e@������������������������       �&�MN��?_            @b@������������������������       �d!Y�B�?             7@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      8@     �B@      7@     �X@      �@     �A@     ��@      .@      @     �S@     �R@     �@     ��@      3@     Pp@     `c@      ,@      ;@      2@      S@     �}@      <@     (�@      (@      @     �Q@      O@     P@     �y@      1@     �j@     �b@      ,@      ;@      2@     �Q@     P|@      :@     X�@       @      @      Q@     �N@     @~@     �x@      1@      j@     �B@      �?       @       @      ,@     @S@      "@     �V@      �?      �?      &@      ,@     �S@     @V@      @     �E@      0@      �?      @       @      ,@      C@       @      >@      �?      �?      @      $@      E@     �E@      @      9@      5@               @                     �C@      �?      N@                      @      @      B@      G@      �?      2@     @\@      *@      3@      0@     �L@     �w@      1@     ��@      @       @     �L@     �G@     `y@      s@      (@     �d@     @\@      *@      3@      0@      L@      w@      ,@     x�@      @       @     �L@     �G@     `y@      s@      (@     �d@                                      �?      @      @       @                                               @               @      @                              @      6@       @      M@      @               @      �?      1@      *@              @       @                              @      @              9@                                              @              �?      �?                              @                      "@                                              �?              �?      �?                                      @              0@                                              @                      @                                      3@       @     �@@      @               @      �?      1@      "@              @      @                                      *@       @      ?@      �?               @      �?      *@      "@              @                                              @               @      @                              @                             �E@      $@      $@      @      7@     �d@      @     �y@      @      @       @      *@     �m@     �`@       @      G@      :@      @       @       @      ,@      T@      @     �b@       @       @      @      @     �[@      P@       @      ;@      6@      @      @       @      &@      Q@      @     �\@               @      @      @     �X@      N@              9@      5@      @      @              "@     �E@      @     �O@               @      �?      @      K@     �D@              4@      �?      �?               @       @      9@              J@                      @              F@      3@              @      @      �?       @              @      (@              A@       @                      @      (@      @       @       @       @      �?       @              @      (@              8@       @                      @      &@       @       @               @                                                      $@                                      �?       @               @      1@      @       @      @      "@     @U@      @     �p@      �?      �?      �?      @     �_@     �Q@              3@      &@      �?       @      @       @      G@      @     �h@      �?      �?      �?      @     �V@      L@              0@       @               @              @       @      �?      1@                                      2@      @              @      "@      �?              @      @      F@       @     �f@      �?      �?      �?      @     @R@      I@              $@      @      @                      �?     �C@              Q@                                     �A@      ,@              @      @      �?                      �?      <@             @P@                                      >@      *@               @               @                              &@              @                                      @      �?              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJaڋAhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             @D|a���?�	           ��@       	                    �?ͽ��a��?�           ʫ@                           �?�k�bZ�?�           8�@                           �?�Z?�"�?o           ��@������������������������       ���ɑ:�?�            �p@������������������������       �C� 3��?�            �v@                            @�X0ki�?�           X�@������������������������       ��d���?           8�@������������������������       ����+��?�            �i@
                            @~1����?�           \�@                            �?T=�N]_�?e           D�@������������������������       ��D��/��?�           �@������������������������       ���f���?�            �t@                           �?:���d��?L           0�@������������������������       �lm����?�            0u@������������������������       ��Rޞ4��?t            `f@                           �?�V��+�?�            @v@                            �?o�ŏ1�?"             I@                           8@�1,D^��?            �@@������������������������       ��&5D�?             1@������������������������       �     @�?             0@������������������������       �|�l�]�?             1@                          �;@0�Ȕ-�?�             s@                            �?ڐf/;�?�            p@������������������������       �/����?'             L@������������������������       �};�r�?v             i@                            �?�-�?��?            �H@������������������������       ��>�>��?             .@������������������������       �l��\��?             A@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `f@      >@      H@      6@     �]@     ؃@      D@     ��@      8@      @     �R@     �Q@     Ȇ@     ��@      4@      p@     `e@      =@      G@      4@     �[@     ��@     �@@     8�@      6@      @      P@     �P@     Є@      ~@      4@      m@     @V@      0@      C@      *@      R@     pr@      6@     �x@      1@      �?      @@     �E@     �q@     �l@      *@     �]@     �@@      @      7@      @      4@      ]@       @     �d@      @              &@      .@      V@     @U@      @      K@      @              @       @      @      F@             �T@      �?               @      "@     �H@      >@      @      6@      ;@      @      1@      @      0@      R@       @     @T@      @              @      @     �C@     �K@       @      @@      L@      &@      .@      @      J@     `f@      4@     �l@      (@      �?      5@      <@     �h@      b@       @      P@     �J@       @      ,@      @     �G@     �a@      1@      e@      (@      �?      (@      ;@     �c@      \@       @      K@      @      @      �?              @      C@      @      N@                      "@      �?     �D@     �@@              $@     �T@      *@       @      @      C@     �r@      &@     ��@      @       @      @@      7@     �w@     @o@      @     �\@      Q@      (@      @      @      >@     �k@      $@     @x@      @      �?      ?@      1@     �p@     �h@      @     @X@      D@      &@       @      @      1@     �f@      @     0t@       @              ,@       @     �j@     �a@       @      N@      <@      �?      @              *@      D@      @     @P@      @      �?      1@      "@     �J@     �J@      @     �B@      ,@      �?       @       @       @      T@      �?     @k@              �?      �?      @      \@      K@              2@       @               @       @      @      M@      �?      b@              �?      �?      @     �L@     �B@              1@      @      �?                      @      6@             @R@                              �?     �K@      1@              �?       @      �?       @       @      "@      D@      @     �`@       @              $@      @     �O@      H@              9@      �?              �?               @       @              1@                      �?              2@       @                      �?                              �?      @              "@                      �?              ,@      �?                      �?                                       @              @                      �?              $@                                                              �?      @              @                                      @      �?                                      �?              �?       @               @                                      @      �?                      @      �?      �?       @      @      @@      @     �]@       @              "@      @     �F@      G@              9@      @      �?      �?       @      @      @@      @     �S@       @              @       @      E@      G@              8@       @      �?      �?       @      @       @      @      $@       @              �?              $@       @              @      @                              @      8@      @     @Q@                      @       @      @@      C@              4@                                                             �C@                      @       @      @                      �?                                                               @                      @       @                              �?                                                              ?@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ	6CThG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@"�e{��?�	           ��@       	                    �?q�Sn��?y           "�@                            @]����?�           ��@                          �1@��x5ZX�?�           ��@������������������������       �?����?�            pp@������������������������       ���H#�?           �@                          �:@ajgH��?           �{@������������������������       �3����?           pz@������������������������       �躍`3�?             1@
                          �9@�M]f#=�?�           ��@                            @���0�?0           ��@������������������������       �|��%��?	           ��@������������������������       �Ggl����?'           `|@                           @�-�� �?q            �h@������������������������       �؋1�K�?X            `c@������������������������       ���ƄIU�?            �E@                           @8�Ț� �?           �{@                           @H��B�?�            �t@                          @@@jȪ^*%�?�            �p@������������������������       �W���'�?�            �l@������������������������       ����(\��?             D@                            �?_k,D	��?#            �M@������������������������       �ףp=
�?             $@������������������������       �{�+h��?            �H@                           @�Ϭ&�S�?I            �[@                            �?�������?-            @P@������������������������       �     ��?             0@������������������������       �ھBNb&�?%            �H@                           @0�;A�L�?            �F@������������������������       �JȬ�@��?            �@@������������������������       �      �?             (@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �f@      A@     �B@      =@     �Y@     ��@      @@     ��@      .@      $@      R@      P@     `�@     ��@      6@     �o@     �c@      >@     �A@      =@     �W@     p�@      =@     ��@      (@       @     �P@     �M@     ��@     @      5@     �l@     �T@      7@      9@      (@      J@      r@      .@     `w@      @      @      A@      >@     �r@     �j@      @     @Z@     �P@       @      5@      (@     �E@      j@      "@     �n@      @       @      =@      >@      i@      d@      @     @U@      4@      �?      $@              0@     �C@      @     �A@      �?      �?      "@      $@      I@     �F@       @      4@      G@      @      &@      (@      ;@      e@      @     `j@       @      �?      4@      4@     �b@     �\@      @     @P@      0@      .@      @              "@     �T@      @      `@              @      @             �X@     �J@              4@      0@      $@      @              "@      T@      @     �_@              @      @             �W@     �I@              4@              @      �?                       @               @                                      @       @                      S@      @      $@      1@      E@     �r@      ,@     0�@      "@      @      @@      =@     px@     �q@      ,@     @_@     �Q@      @      $@      &@     �@@     �q@      *@     p@      "@      @      <@      <@     0u@     �n@      ,@     �[@      J@      @      @      @      =@      j@      *@     Pt@      @      @      8@      4@     �n@     �i@      &@     @W@      3@       @      @      @      @     �R@             @f@      @              @       @     �W@      C@      @      2@      @      �?              @      "@      2@      �?     �G@                      @      �?      J@      D@              ,@      @                      @      "@      *@      �?     �B@                      @      �?      B@     �A@               @              �?                              @              $@                                      0@      @              @      6@      @       @              "@     �Q@      @      d@      @       @      @      @     @V@      C@      �?      8@      4@      @       @               @      L@      @      Z@      @       @      @      @     �P@      >@      �?      7@      3@      @       @              @      F@      @     @U@      @       @       @      @      J@      =@      �?      1@      0@      @       @              @     �C@       @      Q@       @               @      @      H@      =@              (@      @                              �?      @      �?      1@      �?       @                      @              �?      @      �?                              @      (@              3@                       @              .@      �?              @                                                                                                      "@      �?                      �?                              @      (@              3@                       @              @                      @       @                              �?      .@             �L@                       @       @      6@       @              �?       @                              �?      $@              =@                      �?              .@      @              �?                                      �?                      (@                                       @      �?                       @                                      $@              1@                      �?              *@      @              �?                                              @              <@                      �?       @      @       @                                                              @              3@                      �?       @      @       @                                                                              "@                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJY��hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @n�Wej��?�	           ��@                            �?�(]��?�           �@                           !@F��?4           R�@                           �?�	"����?,           6�@������������������������       ��'�ʹD�?6           ��@������������������������       �앇�|��?�           ��@������������������������       ���>4և�?             ,@                           @Pôn���?�           H�@	       
                    �?     �?C            �@������������������������       ���#���?6            @V@������������������������       ��_ͷ���?           pz@                           �?��PkX�?u             i@������������������������       ��GN��?1             V@������������������������       ���H��?D            @\@                           �?޽5A���?�           \�@                           @Ͻ���^�?8           �~@                           @i�����?�            `t@������������������������       �Ԍ/(��?�            Pq@������������������������       ����>�{�?            �H@                           @76ܺe$�?n            �d@������������������������       ���æ�,�?G            �Y@������������������������       �f���n[�?'            �N@                          �3@F��,a�?�           h�@                           @�B�	J�?�            �i@������������������������       � ��5���?d            @c@������������������������       �vL�/�V�?            �J@                           @XC�n��?�            �y@������������������������       ���=ܰ1�?�            �q@������������������������       �Y��&\x�?Q            �`@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@      A@      J@      <@     �Z@     ��@      @@      �@      (@      @      N@     @R@     ؆@     P�@      5@     �p@     `d@      ;@     �B@      :@     �U@     ~@      <@     H�@      "@      @      J@      O@     �@     Px@      3@     �k@     @_@      1@      7@      2@      H@     �w@      7@     x�@      @             �@@      E@     �x@     �p@      $@      b@     �^@      1@      7@      2@      H@     0w@      3@     p�@      @             �@@      E@     �x@     �p@      $@      b@     �M@      @      .@      "@      8@     �f@      "@     `g@      @              2@      7@      b@     �^@      @      T@      P@      (@       @      "@      8@     �g@      $@     0w@      �?              .@      3@     @o@     `b@      @      P@       @                                      @      @      �?                                              �?                      C@      $@      ,@       @      C@      Z@      @     �^@      @      @      3@      4@     @^@     �]@      "@     @S@      A@      @       @       @     �@@     �P@      @     �V@       @      @      ,@      1@     @W@      Q@      @     �L@       @      �?      @      �?      @      *@       @      $@      �?              @      @      3@      @      @      3@      @@      @      @      @      ;@      K@       @     @T@      �?      @      &@      ,@     �R@     @P@       @      C@      @      @      @              @     �B@      �?      ?@       @      �?      @      @      <@      I@      @      4@      �?      @      �?              @      2@      �?      2@       @                              0@      2@       @      @      @              @               @      3@              *@              �?      @      @      (@      @@       @      0@     �H@      @      .@       @      5@     `f@      @     �y@      @      �?       @      &@      k@     �`@       @     �F@      B@      @      *@              &@     @R@      @      b@       @      �?      @      @     �W@      Q@              ;@      9@       @      (@              @     �J@      �?     �T@      �?              @      @      Q@     �F@              7@      7@       @      (@              @      C@      �?     �R@      �?              @      @     �N@     �@@              4@       @                              @      .@              @                                      @      (@              @      &@      @      �?              @      4@       @     �O@      �?      �?      �?       @      :@      7@              @      &@      �?      �?              @      1@              C@      �?      �?               @       @      2@               @              @                       @      @       @      9@                      �?              2@      @               @      *@      �?       @       @      $@     �Z@      �?     �p@      �?              @      @     �^@     @P@       @      2@      @                      �?      @      <@      �?     @S@                      �?      �?     �J@      :@              @      @                      �?      @      0@      �?     �P@                              �?     �D@      3@               @      @                               @      (@              &@                      �?              (@      @              @      @      �?       @      �?      @     �S@              h@      �?               @      @     @Q@     �C@       @      &@      @      �?       @      �?      @      E@             �b@                       @       @      G@      3@              @      �?                                      B@             �E@      �?                       @      7@      4@       @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ<2�4hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @��ۦ��?�	           ��@       	                   �:@��.XS��?�           �@                            �?�6�O��?�           ��@                           @ �{��?           ��@������������������������       �R���*�?�           �@������������������������       ��\�6��?x            �g@                           �?�����y�?�            �@������������������������       ��$�֔�?�           ��@������������������������       �0vh�)C�?           �@
                          �@@B~��E�?�            �x@                          �?@�P�c��?�            �v@������������������������       ����L�?�            �t@������������������������       ����2�?            �B@                          �A@     p�?             @@������������������������       ��ˠT�?             6@������������������������       ��(\����?             $@                           �?#f&->�?�           ��@                           @γWF2G�?�            �t@                           @I�]����?�            �q@������������������������       ��$uf��?�            �o@������������������������       �������?            �@@                          �6@��{�<�?            �E@������������������������       �7��d��?             A@������������������������       ��q�q�?             "@                           @�-:z�?�           ��@                           �?� ��}�?]           ��@������������������������       ��ih>(y�?           �|@������������������������       �Wt���?C            �Z@                           �?�����?x            �g@������������������������       ��:f���?>            �W@������������������������       �%'��]�?:            �W@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `h@     �A@     �C@      @@      Z@      �@      ;@     ��@      2@       @     @W@     �K@     X�@     �@      1@     �p@     �b@      4@      =@      9@     �U@     �}@      8@     ��@      .@      @     �T@     �H@     ��@     �w@      1@     �j@     �_@      1@      9@      4@      S@     0z@      2@     ��@      (@      @     �R@      G@     �~@      u@      .@     @g@     �C@      @      "@       @      1@     `b@      @     �n@       @              1@      @     @f@     �]@      @      =@     �@@      @      "@      @      "@     �\@      @      e@      �?              *@      @     @b@     �Y@       @      5@      @      �?              @       @      @@              S@      �?              @              @@      .@       @       @      V@      $@      0@      (@     �M@      q@      *@     �s@      $@      @      M@     �C@     `s@     �k@      &@     �c@      B@      @      &@      $@      B@     �b@       @      a@       @      @      (@      5@     �a@     @X@      @     �S@      J@      @      @       @      7@     @^@      @     �f@       @              G@      2@      e@     �^@      @     �S@      8@      @      @      @      $@     �J@      @     @`@      @      �?       @      @     �S@      C@       @      <@      5@      @      @      @      $@     �G@      @     @_@      @      �?       @      @     @R@      <@       @      :@      3@      @      @      @      $@     �F@      @      Z@       @      �?       @      @     �P@      :@      �?      :@       @                                       @      �?      5@      �?                              @       @      �?              @                                      @              @                                      @      $@               @      @                                      @              @                                      @       @                                                              @               @                                      �?       @               @      F@      .@      $@      @      2@      e@      @     0w@      @      �?      $@      @     �n@     �`@              J@      $@      @       @       @      @     �G@      �?     �Y@                      @       @     �V@      ?@              >@       @      @       @       @      @     �D@      �?     @V@                       @      �?     @U@      7@              9@       @               @       @      @      D@      �?     �T@                       @      �?     �P@      5@              7@              @                              �?              @                                      2@       @               @       @                                      @              *@                      @      �?      @       @              @       @                                      @              @                      @      �?       @       @              @                                                              @                                      @                              A@      (@       @      @      ,@     @^@       @     �p@      @      �?      @      @     @c@     �Y@              6@      ?@       @      @       @      *@     �V@       @     @g@      �?      �?      @      @      _@     �R@              2@      =@      @      @       @      $@     �Q@      �?     �c@      �?      �?      @       @     �V@     �P@              0@       @      @      �?              @      4@      �?      >@                               @     �@@       @               @      @      @      �?      @      �?      ?@             �T@       @                              >@      <@              @              �?      �?      @      �?      1@             �D@                                      ,@      ,@              @      @      @                              ,@              E@       @                              0@      ,@              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�$hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             �?�:���?�	           ��@       	                     @$*�6H�?G            �@                          �=@ _�����?           ��@                            �?`��v���?�           ̒@������������������������       �����?           `y@������������������������       �M�s���?�           �@                           @Z�x-��?            �I@������������������������       �=[y���?             A@������������������������       �� =[y�?
             1@
                          �0@,8��[`�?0           �}@������������������������       �����H�?             2@                          �=@y��+5�?%           �|@������������������������       �J��.�&�?           0{@������������������������       ����N8�?             5@                          �;@j(uΪ��?Y           �@                            @�xi���?�           8�@                           �?o���?r           �@������������������������       ���8��t�?v             h@������������������������       �z��&���?�           �@                           @�"�B���?K           ��@������������������������       ���s����?E           P�@������������������������       �{�G�z�?             $@                          �<@�7!�H��?�            `o@                           @@�P�a��?%             N@������������������������       �x?r����?             F@������������������������       �      �?             0@                          �>@���\��?w            �g@������������������������       ��1�c��?5            @V@������������������������       �֙]!��?B            �Y@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `i@      C@     �E@      7@      W@     ��@     �A@      �@      1@       @     �U@     �L@     x�@     ��@      .@     �r@     @W@      ;@      =@      "@      K@     �s@      3@     px@      "@      @      A@      @@     `r@     @n@      "@     �d@     @R@      1@      7@      "@      G@      l@      0@     Pp@       @      @      :@      <@      i@     �f@      @     ``@     �P@      1@      7@      "@     �F@     �k@      0@     �m@       @      @      :@      <@     �h@     `e@      @      `@      *@      �?      @       @      (@      T@      @     �Z@                      "@      *@     �Q@      M@       @      >@     �J@      0@      3@      @     �@@     �a@      $@     ``@       @      @      1@      .@     �_@     @\@      @     �X@      @                              �?      @              8@                                      @      "@              @      @                              �?      @              4@                                       @       @              �?       @                                                      @                                       @      @               @      4@      $@      @               @     �V@      @     @`@      �?      �?       @      @     @W@      O@       @      B@                                      �?      �?       @                                              @      @              @      4@      $@      @              @     @V@      �?     @`@      �?      �?       @      @     �V@     �K@       @      @@      0@      $@      @              @     �U@      �?     �_@      �?      �?       @      @     @T@     �K@              @@      @                                       @              @                                      "@               @             �[@      &@      ,@      ,@      C@     pu@      0@     ȅ@       @      @     �J@      9@     �z@     @r@      @     @`@     @Z@      "@      ,@      ,@      B@     �r@      *@     X�@      @      �?      I@      8@     �w@     `q@      @      ]@     �V@      @      *@      @      =@     �k@      "@     w@      @      �?      H@      3@     pp@     `k@      @     �X@      ,@               @       @      @      ,@       @     �L@                       @       @      B@      8@              <@     @S@      @      &@      @      :@      j@      @     �s@      @      �?      D@      1@     `l@     `h@      @     �Q@      ,@      @      �?      @      @     �R@      @     @k@                       @      @      ^@     �M@              1@      ,@      @      �?      @      @      R@      @      k@                       @      @     �]@      K@              1@                                              @              �?                                      �?      @                      @       @                       @     �F@      @     �[@      @       @      @      �?      E@      ,@      @      ,@              �?                              ,@              :@                                      "@       @       @                      �?                              (@              0@                                      @       @       @                                                       @              $@                                      @                              @      �?                       @      ?@      @      U@      @       @      @      �?     �@@      @      �?      ,@      @      �?                              .@              F@      @              �?              0@       @              @       @                               @      0@      @      D@      �?       @       @      �?      1@      @      �?      &@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @!�نՖ�?�	           ��@       	                   �<@`���?�           2�@                           �?���-�?q           ��@                            �?G�!����?�            `u@������������������������       �����g�?^             b@������������������������       ���D)4�?�            �h@                          �1@��]�0�?�           �@������������������������       �n��y*d�?           �|@������������������������       ���2m7�?�           ��@
                           �?�x���t�?|            @j@                            �?u��A���?%             N@������������������������       ��q�q�?             8@������������������������       ��������?             B@                           @�R(Z��?W            �b@������������������������       ���8u���?<            �Y@������������������������       ���8��x�?             H@                          �;@"w_F>��?�           ��@                          �5@�R�"�?d           ��@                           @�qg	�9�?u           ��@������������������������       ��B�iߗ�?9           �|@������������������������       ��'�i�n�?<            @X@                           �?�qǵ�?�             x@������������������������       ���(\��?e             d@������������������������       ������?�             l@                          �=@     ��?O             `@                           �?~�:pΈ�?             I@������������������������       �q�{���?             5@������������������������       ����ϭ�?             =@                           �?�Y� ���?0            �S@������������������������       �΃�\W�?             =@������������������������       ���_�q�?            �H@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @i@      7@      J@      >@     @`@     ��@      C@     0�@      ,@      @     �U@     �K@     ؇@     p@      0@     �p@     @c@      0@      E@      8@      Z@     P|@      B@     8�@      (@      @     �R@     �G@     `�@     �x@      ,@     �l@     �b@      .@      C@      8@     �Y@     �z@     �@@     p�@      "@      @     �P@     �F@     �~@      x@      (@     �j@      1@      @       @      @      &@     �@@             �T@       @              ,@      @     �T@      G@              D@      @      �?               @       @      0@              F@                      "@      �?     �D@      .@              @      &@       @       @       @      "@      1@             �C@       @              @      @      E@      ?@             �@@     ``@      (@      B@      4@      W@     �x@     �@@     ؀@      @      @      J@     �D@     �y@      u@      (@     �e@      >@       @      @      �?      7@     �W@      ,@     @U@                      "@      &@     �Q@     �S@      �?      @@     @Y@      $@      >@      3@     @Q@     �r@      3@     `|@      @      @     �E@      >@     u@     @p@      &@     �a@      @      �?      @              �?      <@      @     @V@      @               @       @     �@@      *@       @      1@      @      �?      @              �?      @              >@                       @              @      @              �?                                      �?      �?              4@                                      �?                      �?      @      �?      @                      @              $@                       @              @      @                                                              6@      @     �M@      @              @       @      =@       @       @      0@                                              0@      @      ?@      @              @       @      5@      @       @      0@                                              @              <@                      @               @      @                      H@      @      $@      @      :@     `f@       @     Px@       @              (@       @     �m@     �Z@       @      B@     �D@      @      "@      @      7@     �c@       @     Pt@       @              (@      @      k@      Z@              A@      <@       @      @      @      4@      R@      �?     �i@      �?               @      @      ]@      P@              :@      9@       @      @      @      4@      M@      �?     �c@      �?              @      @     @Y@     �M@              4@      @                      @              ,@              H@                      @              .@      @              @      *@      @      @              @      U@      �?     @^@      �?              @      �?      Y@      D@               @      &@      �?      @              �?     �F@      �?     �D@      �?              �?              C@      0@              �?       @      @                       @     �C@              T@                      @      �?      O@      8@              @      @              �?              @      7@              P@                              �?      7@       @       @       @      @              �?                       @              ?@                                      @       @               @      @              �?                      �?              &@                                       @      �?               @                                              @              4@                                      �?      �?                      @                              @      .@             �@@                              �?      4@               @              @                              @      @              $@                              �?      @               @              �?                                      "@              7@                                      0@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�]NKhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�<�Od��?�	           ��@       	                   �1@����+�?P           ��@                          �0@��4���?�            �s@                           �?�t۟=��?I            @[@������������������������       �և���X�?#             L@������������������������       �>α�
��?&            �J@                           �?��*���?�            �i@������������������������       ��A�f���?#             I@������������������������       �j����?b            �c@
                          �3@~O&�/��?�           Ԗ@                           @��#Vn��?�             w@������������������������       �.^���?�?�            pp@������������������������       �6�'�q�?D            @Z@                          �7@>��d&�?�           �@������������������������       �5wrxV�?{           ��@������������������������       ��l n��?-           `~@                            @ �j�.��?5           ��@                            �? J�B�?�           ��@                          �2@&d� ���?�           d�@������������������������       ���C��?�            Pr@������������������������       ��]Q��?           ��@                          �2@Xه7"��?�            �x@������������������������       �Έ����?=             Y@������������������������       �����?�            �r@                           �?�@�6���?�           ��@                           @�1��k�?a             c@������������������������       ���'��?Y            @a@������������������������       �^N��)x�?             ,@                           �?�!م���?&           �}@������������������������       �^���sf�?�            `r@������������������������       �0��k���?j            �f@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@     �C@      C@      >@     @X@     ��@      >@     p�@      *@      @      W@      O@     ��@     @�@      7@      p@     @Z@      3@      9@      .@     �N@     �p@      0@     {@      @      @     �J@      ?@     �t@     �p@      $@      a@      2@      @      "@              5@     �E@      @      K@              �?      $@      (@      H@      M@       @      =@       @      �?      �?              (@      ,@      @      1@                      @      @      4@      5@      �?       @              �?                      $@       @      �?      "@                      @      �?      &@      .@               @       @              �?               @      (@       @       @                       @       @      "@      @      �?      @      0@      @       @              "@      =@      @     �B@              �?      @      "@      <@     �B@      �?      5@      @              @              �?      @      �?      .@                       @      �?      @      @               @      (@      @       @               @      8@       @      6@              �?       @       @      9@     �@@      �?      *@     �U@      .@      0@      .@      D@     �k@      $@     �w@      @      @     �E@      3@     �q@      j@       @     �Z@      ,@      @      @      �?      "@      E@      �?     �^@              �?      "@      @     �S@     �G@      @      8@      @      @      @      �?      "@      @@             �X@              �?      @      @     �H@      >@       @      0@       @                                      $@      �?      7@                      @      @      =@      1@      @       @     @R@      $@      (@      ,@      ?@     �f@      "@     p@      @      @      A@      *@     �i@      d@      @     �T@      ?@      @      "@      @      7@     �Y@      @      ^@      @       @      8@      (@     �^@     @Y@       @     �B@      E@      @      @      "@       @     �S@       @      a@      �?      �?      $@      �?     �T@      N@      �?      G@     @W@      4@      *@      .@      B@     �t@      ,@     X�@      @       @     �C@      ?@     �z@     �q@      *@      ^@     @R@      1@      $@      &@      >@     �l@      (@     �z@      @       @     �A@      8@     �r@     `l@      *@      X@      E@      0@      @       @      ,@     @f@       @     �u@      @              .@      (@     �l@     �c@      @     �O@      2@      �?                      @     �H@      �?     �[@                      @      @      J@      C@       @      $@      8@      .@      @       @      &@      `@      @      n@      @              (@      @     `f@      ^@      @     �J@      ?@      �?      @      @      0@     �J@      @     �R@               @      4@      (@     �P@     @Q@      @     �@@      "@               @      �?      �?      5@       @      &@                      @      @      @      :@      @      *@      6@      �?       @       @      .@      @@       @     �O@               @      0@      "@     �O@     �E@      @      4@      4@      @      @      @      @      Z@       @     0p@      �?              @      @     �`@     �M@              8@      @                      �?      �?      "@             @P@                      @      �?     �B@      2@              *@      @                      �?      �?      @             �O@                      @              @@      1@              &@      �?                                       @               @                              �?      @      �?               @      0@      @      @      @      @     �W@       @     @h@      �?              �?      @     �W@     �D@              &@      "@      @      �?      @      @      L@       @     @]@      �?                      @     �H@      @@              &@      @               @              �?     �C@             @S@                      �?              G@      "@                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�=�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @�6*���?�	           ��@       	                   @@@c�:����?q           d�@                           �?6��>$~�?c           �@                            @�O�3�?�           ��@������������������������       �pQ��0��?           �z@������������������������       ��O�偯�?�            Pr@                          �4@o�y3ҍ�?�           ��@������������������������       ����n��?n           ��@������������������������       ��3��?-           @@
                           �?@�"s�?             =@������������������������       �P�|�@�?             1@������������������������       ��q�q�?             (@                           �?h����?>           `�@                           @�ee~��?B           ��@                           @�@��\,�?            |@������������������������       �x���`F�?f            �c@������������������������       �x7���q�?�            0r@                            @QM�ıx�?$            }@������������������������       �)S�����?�            `x@������������������������       �AD˩�m�?4            �R@                          �<@�H+���?�           x�@                          �0@p�00sV�?�           ��@������������������������       ���_�}�?(             Q@������������������������       ���Qa7�?�           ��@                            �?��p6��?Q            �_@������������������������       ��-Xm�?            �D@������������������������       ��
)8G�?7            @U@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @g@      9@      D@      <@      X@     ��@      E@     �@      2@      @     �Q@      R@     ��@     ��@      0@     `q@     �X@      *@      =@      1@     �H@     0s@      $@     @       @      @      <@      >@     �x@     �g@      @     `a@     @X@      *@      =@      1@     �E@     0s@      $@     0~@      @      @      <@      >@     �x@     �g@      @      a@      =@       @      .@      @      1@     @[@       @     @l@      �?              1@      "@      a@     @U@             �N@      3@       @       @       @      0@      N@      �?     �[@      �?              ,@      "@      W@     �G@              D@      $@              @      @      �?     �H@      �?     �\@                      @              F@      C@              5@      Q@      @      ,@      &@      :@     �h@       @     p@      @      @      &@      5@      p@     @Z@      @     �R@     �E@      @      @      @      (@     �_@      @     �\@      �?      @      @      1@     �`@     �G@      @      C@      9@               @      @      ,@     �Q@       @     �a@      @      �?      @      @     �^@      M@             �B@      �?                              @                      ,@       @       @                                      �?      @                                      @                      @               @                                      �?      @      �?                               @                      @       @                                                              V@      (@      &@      &@     �G@     �u@      @@     @�@      $@      �?     �E@      E@     @w@     `u@      (@     `a@      G@      $@      @       @      9@      d@      *@     @l@      @      �?      .@      8@     `c@     �b@      @      R@      A@       @      @      �?       @     �V@       @     �X@       @      �?      @      @      M@      S@      �?     �F@      *@      �?                      @      =@             �G@                      @       @      0@      =@      �?      *@      5@      @      @      �?      @     �N@       @      J@       @      �?      @      @      E@     �G@              @@      (@       @       @      �?      1@     �Q@      @     �_@      @               @      1@     @X@      R@      @      ;@      (@       @       @      �?      ,@     @P@      @     �W@      @              @      1@     �R@     �P@      @      6@                                      @      @              @@                      �?              7@      @              @      E@       @      @      "@      6@     �g@      3@     `v@      @              <@      2@      k@     @h@      @     �P@     �D@       @      @      "@      6@      d@      1@      s@      @              <@      2@      g@     �g@      @      P@      @                       @              @              $@                              �?      1@      ,@              &@      A@       @      @      @      6@     `c@      1@     �r@      @              <@      1@      e@     �e@      @     �J@      �?                                      =@       @      J@       @                              @@      @              @                                              @              0@       @                              (@      @                      �?                                      6@       @      B@                                      4@      �?              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��'hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @B ۋ�{�?�	           ��@       	                   �1@�������?�           �@                           @_"�z�?'           �|@                           @:x�����?�            �u@������������������������       �pi.Y�M�?�            0s@������������������������       ���ճC��?             F@                           @��0�m��?C            @Z@������������������������       �     ��?'             P@������������������������       �������?            �D@
                            �?�Fa���?�           ��@                           !@ѣ��Q/�?^           \�@������������������������       ��ع�L+�?V           �@������������������������       �     @�?             0@                          �7@DV�����?]           H�@������������������������       �6�g4���?�            �v@������������������������       ��h��)��?v            �g@                          �2@�=����?�           �@                           �?�
���?�            �p@                           �?_�g�J�?U            �`@������������������������       �"lxz�,�?              I@������������������������       �������?5            �T@                           @"�A�L�?Z             a@������������������������       �$I�$I��?,            �Q@������������������������       ��0��?.            �P@                          �;@�����_�?�           ��@                           �?ט���?�           �@������������������������       �K	�{�?�            Pr@������������������������       ����_��?�            �w@                           @)O���?V             b@������������������������       ���7f���?O            @`@������������������������       �s
^N���?             ,@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        j@      E@      F@      7@     �[@     X�@      @@     ��@      .@      @     @V@     �L@     �@     0}@      .@     Pp@     �c@      >@      >@      5@      U@     `~@      :@     ��@       @      @      T@      I@     @@     @v@      ,@     �k@      B@      @      @      �?      0@     �W@      &@     �T@       @      �?      *@       @     �Q@     �Q@      �?      E@      ?@       @       @      �?      .@     @S@      @      L@                      *@      @     �J@      H@              D@      7@       @       @              .@      R@      @     �I@                      "@      @      I@     �E@              <@       @                      �?              @              @                      @      �?      @      @              (@      @      �?       @              �?      1@      @      ;@       @      �?              �?      2@      6@      �?       @      @      �?      �?                      .@      @       @       @                      �?      ,@      (@      �?              �?              �?              �?       @              3@              �?                      @      $@               @     �^@      ;@      :@      4@      Q@     �x@      .@     ��@      @      @     �P@      E@     �z@     �q@      *@     `f@      W@      5@      *@      2@     �G@     @t@      &@     8�@      �?              E@      3@      v@      h@       @      _@      W@      5@      *@      2@      G@     �s@      "@     (�@      �?              E@      3@     �u@     �g@       @      _@                                      �?       @       @       @                                      �?       @                      >@      @      *@       @      5@      Q@      @      ^@      @      @      9@      7@     @S@     �W@      @     �K@      0@       @      *@       @      .@      G@      �?      Q@      @      @      4@      5@      D@      R@             �D@      ,@      @                      @      6@      @      J@               @      @       @     �B@      6@      @      ,@      I@      (@      ,@       @      :@     �d@      @     `w@      @              "@      @     �p@     �[@      �?      D@      @              �?      �?      @      <@       @     @W@                      @      @     �V@      :@              "@       @              �?      �?      @      *@              K@                       @      �?      =@      3@              @      �?                                       @              <@                                      ,@      @              �?      �?              �?      �?      @      &@              :@                       @      �?      .@      .@              @      @                                      .@       @     �C@                      �?       @      O@      @              @      @                                      @              .@                                      C@      @               @      �?                                      "@       @      8@                      �?       @      8@       @               @     �E@      (@      *@      �?      4@      a@      @     �q@      @              @      @     �e@     @U@      �?      ?@     �A@      (@      $@      �?      ,@     �[@      @     �k@      @              @      @     �a@     �T@      �?      9@      6@      @      @              (@      K@      @     @T@       @              @       @      M@      A@              @      *@      @      @      �?       @     �L@      �?     �a@       @              �?       @     @U@      H@      �?      3@       @              @              @      :@              M@      @                              ?@      @              @       @                               @      8@              L@      �?                              ?@      @              @                      @              @       @               @       @                                                      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�0hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @�ϳ�xv�?�	           ��@                            �?@n�����?�           ޥ@                           @1�]���?�           D�@                           @i�[�N��?�           ��@������������������������       �3�*���?6           �}@������������������������       ��n#،��?J            �@������������������������       �ŕ�(�?             5@                           �?cc��J�?a           x�@	       
                   �;@�+�9<�?�             m@������������������������       ���y�
�?x            �g@������������������������       ��.�袋�?             F@                           @u��D:�?�           ԗ@������������������������       �v�(Z�?|           ̕@������������������������       ������?S            @`@                          �2@$�a��7�?�           h�@                           @Y��]�?�            `p@                           @��9�-��?x             g@������������������������       �ؒꮃ�?X            @a@������������������������       �i�5���?              G@                           �?��:�^��?6            �S@������������������������       �      �?             4@������������������������       ���hha��?+             M@                           �?�=�'��?!           ��@                           @��8�<T�?�            @w@������������������������       �tn�$�a�?�            �q@������������������������       � 9�����?;             V@                           �?n�����?+            ~@������������������������       ��˹�m�?2             S@������������������������       ��|F��?�            @y@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      7@      I@      ?@     �\@     ��@      6@     ��@      2@      @      Q@      R@     `�@     �@      .@     �n@     `d@      2@     �B@      :@     @V@     �~@      5@     0�@      (@      @     �L@     �L@     �~@     �w@      *@     �h@     �I@      @      @      (@      6@     �g@      *@      u@      @              3@      0@     �i@     �[@      @     �I@     �H@      @      @      (@      1@     `f@      *@     �t@      @              3@      0@     @i@     �[@      @     �I@      <@      @       @       @      *@     @X@      @      c@      �?               @      @     �X@     �A@      �?      3@      5@       @      @      @      @     �T@      "@     �f@      @              &@      "@      Z@     �R@      @      @@       @                              @      "@              @                                       @                              \@      *@      ?@      ,@     �P@      s@       @     `y@       @      @      C@     �D@     �q@     �p@      "@     `b@      *@      @       @      @      &@      ;@             �E@       @               @             �K@     �B@       @      ;@      @      �?       @      @      &@      3@             �A@       @              @              G@      >@       @      ;@       @       @                               @               @                       @              "@      @                     �X@      $@      =@      &@      L@     Pq@       @     �v@      @      @      >@     �D@     �l@      m@      @      ^@     @X@      $@      <@      &@      K@     0p@      @     �s@      @      @      ;@      D@      k@     @j@      @     @Z@       @              �?               @      2@      �?      I@                      @      �?      .@      6@              .@     �E@      @      *@      @      9@      f@      �?     �w@      @       @      &@      .@      p@     �_@       @      G@      @      �?      @      @       @     �A@      �?      R@                      @       @     �T@      ;@              ,@      @              �?      @      @      <@             �E@                      @      �?     @Q@      2@              "@      @              �?      �?      �?      7@              A@                      �?              L@      ,@               @      �?                       @       @      @              "@                       @      �?      *@      @              @      �?      �?      @              @      @      �?      =@                       @      �?      *@      "@              @                      @              @                      @                                              @              �?      �?      �?                              @      �?      6@                       @      �?      *@      @              @      B@      @       @       @      1@     �a@             @s@      @       @      @      *@      f@     �X@       @      @@      7@      @      @              *@     �Q@             �Y@      @      �?      @      @     �R@      I@      �?      2@      7@      @      @              @      M@             �P@      @      �?              @     �O@      D@      �?      &@                      �?              @      *@             �A@                      @              &@      $@              @      *@      �?       @       @      @     �Q@             �i@      @      �?       @      $@     �Y@     �H@      �?      ,@      @              �?                      ,@              3@                                      1@      1@              �?      @      �?      �?       @      @      L@             `g@      @      �?       @      $@     @U@      @@      �?      *@�t�bub��     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJDh�NhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?M�i8���?�	           ��@       	                   �?@�$<g3�?b           ě@                            @Z����8�?N           4�@                           !@���}��?           �@������������������������       ����$��?           �@������������������������       �      �?              @                           @�񞝨>�?7           H�@������������������������       ������?�            pu@������������������������       ���j��M�?f            @f@
                            �?~X�<��?             B@������������������������       �hE#߼�?             .@������������������������       �c>���?             5@                            @�<�w��?b           ��@                            �?{���e�?�           ؗ@                          �@@*t:"��?�           4�@������������������������       �����!��?�           �@������������������������       ��������?             (@                          �4@��?�            �v@������������������������       �^��"��?t            `e@������������������������       �1����?�            �g@                          �;@~�����?�           �@                           @��T�l��?L           ��@������������������������       �j*;�v��?E            �@������������������������       �      �?             (@                           @N<4����?6            �T@������������������������       �dR3?т�?            �D@������������������������       �0�@g���?            �D@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       `k@      @@      =@      9@     @[@     ��@     �@@     �@      0@       @     �R@      P@     ��@     8�@      .@     �o@     @]@      0@      5@      (@      S@      t@      3@     `y@      *@      @     �@@      >@     �t@     �l@      @      a@     @\@      0@      5@      (@      S@     �s@      3@     `x@      &@      @     �@@      >@     �t@     �k@      @      a@     @T@      @      0@      (@     �M@     �k@      2@      n@      $@      @      6@      ;@     `l@     �c@      @     @[@      T@      @      0@      (@      M@     �k@      .@      n@      $@      @      6@      ;@     `l@     �c@      @     @[@      �?                              �?       @      @                                                      �?                      @@      "@      @              1@     �W@      �?     �b@      �?      �?      &@      @     �Z@     �N@      �?      <@      *@              @              &@     �Q@      �?     �V@                      &@      �?     �U@      C@              .@      3@      "@                      @      8@             �M@      �?      �?               @      4@      7@      �?      *@      @                                      @              0@       @                               @      "@                                                              �?              &@                                              @                      @                                       @              @       @                               @      @                     �Y@      0@       @      *@     �@@     �u@      ,@     `�@      @       @     �D@      A@     �z@      r@       @      ]@     @V@      *@      @      "@      >@     �o@      (@     �{@      @      �?      C@      :@     0r@     �i@      @     @Y@     @P@      &@      @      @      ,@     �h@      &@     `w@       @              8@      ,@     `l@     �b@       @     �O@     @P@      &@      @      @      ,@     �g@      &@     Pw@       @              8@      ,@     @l@     �b@       @     �O@                                              $@              �?                                      �?                              8@       @       @       @      0@     �K@      �?     �P@      �?      �?      ,@      (@      P@     �L@      @      C@      .@              �?              @      ?@              4@                      $@      @      4@     �@@      �?      <@      "@       @      �?       @      $@      8@      �?     �G@      �?      �?      @      @      F@      8@      @      $@      *@      @      @      @      @     �W@       @     `n@              �?      @       @     �`@     �T@      �?      .@      (@      @      @      @      �?     @Q@       @     @j@                      @       @     �^@      S@      �?      *@      (@      @      @      @      �?      P@       @     @j@                      @       @     @^@     �Q@      �?      *@                                              @                                                       @      @                      �?                               @      :@             �@@              �?                      $@      @               @      �?                               @      @              6@              �?                      @      @               @                                              6@              &@                                      @       @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�!JhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @���b�?�	           ��@       	                    �?=i���?�           ��@                            �?�6�0[�?           ��@                          �?@8���?M           �@������������������������       �+/�ɯ#�??           h�@������������������������       �
ףp=
�?             4@                           �?\����?�            `r@������������������������       ������H�?             ;@������������������������       ��2�O��?�            �p@
                           @5j��	P�?�           \�@                           �?:FR^jv�?�           @�@������������������������       ������?I            �\@������������������������       ���!)1�?c           ��@                            �?��(��?           x�@������������������������       ��r��M�?�           �@������������������������       ��.*��?�            �i@                           @b�\h1��?�           ,�@                           �?;�#���?$           x�@                           @�����3�?           �y@������������������������       �����(�?�            Ps@������������������������       ���y��?A             Y@                          �2@��޳��?!           `}@������������������������       ���F���?T            �a@������������������������       �!���/��?�            �t@                           �?�u_��?�            �k@                           @     ��?             @@������������������������       ��3_<�?             5@������������������������       �}��7�?             &@                          �5@��E�B��?z            �g@������������������������       �-B����?3             U@������������������������       ��WV��?G             Z@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      @@     �@@      5@      \@     ��@      A@     �@      9@      "@     @R@     �M@     p�@     @      2@     @n@     �c@      3@      9@      0@     @W@     �}@      >@     ��@      5@      @     �M@     �G@     `@     �w@      0@      j@      T@      "@      2@       @      J@     �k@      ,@     pr@      ,@      @      <@      4@      i@     �e@      $@     @[@     �Q@      @      .@      @     �C@     �f@       @     �m@      "@      �?      1@      $@      c@     �_@      @     @R@     �Q@      @      .@      @     �C@     �f@       @     `l@      "@      �?      1@      $@     �b@     �^@      @     @R@                                                              &@                                      @      @                      "@      @      @       @      *@      C@      @     �L@      @      @      &@      $@      H@     �F@      @      B@              �?      �?                      �?              @      @                               @       @              "@      "@      @       @       @      *@     �B@      @     �I@              @      &@      $@      G@     �E@      @      ;@      S@      $@      @       @     �D@     0p@      0@     �|@      @       @      ?@      ;@     �r@     @j@      @     �X@     �D@      @      �?      @      5@     �]@      @      g@       @              *@      ,@     @b@     �S@       @      G@      @      �?              �?      @      .@              6@                       @      @      ;@      (@              6@      B@       @      �?       @      0@     �Y@      @     @d@       @              &@      &@     �]@     �P@       @      8@     �A@      @      @      @      4@     �a@      "@     0q@      @       @      2@      *@     `c@     ``@      @     �J@      :@      @      @      @      $@     @[@      @     `m@      @              "@      @     �`@     �U@      �?      @@      "@      �?      �?      �?      $@      @@       @      D@      �?       @      "@      "@      4@     �F@      @      5@      E@      *@       @      @      3@      g@      @     �x@      @       @      ,@      (@      o@     �\@       @      A@      ?@       @      @      @      3@     �_@      @     �s@      @       @      $@      "@     @j@     �W@      �?      =@      4@      @      @      �?      $@     �R@      @     �Z@      �?              $@      @     �W@     �N@      �?      *@      3@      �?      @              @     �O@      @     �R@      �?              @      @     �Q@     �G@      �?      (@      �?      @      �?      �?      @      &@              ?@                      @              8@      ,@              �?      &@      �?      @      @      "@     �J@      �?     �j@      @       @              @     �\@     �@@              0@      @               @      @       @      .@              H@                              �?     �H@      $@              @      @      �?      �?      �?      @      C@      �?     �d@      @       @              @     �P@      7@              "@      &@      @      �?                      M@             @R@                      @      @      C@      5@      �?      @      @                                       @              @                                      @      $@                      @                                      @              @                                      @       @                                                              @              @                                      �?       @                       @      @      �?                      I@             �P@                      @      @      A@      &@      �?      @      @      @                              1@              @@                      @       @      .@      @              @      @      �?      �?                     �@@              A@                              �?      3@       @      �?       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���(hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @[K��^��?�	           ��@       	                     �?��J��?�            �@                            �?KFx���?           T�@                           �?=�c>���?o           �@������������������������       �JDO�F��?d            `c@������������������������       ��h6)�?           0�@                          @A@E:Kd	�?�           $�@������������������������       �PA��?�           �@������������������������       �      �?              @
                           �?�3Ē(��?�           ��@                           @8��=���?�            @u@������������������������       �i�{#.�?�            `s@������������������������       �
ףp=
�?             >@                           @�t2��?�             x@������������������������       �<�͑7��?�            �s@������������������������       ��z���n�?)            @Q@                           �?|Ѳp�!�?�           $�@                           @Ac�oH"�?)           0}@                           @�#S�w�?�            �r@������������������������       ��K �i�?�            �i@������������������������       ���8��x�?6             X@                           @�	dN��?e            �d@������������������������       ���g�K�?S            �`@������������������������       � \��M�?             A@                          �;@���7�?�           ��@                           @K�Pr�v�?d           @�@������������������������       �('&Η�?
           �y@������������������������       �4T2���?Z            @a@                          @@@dJ�dJ��?5            �S@������������������������       ��?�(ݾ�?%             J@������������������������       ��q-�?             :@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @h@      ;@     �E@      =@     @]@     Є@      9@     ��@      6@      "@     �R@     �M@     ��@     `@      8@     �p@     �a@      5@      A@      9@     @X@     0~@      6@     ��@      4@      @     �K@      J@     �@     @w@      6@     �k@     �X@      0@      9@      2@     @Q@     �v@      1@     ��@      ,@      @     �C@      9@      x@     pp@      "@      b@     �D@       @      @      "@      :@     �e@      @     �s@      @              (@      &@     �g@     �_@       @      N@      @      �?              �?      @      0@             �R@                       @              8@      *@              *@     �A@      @      @       @      6@     �c@      @     @n@      @              $@      &@     �d@     �\@       @     �G@      M@       @      3@      "@     �E@      h@      (@     �q@       @      @      ;@      ,@      h@      a@      @     @U@      M@       @      3@      "@     �E@     �g@      (@     �q@       @      @      ;@      ,@     �g@     �`@      @     @U@                                              @                                                      @      �?                      F@      @      "@      @      <@     �]@      @      a@      @      @      0@      ;@     �^@     @[@      *@     @S@      5@      @      @      �?      ,@     �K@       @      L@      @      @      @      0@     �H@      N@       @     �C@      5@      @       @      �?      ,@     �J@       @     �E@      @      @      @      0@      G@      J@       @      C@                       @                       @              *@      �?                              @       @              �?      7@       @      @      @      ,@     �O@      @      T@              �?      *@      &@     @R@     �H@      @      C@      0@       @      @      @      $@     �K@      @     @P@              �?      (@      &@     �H@      G@      @      @@      @              �?              @       @              .@                      �?              8@      @              @     �I@      @      "@      @      4@     �f@      @     Px@       @       @      3@      @     @l@     @`@       @      F@      7@      @      @      �?      &@     �T@       @     �a@      �?      �?      ,@      @     �U@     @P@      �?      :@      0@              @      �?      $@     @P@      �?     �S@                      *@       @      J@     �D@              2@      &@              @      �?      @      @@      �?      L@                      $@              D@     �@@              *@      @                              @     �@@              6@                      @       @      (@       @              @      @      @       @              �?      1@      �?     �O@      �?      �?      �?       @     �A@      8@      �?       @      @      @       @              �?      $@      �?     �K@      �?      �?      �?       @      9@      5@      �?      @      @                                      @               @                                      $@      @               @      <@      @      @      @      "@     @Y@      �?      o@      �?      �?      @      @     `a@     @P@      �?      2@      ;@      @      @      @      @     �S@      �?      j@                      @      @      `@     @P@      �?      1@      8@       @      @      @      @     �J@      �?     �d@                      @       @      Y@      B@              ,@      @      �?                      �?      9@              F@                      �?      �?      =@      =@      �?      @      �?                               @      7@             �C@      �?      �?                      $@                      �?                                              6@              9@      �?                              @                      �?      �?                               @      �?              ,@              �?                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJƮ�hhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @f"��I��?�	           ��@       	                     �?,+A��?�           ֥@                          �=@CI�`&�?�           ��@                           @��r#I�?z           8�@������������������������       �"`1
��?�           `�@������������������������       ��3#����?�            `k@                          �>@|�l�]�?'             Q@������������������������       �     ��?             0@������������������������       �θ	j*�?             J@
                           @zۧ�i�?L            �@                            �?u%Y
��?�           d�@������������������������       �*/#Hc(�?a           ��@������������������������       �Uy�y�?�           0�@                           @���giu�?\            �d@������������������������       �騷}*_�?L            �`@������������������������       �     `�?             @@                          �;@%��+���?�           x�@                           �?���j�
�?`           ��@                          �0@(���;T�?
            {@������������������������       ��
t�F��?
             1@������������������������       ������?            z@                          �9@}����?V           �@������������������������       ���َ��?6           �~@������������������������       �����[�?              K@                           @)�bpN��?W            `a@                          @@@���]%�?J            @^@������������������������       � �K@��?<            �X@������������������������       �x�W��#�?             7@������������������������       �����K�?             2@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      :@     �C@      9@      Z@     h�@      <@     ��@      0@      @      U@     @P@     H�@     ��@      4@     p@     @e@      6@      >@      5@     �T@     �~@      7@     ��@      *@      @      Q@      N@     �|@     �x@      3@     �j@      O@      @      @      "@      5@      k@      $@     �s@      @              6@      (@      f@     �a@      @      N@      O@      @      @      "@      3@     `j@      "@     �q@      @              6@      &@     @d@     �`@      @     �M@     �I@      @      @      @      .@     @d@       @     �i@      @              6@       @     �`@     @Z@             �I@      &@       @               @      @     �H@      �?      T@                              @      <@      <@      @       @                                       @      @      �?      @@                              �?      .@      $@              �?                                              �?              *@                                       @                                                               @      @      �?      3@                              �?      *@      $@              �?      [@      .@      :@      (@      O@     0q@      *@     Py@      $@      @      G@      H@     �q@      o@      0@      c@     @Z@      .@      7@      (@      O@     �o@      (@     �u@      "@      @      E@     �G@     Pp@     �j@      0@      a@      N@      @      1@      @      C@     �d@      "@     �l@      @      �?      1@      4@     �e@     �]@      @     @S@     �F@      $@      @      @      8@      V@      @     �^@      @      @      9@      ;@     �U@     �W@      $@      N@      @              @                      7@      �?      K@      �?              @      �?      9@     �B@              .@      �?              @                      2@             �F@      �?              @      �?      3@      =@              ,@       @                                      @      �?      "@                                      @       @              �?      I@      @      "@      @      5@      d@      @      y@      @              0@      @     @o@      b@      �?     �F@      E@      @      @      @      3@      a@      @     Pu@      �?              0@      @      l@     `a@             �B@      ;@      @      @      �?      *@      T@      @     �\@                      (@             @W@      O@              4@       @                              @      �?              �?                      �?                      @              @      9@      @      @      �?      $@     �S@      @     @\@                      &@             @W@     �L@              0@      .@               @      @      @     �L@      �?     `l@      �?              @      @     ``@     @S@              1@      .@               @      @      @      L@      �?     @j@      �?              @      @     �Y@     @R@              .@                                      �?      �?              1@                                      =@      @               @       @              @               @      8@             �M@       @                      �?      :@      @      �?       @       @                               @      7@             �K@      �?                      �?      3@      @      �?      @      @                              �?      7@             �F@      �?                      �?      (@      @      �?      @       @                              �?                      $@                                      @                      @                      @                      �?              @      �?                              @      �?              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @y1����?�	           ��@       	                   �0@�[�NX�?           6�@                           @�BE���?z            @g@                           @K�$;z�?7            @V@������������������������       �4$����?+            �P@������������������������       �|�!*�?             7@                           @9�5�3�?C            @X@������������������������       ��<ݚ�?             B@������������������������       �l�(�|�?+            �N@
                           �?xQ�����?�           ¤@                          �=@d.��e�?�           ��@������������������������       �~	�9�~�?�           Đ@������������������������       ��֤����?            �H@                            �?�q��N��?�           ��@������������������������       ���x���?�           D�@������������������������       ��j�P��?�            �v@                           @@�L�'��?�           ��@                           �?�L%����?C           �~@                           @d��m�?�            �s@������������������������       �G�9��?�            �k@������������������������       ����[Ж�?D            @X@                           �?�[0$��?r            �e@������������������������       ��� ��?&             I@������������������������       ��yȔA�?L            @_@                           @�=v�A�?q           �@                           �?��'kM�?           �z@������������������������       �Tܿ^�?7            �T@������������������������       ��1��Ao�?�            �u@                           @�a��H��?c            �b@������������������������       �n�_hD��?Z            �`@������������������������       �     @�?	             0@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      :@      B@      ?@     @[@     �@      A@     t�@      0@      $@      O@     �R@     ��@     Ȁ@      >@     Pp@      d@      2@      >@      :@     @V@     �~@      =@     ��@      .@      @     �J@     �P@     ~@     �y@      ;@     �j@       @      �?       @       @       @     �A@      @      6@      �?      �?      @      "@      B@      B@       @      0@      @              �?              @      "@       @      @                      �?      "@      8@      7@       @      @      @              �?                       @       @      @                      �?      @      0@      6@              @                                      @      �?              @                              @       @      �?       @              @      �?      �?       @      @      :@       @      0@      �?      �?       @              (@      *@              $@      �?      �?      �?       @       @      $@              @                      �?              $@      �?              @      @                              @      0@       @      *@      �?      �?      �?               @      (@              @      c@      1@      <@      8@     @T@     p|@      9@     ��@      ,@      @      I@      M@     �{@     pw@      9@     �h@      S@      &@      2@      ,@     �B@      j@      .@     0p@       @      @      0@      ;@     `d@      d@      "@     @X@      R@      &@      2@      ,@     �@@     �i@      .@     �l@       @      @      0@      ;@     @d@      c@      "@      X@      @                              @      @              =@                                      �?      @              �?     @S@      @      $@      $@      F@     �n@      $@     �{@      @       @      A@      ?@     �q@     �j@      0@     �Y@     �L@      @      @      "@      ;@     @i@       @     �v@      @              *@      7@      l@     @c@      "@     �N@      4@      �?      @      �?      1@     �F@       @     @S@      �?       @      5@       @     �L@     �N@      @     �D@     �E@       @      @      @      4@     �b@      @     �x@      �?      @      "@       @     `n@     �_@      @      G@      0@       @      @       @      @      E@       @     @h@               @      @       @     �`@      L@              9@      &@       @                      @      <@       @     �]@                      @       @     @T@      E@              6@       @                              @      5@       @     �V@                      �?      �?      K@      A@              (@      "@       @                              @              =@                      @      �?      ;@       @              $@      @              @       @      @      ,@             �R@               @      �?             �I@      ,@              @      @              @      �?      �?      @              2@                                       @      &@              �?       @              �?      �?       @      &@             �L@               @      �?             �E@      @               @      ;@      @      �?      @      *@     @[@      @     �h@      �?      �?      @      @     �[@     �Q@      @      5@      :@      @      �?      @      @     �V@      @      a@              �?      �?      @      T@     �K@      @      &@      @                                      0@      �?      ;@                      �?              $@      3@              @      6@      @      �?      @      @     �R@       @     �[@              �?              @     �Q@      B@      @      @      �?      �?                      @      2@              O@      �?               @              ?@      .@              $@      �?      �?                      @      1@              M@      �?               @              9@      ,@              @                                              �?              @                                      @      �?              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJM��#hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                            �;@9L��r�?�	           ��@       	                    �?m��O#��?�           �@                           �?���4BE�?�           ��@                          �0@ 	a��<�?�             m@������������������������       ��Q����?
             4@������������������������       �I�����?�            �j@                          �1@�!��<�?f           ��@������������������������       ��Wb���?�            �m@������������������������       ���H`V�?�           <�@
                           @��=
��?�           x�@                          �3@i��ӳ�?�           ��@������������������������       �:Eh�v�?�            Px@������������������������       �+��-k��?�           �@                          �1@��^�f�?�           ��@������������������������       ��z�^�?r            �e@������������������������       ���~,G�?~           X�@                           @���|*f�?           P|@                           @�e��!�?�            �x@                            �?[B�C~��?�            s@������������������������       �>!,u%@�?.            @T@������������������������       �/����?}             l@                          �<@e���?@            �W@������������������������       ��k���?             ;@������������������������       �aQŜk�?-            �P@                           @rJ�:��?#             K@                           �?�~����?            �E@������������������������       �9��8���?             8@������������������������       ����y4F�?             3@������������������������       ��C��2(�?             &@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@      A@     �F@      7@     @U@     ��@      C@      �@      6@      $@      T@     @P@     ��@     `�@      1@     pp@     �g@      ;@      D@      7@     �R@     ��@     �A@     ��@      2@       @     �Q@     �N@     ��@     �~@      ,@     �l@     �T@      1@      =@      $@      H@      q@      3@     �v@      ,@      @      A@     �@@     pq@      l@       @     �`@      "@      @      @      �?       @      >@       @     �O@      "@              @      @      D@      ;@              7@                       @                       @                                      �?      �?      @      $@                      "@      @      @      �?       @      <@       @     �O@      "@              @      @      B@      1@              7@     @R@      ,@      6@      "@      D@     �n@      1@     �r@      @      @      ;@      =@     �m@     �h@       @     �[@      3@      �?      @      �?      @     �E@      @     �A@              �?      @      @      D@      ?@       @     �A@      K@      *@      .@       @     �@@      i@      (@     �p@      @      @      5@      8@     �h@     �d@      @     �R@      [@      $@      &@      *@      :@     0r@      0@     ��@      @       @      B@      <@     �w@     �p@      @      X@     @R@      @       @       @      (@      d@      @     @v@       @      �?      2@      1@     p@     �b@      @      H@      <@              @      �?      @     �D@      @     @`@                      @      @     �Z@      F@      @      (@     �F@      @      @      @      @      ^@      @     @l@       @      �?      (@      ,@     �b@     @Z@              B@     �A@      @      @      @      ,@     @`@      $@      n@       @      �?      2@      &@     @^@      ]@      �?      H@      ,@      �?              �?              B@      �?      N@                              @      3@      @@              @      5@      @      @      @      ,@     �W@      "@     �f@       @      �?      2@       @     �Y@      U@      �?      E@      &@      @      @              &@     �P@      @      h@      @       @      $@      @     �P@      A@      @      A@      &@      @      @              &@     �M@      @     �c@      @       @      "@      @      M@     �@@      @      A@      @      @      @               @     �D@      @     ``@      @       @      @      @      B@      :@      @      :@      �?                              @       @      @     �G@                      �?              @      @               @      @      @      @              @     �@@              U@      @       @      @      @      @@      4@      @      2@      @                              @      2@              :@      �?              @              6@      @               @      @                                      @               @                                      @                      @                                      @      ,@              2@      �?              @              2@      @               @                                              @              B@                      �?      �?       @      �?                                                              @              :@                      �?      �?      @      �?                                                              @              &@                      �?      �?      @      �?                                                                              .@                                      @                                                                                      $@                                      �?                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���WhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             !@�ŰzԒ�?�	           ��@       	                   �<@�����?�	           `�@                          �0@��u�@��?�           ��@                           �?�{���?�            �l@������������������������       �\9̜%�?O            �`@������������������������       ��q�ql�?=             X@                           @sdW�v��?I           �@������������������������       ��$v��j�?�           �@������������������������       ��١f!��?}           �@
                           �?^QB�1t�?�            `u@                           @YGn��m�?M            �`@������������������������       �6�>W[��?:             Y@������������������������       �\x ~�c�?            �@@                          @A@��4�[��?�             j@������������������������       �yַ���?x            �g@������������������������       �^Cy�5�?             3@������������������������       ���ZӼ��?             9@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      =@      B@      :@     @^@     ��@      @@      �@      (@      @      T@     @P@     ��@     �@      7@     �p@     �g@      =@      B@      :@     @^@     8�@      ?@     �@      (@      @      T@     @P@     ��@     �@      7@     �p@      f@      =@     �A@      :@     �Z@     ��@      ?@     ��@      "@      @     �R@     �N@     �@     �@      5@     �o@       @      �?      �?       @      "@     �B@      @     �F@      �?      �?      "@      @      =@      E@      �?      <@      @      �?      �?      �?      "@      2@      @      6@      �?      �?       @      @      1@      9@      �?      (@      @                      �?              3@              7@                      �?      @      (@      1@              0@      e@      <@      A@      8@     �X@     X�@      8@     @�@       @      @     @P@      K@      �@     �|@      4@      l@     �X@      @      4@      ,@     �I@     �p@      @     0{@      �?      �?      7@      5@     0s@      f@      @      Y@     �Q@      5@      ,@      $@     �G@     r@      3@     P}@      @      @      E@     �@@     u@     �q@      ,@     @_@      ,@              �?              ,@     �K@             �a@      @      �?      @      @      J@     �B@       @      (@      $@              �?              &@      &@             �L@       @              @      �?      *@      4@      �?      @       @              �?               @      &@             �G@       @              @      �?      @       @      �?      @       @                              @                      $@                                      @      (@                      @                              @      F@              U@      �?      �?      @      @     �C@      1@      �?      "@      @                              @      E@             �S@      �?      �?      @      @      =@      .@      �?      "@                                               @              @                                      $@       @                                                              (@      �?      @                                              @                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJg-�qhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?��(���?�	           ��@       	                    �?��tF�Y�?J           D�@                          �:@��H��w�?j           Ё@                           @~�6��w�?           �|@������������������������       ��G�u�?
           �z@������������������������       �[*�c
�?             ?@                          �=@�)�Ђh�?L            �[@������������������������       ��Z�R��?.            @Q@������������������������       �0,Tg��?             E@
                          �;@ȓWjD�?�           \�@                          �1@q\[�?�           �@������������������������       �U�{���?�            @n@������������������������       �D��G�?           ��@                          �<@����vg�?4            @U@������������������������       �     ��?             @@������������������������       ��bv�X��?!            �J@                            @�[y!��?L           �@                           @���W�?�           H�@                          �1@�ܻ�yX�?�           @�@������������������������       �:(�~�?>            �W@������������������������       �o?(�;V�?p           P�@                            �?��X�8�?           P�@������������������������       ��T�*�?�           Ȅ@������������������������       �z�"_7�?�             j@                           @V�~2���?�           0�@                          �4@@�T2��?            |@������������������������       �"����3�?�             j@������������������������       �0sKbCH�?�             n@                           �?�h�T�?g            �d@������������������������       �)O���?             2@������������������������       �
� :f��?W            @b@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@      >@      H@      @@      Z@     ��@     �D@     `�@      0@       @     �S@      O@     ��@     �~@      3@     �p@     �\@      0@     �@@      *@     �R@     �t@      7@     @x@      $@      @      E@      <@     @s@      k@      &@     �`@      A@       @      3@      @      2@      [@      @     �_@      @      �?      3@      @     @V@     �R@      @      J@      =@      @      .@      @      0@      W@       @      V@      @      �?      &@      @     �R@      Q@       @     �E@      <@      @      *@      @      .@     @V@       @      U@      @      �?      &@      @     �O@     @P@       @      C@      �?               @              �?      @              @                                      (@      @              @      @      @      @       @       @      0@      �?      C@                       @              ,@      @      �?      "@      �?      @      @       @      �?      "@      �?      7@                       @              @      @              @      @                              �?      @              .@                                      $@       @      �?       @      T@       @      ,@       @      L@     �k@      4@     `p@      @      @      7@      5@     `k@     �a@       @     @T@     @R@       @      (@       @     �K@      k@      4@     �l@      @      @      7@      5@      i@     �`@       @     @R@      0@      @      @              2@      K@       @     �@@              @      @      @     �A@      @@       @      4@     �L@      @      @       @     �B@     @d@      (@     `h@      @              3@      .@     �d@     �Y@      @     �J@      @               @              �?      @              A@                                      2@      "@               @      @               @                      @              (@                                      @                      @      @                              �?       @              6@                                      .@      "@              �?      Y@      ,@      .@      3@      >@     �t@      2@     ��@      @      @      B@      A@     �z@      q@       @     �`@     @T@      (@      $@      0@      :@     �m@      .@     �}@      @      @     �A@      :@     �q@      j@      @     �]@     �G@      @      @       @      &@     �X@      @     �h@      @              *@      (@     �b@      R@      @     �H@      &@                                      :@              7@                      �?       @      4@      @              @      B@      @      @       @      &@     @R@      @      f@      @              (@      $@      `@     @P@      @     �F@      A@      @      @       @      .@     �a@      (@     q@              @      6@      ,@     �`@      a@      @     @Q@      3@      @       @      @      $@     �Z@      @     `n@                      *@       @     �Z@     �Y@             �C@      .@      �?      @       @      @      A@      @      >@              @      "@      @      <@      A@      @      >@      3@       @      @      @      @     �W@      @     �o@      @              �?       @     �a@     �O@      �?      ,@      ,@      �?      @      @      @     �I@      @     @i@      �?                      @     �[@     �D@               @      "@              @      @      �?      ;@       @     @S@      �?                              M@      6@              @      @      �?      �?              @      8@      �?     @_@                              @     �J@      3@              @      @      �?                             �E@              I@       @              �?       @      ?@      6@      �?      @      �?                                       @              @                                       @      "@                      @      �?                             �D@              G@       @              �?       @      =@      *@      �?      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ3BwhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@����Ng�?�	           ��@       	                    �?�l2�w�?}           �@                           �?�=WQ>�?�           ؘ@                            @�F�4�D�?�            �m@������������������������       ��j])�S�?Z            `c@������������������������       ���1ʂ��?3            @T@                           @��~�vO�?S           (�@������������������������       ��>�$?�?:           �~@������������������������       �p�>T�L�?           �@
                           @�@���?�           @�@                            @:JNh���?�           T�@������������������������       �y�Sy�?s           �@������������������������       �]?n#k��?=            @                            �?"Q)Ho�?�            �w@������������������������       �6D3睠�?�            �j@������������������������       ��/�K.��?i            �d@                           �?��Iګ�?           0|@                            �?    �,�?�             p@                           �?C��H��?O            ``@������������������������       �AU� 9�?             �L@������������������������       ��_� ���?/            �R@                           �?�F ^�/�?O            @_@������������������������       �� �?            �I@������������������������       ������?1            �R@                           @�5�l��?}            `h@                           �?O���<�?p            �e@������������������������       �p�����?2            �R@������������������������       ��3�*��?>            �X@                           @؇���X�?             5@������������������������       ��<ݚ�?             "@������������������������       ��8��8��?             (@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      ;@      B@     �B@     �[@     (�@      ?@     ,�@      4@      $@     @P@      P@     ��@     �@      4@     @p@     �e@      6@      A@     �B@     �X@     ȁ@      >@     ��@      .@      @      K@      M@     Ѓ@     �}@      .@     �l@     �S@      ,@      <@      7@     �Q@     r@      3@     x@      *@      @      =@     �@@     �p@     �j@      &@      ]@      $@       @       @      �?      $@      :@      �?     �R@      @              @      @     �I@      5@              6@      @       @       @      �?      @      *@      �?     �H@      @              @      @      A@      *@              .@      @                              @      *@              9@                              �?      1@       @              @      Q@      (@      :@      6@      N@     pp@      2@     ps@      "@      @      7@      ;@     �j@      h@      &@     �W@      <@      @      $@      $@      3@      W@      (@      \@       @       @      @      @     �Q@     �U@       @     �@@      D@       @      0@      (@     �D@     `e@      @     �h@      @       @      3@      5@     �a@     �Z@      "@     �N@      X@       @      @      ,@      =@     �q@      &@     x�@       @      @      9@      9@      w@     �p@      @      \@     @S@      @      @      ,@      5@     �l@      "@     }@      �?      @      6@      3@     `s@     �k@      @     @U@      O@      @       @      &@      *@     `e@      @     �p@              @      5@      *@     �f@      e@      @     @P@      .@              �?      @       @     �M@       @     �h@      �?              �?      @      `@     �K@      �?      4@      3@      �?      @               @      I@       @     �c@      �?              @      @      N@     �D@              ;@      @      �?      �?              @      1@       @     �Z@      �?               @      @      B@      3@              1@      .@               @              @     �@@              J@                      �?      �?      8@      6@              $@      6@      @       @              (@      S@      �?     `c@      @      @      &@      @      V@      <@      @      @@      ,@      @       @              @      H@      �?     �U@      @      @      $@      @      A@      .@      @      5@      @      @       @               @      4@              A@                      $@              5@      *@              3@      @      @       @               @      @              &@                      $@              @      �?              *@       @                                      ,@              7@                                      1@      (@              @      "@                              @      <@      �?      J@      @      @              @      *@       @      @       @      @                               @      *@              ,@      @                      @      @      �?      �?               @                              �?      .@      �?      C@              @                      @      �?      @       @       @                              @      <@             @Q@       @              �?       @      K@      *@              &@       @                              @      <@             �I@       @              �?       @     �I@      *@              &@      @                              @      @              <@                                      0@      @               @      @                              @      5@              7@       @              �?       @     �A@      @              @                                                              2@                                      @                                                                                      @                                       @                                                                                      &@                                      �?                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�3ZhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @v��b�?�	           ��@       	                     �?Τ*����?�           R�@                           �?������?�           ��@                           @'b�z��?            |@������������������������       �t�E]t�?�            @s@������������������������       ��ݟ�ߦ�?b            �a@                           @�w?ȉ�?           P�@������������������������       ��q�=�r�?:           �~@������������������������       ���G-l�?E            �^@
                            �?~��`�7�?T           ��@                           �?w��V���?�           ܐ@������������������������       �{�G�N�?�             t@������������������������       ���K�6H�?�           ��@                           @�$����?�           0�@������������������������       �^#;���?;           Ѐ@������������������������       ��G�Z���?r            �e@                           @�p��!�?�           ��@                          �<@�r�{��?           H�@                           �?xN��/�?�           ؆@������������������������       �~��b)�?�            pu@������������������������       ���XD0��?�            @x@                          �=@l+�X�,�?1            �S@������������������������       ��0�~�4�?             6@������������������������       ��$I�$I�?$             L@                           �?�}/��I�?�            �n@                          �1@�(&����?]            `a@������������������������       �     @�?	             0@������������������������       ����%���?T            �^@                          �4@�5?,R�??             [@������������������������       ��8����?            �J@������������������������       �::P��P�?#            �K@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        f@     �A@      E@      <@     �X@     0�@      9@     ��@       @      @     @R@     �N@     ��@     p�@      1@     Pp@     �a@      6@     �@@      7@     �S@     �~@      5@     Ї@      @      @      P@     �I@     �@     �y@      ,@      l@      G@      $@      @      ,@      7@     �c@      "@     0w@      �?              1@      0@     �i@     �a@      @     �G@      2@      @      @      @      (@     �R@       @     @b@      �?              &@       @     �S@     �N@              =@      $@              @      @      "@      H@             �[@                      @      @     �J@     �A@              5@       @      @                      @      :@       @     �A@      �?              @      �?      9@      :@               @      <@      @       @      $@      &@      U@      @      l@                      @       @      `@      T@      @      2@      :@      @       @      @      @     @R@      @      e@                      @       @     @Z@     �P@      �?      &@       @                      @      @      &@             �L@                                      8@      *@       @      @     �W@      (@      <@      "@     �K@     �t@      (@     px@      @      @     �G@     �A@      s@     �p@      &@      f@     �I@      �?      2@      @      @@     �l@      @     pp@      �?              8@      1@     @i@     �`@      @      V@      0@      �?      $@      �?      ,@      L@             �R@      �?              0@      @      F@     �H@             �@@     �A@               @      @      2@     �e@      @     �g@                       @      *@     �c@     �U@      @     �K@     �E@      &@      $@      @      7@     �Y@      @      `@      @      @      7@      2@      Z@     �`@      @     @V@      C@      "@       @      @      2@     �S@      @     @X@      �?      @      1@      &@      T@      V@      @      S@      @       @       @              @      8@      �?      ?@       @              @      @      8@     �G@      @      *@     �B@      *@      "@      @      5@     `g@      @     pv@      @       @      "@      $@     @n@     �\@      @     �B@      ?@      @       @      @      2@     �`@      @     �q@      �?       @       @      @     �f@     �U@       @      >@      ;@      @       @      @      *@     �_@      @     `n@                       @      @     �e@     �U@              ;@      3@      @      @      �?      @      R@      @     @S@                      @      �?      V@     �E@              0@       @      �?       @      @      @      K@      �?     �d@                      @      @      U@     �E@              &@      @                              @      @             �E@      �?       @                      $@      �?       @      @                                               @              3@                                                              �?      @                              @      @              8@      �?       @                      $@      �?       @       @      @      @      �?              @      K@             @R@       @              �?      @      N@      <@      �?      @       @              �?              �?      ;@              L@                              @      >@      .@      �?      @                                      �?      @              "@                                                                       @              �?                      5@             �G@                              @      >@      .@      �?      @      @      @                       @      ;@              1@       @              �?      �?      >@      *@              @      @      @                       @       @              ,@                      �?      �?      (@       @              @              �?                              3@              @       @                              2@      &@              �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ/�khG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@z�,�c��?�	           ��@       	                    �?�v��?�           :�@                            @	�82�B�?�           ,�@                           �?��Б��?�           P�@������������������������       ��-8Hth�?M            �^@������������������������       ����\w�?~           Ȏ@                          �6@�_�hd�?           p{@������������������������       �_'��?�            pt@������������������������       �s
^N���?G             \@
                            @0�����?�           H�@                            �?�t�����?w           �@������������������������       ����i��?�           h�@������������������������       �3(&���?�             v@                           �?�1f ��?T           ��@������������������������       �݌��Ӏ�?�            0u@������������������������       �h������?{            �h@                            �?*�����?           �z@                           @�s8ޮM�?�            `m@                           �?2q�{��?l             e@������������������������       ���]^m�?>             W@������������������������       �2��k�?.             S@                          @@@�O��Ip�?+            �P@������������������������       ��!��}�?%            �L@������������������������       ���Q��?             $@                          �@@�a��"��?             h@                           �?l���s;�?s            `f@������������������������       ���0�*�?0            �R@������������������������       �ֻ���3�?C             Z@                           �?/����?             ,@������������������������       �      �?              @������������������������       �      �?             @�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      C@     �B@      =@      Z@     ��@      ?@     ܐ@      0@      @     @R@     �K@     ��@     �@      *@      p@     �g@      ;@     �A@      =@     �X@     (�@      ?@     Ќ@      (@      @      Q@      J@     h�@     �@      &@     @m@     �W@      *@      9@      .@      Q@     �s@      5@      t@      @      @      <@      7@     �q@      j@      @      _@      S@      @      1@      ,@     �J@     �k@      2@     �j@      @      @      8@      3@     �g@     `b@      @     @Y@      @      @      �?      �?      &@      .@      �?      =@       @              @       @      9@      @              .@     @Q@      @      0@      *@      E@     �i@      1@     �f@      @      @      4@      1@     `d@     �a@      @     �U@      3@      @       @      �?      .@     �V@      @      [@              �?      @      @     �W@     �N@              7@      $@      @      @      �?      *@      L@      @     �X@              �?      @      @     �Q@      C@              4@      "@      @      @               @     �A@              "@                                      8@      7@              @     @W@      ,@      $@      ,@      >@     �r@      $@     Ђ@      @       @      D@      =@     0w@     �r@      @     �[@     �S@      &@      $@      &@      :@     �l@      @     `x@      @       @     �B@      4@     �n@     @l@      @     @W@      J@      @      �?       @      4@     �e@      @     pt@      @              .@      *@     @i@     �d@      @     �K@      :@      @      "@      @      @     �L@             �O@      @       @      6@      @      F@     �N@      @      C@      .@      @              @      @     �Q@      @     �j@                      @      "@     @_@      R@              1@      "@                      @      @     �G@      @     �`@                      @      @      P@      I@              0@      @      @                              7@             �S@                               @     �N@      6@              �?      3@      &@       @              @     �U@             �c@      @      �?      @      @      Q@     �C@       @      8@      &@      &@      �?              @      H@             �P@       @              @      @      D@      ?@              ,@      &@      &@      �?              @     �C@              C@       @               @              =@      3@              *@      @      &@      �?              @      8@              8@                       @               @      @              @      @                                      .@              ,@       @                              5@      (@              @                                              "@              =@                       @      @      &@      (@              �?                                              @              =@                       @              &@       @              �?                                              @                                              @              @                       @              �?              @     �C@             �V@       @      �?      �?              <@       @       @      $@      @              �?              @     �C@              T@       @      �?      �?              9@       @       @      $@      @              �?                      ,@              >@      �?                              ,@      @              @                                      @      9@              I@      �?      �?      �?              &@      @       @      @      �?                                                      $@                                      @                                                                                      @                                       @                              �?                                                      @                                      �?                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJa΁;hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @n\`���?�	           ��@       	                     @\�ե���?-           ^�@                          �0@�ӈ��?l           ؛@                           @\��cy��?J            �_@������������������������       ���3@��?!            �M@������������������������       �\ͷ���?)            �P@                           �?�1��?"           ��@������������������������       �ޓ�݄P�?�           (�@������������������������       ���!����??           ��@
                          �4@��+J0�?�           ȅ@                           @�Z.��?�             r@������������������������       �[�Q}�D�?�            @h@������������������������       ���8��(�?A             X@                           �?Z��e8C�?�            py@������������������������       ��F���?y             h@������������������������       ��DS�T�?�            �j@                           �?�s1�l�?�           h�@                          �;@_>f|�?z           8�@                           @+���L�?Q           �@������������������������       ���3+ax�?           �y@������������������������       ��-���1�?A             Y@                           @ �Pm��?)            @Q@������������������������       �     ��?             0@������������������������       ���%�z�?            �J@                          �;@�oV.��?6           ��@                            @Qs>�E�?�           Ѕ@������������������������       �2�y�e��?\           �@������������������������       �
��U�z�?~            �f@                            @Z�_8-��?\             c@������������������������       �`Y�K�?@             Z@������������������������       �V�.��0�?            �H@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @i@     �@@     �D@      7@     �Z@     ��@     �@@     L�@      ?@      &@     �S@     �Q@     ��@     @�@      6@     q@     �a@      5@      B@      *@     @T@     @z@      0@     `�@      1@       @      E@     �D@     �}@     �q@      ,@      g@     �\@      1@      ;@      &@      O@     �t@      ,@     0{@      *@      @     �A@      ?@     �s@     �j@      ,@      b@      @      @      �?       @      @      <@      @      .@      @      �?      @              8@      ,@              0@                      �?               @      (@      @      @                      �?              4@      @              @      @      @               @      @      0@              "@      @      �?       @              @      @              $@     @[@      ,@      :@      "@      L@     �r@      $@     @z@      $@      @      @@      ?@     Pr@     �h@      ,@      `@     �F@      @      3@      @      C@     `a@      �?     �e@       @      @      *@      5@      _@     �U@       @      K@      P@       @      @      @      2@      d@      "@     �n@       @       @      3@      $@      e@     �[@      (@     �R@      ;@      @      "@       @      3@      W@       @      o@      @       @      @      $@     �c@     @R@              D@      .@       @      @       @      @     �D@             @S@                      @      @     @U@      @@              .@      $@              @       @      @      >@             �F@                      @      @     �J@      :@              *@      @       @                      @      &@              @@                       @              @@      @               @      (@       @      @              (@     �I@       @     �e@      @       @      �?      @      R@     �D@              9@      "@              @              "@      ?@       @     �F@      @                      �?      A@      ?@              5@      @       @                      @      4@             �_@               @      �?      @      C@      $@              @      N@      (@      @      $@      :@     �m@      1@     pz@      ,@      @      B@      >@     �l@     `m@       @      V@      ?@      "@      @      �?      "@     �X@      &@     `b@      "@      @       @      1@      U@     @Y@      @     �G@      ;@      "@      @      �?       @      W@      &@     @\@      "@      @      @      1@     �S@     �V@      @      D@      8@      "@      @      �?      @     �R@      $@     �U@      "@      @      @      0@     �M@     @S@      @      <@      @              �?              @      2@      �?      ;@                              �?      4@      ,@              (@      @                              �?      @              A@                      �?              @      $@      �?      @      �?                              �?       @              @                      �?              @              �?      @      @                                      @              ?@                                       @      $@              @      =@      @      �?      "@      1@     �a@      @     @q@      @              <@      *@      b@     �`@      @     �D@      =@      @      �?      "@      .@      Z@      @     �j@      @              :@      &@     �[@     @_@      @     �C@      5@      �?      �?      "@      (@     �R@      @     �a@      @              8@      "@     @U@     �V@       @      B@       @       @                      @      >@             �Q@                       @       @      :@      A@       @      @                                       @      B@              P@       @               @       @      A@      "@               @                                       @      *@             �H@                       @       @      ;@      @               @                                              7@              .@       @                              @       @                �t�bub�"     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�ϟhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@~���d��?�	           ��@       	                     @#�Zz���?s           B�@                            �?J���?           ��@                           �?`Nh���?j           �@������������������������       ���4�]�?�           �@������������������������       ��*�.)�?~           |�@                           @``Z+/��?�           ��@������������������������       ��4�B��?a           (�@������������������������       �F/.�?7            @V@
                           �?� �E>�?q           �@                           @
F<<�?           �{@������������������������       �DL#���?�            0s@������������������������       �iA� �?X            �a@                           @���5��?b           �@������������������������       ��N����?�            �u@������������������������       ��p?�[��?�            �h@                            @ӹ�	��?           �z@                          �=@#�� ���?�            �q@                           @
��@k�?Y            �`@������������������������       �s�n_Y��?D             Z@������������������������       ���L�*`�?             ?@                            �?�����?\            `b@������������������������       ��*Kf�?K             _@������������������������       ���Z�Y�?             7@                          �=@�>��3��?\            �a@                           @      �?'             P@������������������������       �      �?             H@������������������������       �     @�?             0@                          @@@8�Z$�?5            �S@������������������������       �QA�!��?$             K@������������������������       ���8��8�?             8@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @i@      C@      J@      7@     �W@     0�@     �@@     x�@      0@      "@      S@      N@     ��@     ��@      5@     `l@     �g@     �@@      I@      7@     @V@     ��@      =@     �@      *@       @     �P@      M@     0�@     �~@      3@     �i@     @d@      <@      ?@      4@     @Q@     �z@      5@     Ё@      &@      @      N@      H@      ~@     �w@      2@     �d@     �]@      5@      1@      0@     �F@     Pu@      0@     `}@      @      �?     �D@      =@     �v@     �o@      &@      [@      L@      $@      .@      @      7@     �b@      "@     �d@      @      �?      8@      .@      d@     �W@      @      N@      O@      &@       @      "@      6@     �g@      @      s@      �?              1@      ,@     �i@      d@      @      H@      F@      @      ,@      @      8@     �T@      @      Y@      @      @      3@      3@     �]@      `@      @      L@      B@      @       @      @      3@      R@      @      T@      @      @      2@      3@     �X@     �]@      @      H@       @              @      �?      @      &@              4@                      �?              4@      "@               @      <@      @      3@      @      4@     �f@       @     �t@       @       @      @      $@     �l@      [@      �?     �D@      *@      @      2@       @      ,@     �X@      @     @^@               @      @      �?     �U@      J@              ;@      (@      �?      2@              &@     �R@      @     �Q@               @      @      �?      M@     �B@              0@      �?       @               @      @      8@       @      I@                      �?              =@      .@              &@      .@       @      �?      �?      @     @U@      @     �i@       @              @      "@     �a@      L@      �?      ,@      "@      �?      �?      �?      @      G@             �`@       @               @      @     @Y@     �A@              &@      @      �?                       @     �C@      @     @R@                      �?      @      D@      5@      �?      @      (@      @       @              @     �Q@      @     �c@      @      �?      "@       @      V@     �D@       @      6@       @      @       @              @      D@      @     �V@      �?              "@      �?     @P@      A@              4@      @      @       @              �?      3@              A@                       @              A@      ,@              ,@      @      @       @              �?      &@              :@                       @              7@      *@              ,@      @                                       @               @                                      &@      �?                       @       @                       @      5@      @      L@      �?              �?      �?      ?@      4@              @               @                       @      4@       @     �F@      �?                              >@      1@              @       @                                      �?       @      &@                      �?      �?      �?      @              �?      @                              @      ?@             �P@       @      �?              �?      7@      @       @       @      @                                      (@              C@                                      @      @              �?      @                                      @             �@@                                      @      @                                                              @              @                                       @       @              �?      �?                              @      3@              <@       @      �?              �?      2@       @       @      �?      �?                               @      1@              *@       @                      �?      ,@       @       @                                              �?       @              .@              �?                      @                      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ%�@hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?<^1���?�	           ��@       	                    @ ���$�?F           l�@                           �?�5��*�?�           ��@                          �0@$���_��?W           h�@������������������������       �d�����?             3@������������������������       ��{�+P��?K           Ѐ@                            @��f��?�           ؐ@������������������������       ��dd�*�?           ��@������������������������       ��ܶ?Vr�?�            @l@
                            �? d��0u�?K             ^@                           �?0�����?             B@������������������������       ��q�q�?             "@������������������������       �d�ϙ�?             ;@                          �8@lv�"��?8             U@������������������������       �     H�?*             P@������������������������       ��G�z�?             4@                            @�A��?b           ܠ@                          �;@23���?�           $�@                            �?Lb;����?a           x�@������������������������       ��pi�� �?|           P�@������������������������       ��wS���?�            @w@                           @4��d6��?v            `e@������������������������       �����#�?O            @]@������������������������       ��6�3�?'             K@                           �?�d�́��?�           (�@                           �?�	,UP��?�             w@������������������������       �_�(6n�?<            �W@������������������������       ��A�S�?�             q@                          �2@\"�b���?�            �n@������������������������       ���b��?2            �S@������������������������       ����&Z�?h            �d@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@     �C@     �C@      >@      Z@     0�@      D@     8�@      6@      "@     �X@      M@     ��@     @~@      3@      q@      Y@      ;@      8@      3@     �O@      u@      2@     z@      1@       @      @@      >@     `t@     �g@      @     �a@     �V@      ;@      4@      3@      N@      t@      2@      x@      .@       @      @@      =@     �r@      f@      @      `@     �D@      0@      (@      "@      (@      Z@      @     �^@      $@      �?      0@      @      U@     �O@      �?     �M@                      �?                      �?                                      �?              @      $@               @     �D@      0@      &@      "@      (@     �Y@      @     �^@      $@      �?      .@      @      T@     �J@      �?     �L@      I@      &@       @      $@      H@     @k@      ,@     `p@      @      @      0@      :@     �j@     @\@      @     @Q@     �G@      @      @      "@     �A@     @e@      *@     @h@      @      @      .@      7@     `d@     @V@      @     �O@      @      @      �?      �?      *@      H@      �?      Q@                      �?      @      J@      8@              @      "@              @              @      ,@             �@@       @                      �?      ;@      .@              (@      @               @              @                      @                                      $@       @              @                                                              @                                      @                              @               @              @                      @                                      @       @              @       @               @                      ,@              :@       @                      �?      1@      *@              @       @               @                      *@              $@       @                      �?      0@      *@              @                                              �?              0@                                      �?                       @      X@      (@      .@      &@     �D@     `u@      6@     h�@      @      �?     �P@      <@     �x@     Pr@      (@     �`@     @R@      $@      "@       @     �A@      o@      4@     `z@      @      �?      O@      6@     q@     �m@      (@      [@      Q@      @      "@      @     �A@      k@      2@     �v@       @      �?      M@      2@      n@      l@      &@     �W@     �G@      @      @      @      1@     `e@      .@     �s@      �?              >@      @     �g@     @`@      @     �L@      5@      �?      @       @      2@     �F@      @     �H@      �?      �?      <@      &@      J@     �W@      @      C@      @      @              �?             �@@       @      M@      @              @      @      @@      (@      �?      *@      @      @              �?              7@       @      >@      @              �?      @      =@      @      �?      *@                                              $@              <@                      @      �?      @      "@                      7@       @      @      @      @     @W@       @     pp@                      @      @     �^@     �L@              8@      *@      �?      @      @      @     �F@       @     �c@                      @      @      P@     �E@              5@      @              @              �?      &@      �?      A@                                      ,@      .@               @       @      �?              @       @      A@      �?     @_@                      @      @      I@      <@              *@      $@      �?      �?              @      H@              Z@                      �?      �?     �M@      ,@              @      @                                      0@              ;@                      �?              8@      @                      @      �?      �?              @      @@             @S@                              �?     �A@      $@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ\�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�Bx         
                    �?0,��Rb�?�	           ��@       	                    !@�&�l�?M           X�@                          �=@%wO*
�?G           4�@                          �0@�!��?           �@������������������������       ��DXx_�?H            �\@������������������������       �`L����?�           L�@                            �?��L��?-            �Q@������������������������       ���M���?             A@������������������������       �/��.���?            �B@������������������������       �B{	�%��?             "@                            @��)e��?t           f�@                          �1@'w�g�?�           ��@                           @{u=49J�?�            �l@������������������������       �u�f�H �?`            �a@������������������������       ��t[p���?4            �U@                            �?��'`�P�?I           (�@������������������������       �L?܌��?~           <�@������������������������       ��Q.7�X�?�            �s@                           �?�)n��?�           (�@                           @*Mp���?@            �Y@������������������������       ��	"P7��?0             S@������������������������       ��1G����?             :@                           @ɉ�:��?W           ��@������������������������       �5&�3�?�            ps@������������������������       ����Kϟ�?�             m@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        l@      3@      @@      <@     �W@     @�@      C@     ��@      6@      "@     �P@      N@     ��@     ~@      :@     �m@     @^@      "@      6@      &@     �H@     �s@      6@      z@      1@      @      =@      ?@     �r@     @h@      &@     �`@     �]@      "@      6@      &@      H@     �s@      3@      z@      1@      @      =@      ?@     �r@     @h@      &@     ``@     �Z@      "@      6@      &@      E@     s@      3@     Px@      0@      @      =@      ?@     pr@      g@      $@     @`@      @              @              @      *@       @      1@      @              @      @      4@      2@      �?      &@     �Y@      "@      3@      &@     �A@     @r@      &@     @w@      (@      @      9@      :@     0q@     �d@      "@     �]@      &@                              @      @              ;@      �?                              @      $@      �?      �?       @                               @      �?              6@                                       @      @              �?      "@                              @      @              @      �?                              @      @      �?              @                              �?      �?      @                                                                      �?     �Y@      $@      $@      1@     �F@     �v@      0@     x�@      @       @      C@      =@     �|@     �q@      .@     �Z@     �U@      @      @      ,@     �E@      p@      (@     0|@      @       @     �B@      6@      t@     �j@      *@      W@      0@      �?      �?       @             �J@       @     �L@                      $@      @      =@      F@      �?      @      *@              �?                      C@       @      B@                      @      @      8@      *@              @      @      �?               @              .@              5@                      @      �?      @      ?@      �?      @     �Q@      @      @      (@     �E@     `i@      $@     �x@      @       @      ;@      1@     0r@     @e@      (@     @U@      E@      @      @      $@      6@     @f@       @     �s@      @              1@      &@     �l@      `@       @     �J@      =@               @       @      5@      9@       @     @S@      �?       @      $@      @     �N@     �D@      @      @@      0@      @      @      @       @     �[@      @     �p@                      �?      @      a@     @R@       @      .@      @               @              �?      6@      �?      >@                                      *@      4@              @      @               @              �?      1@      �?      7@                                      (@       @              @      �?                                      @              @                                      �?      (@                      "@      @      �?      @      �?     @V@      @     �m@                      �?      @      _@     �J@       @      "@      @      �?      �?      @      �?     �A@             �b@                      �?      @     �R@      >@              @      @       @                              K@      @     �V@                              �?      I@      7@       @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��{fhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @QL�ԙP�?�	           ��@       	                   �=@B�ED���?�           ��@                            �?�y�����?�           Ф@                            �?R|N��l�?�           ��@������������������������       �0�9���?o           ��@������������������������       ��:�ҍ��?�           ��@                          �1@�I{���?�           Ѓ@������������������������       �Z1x{���?W             `@������������������������       �$�Se��?G           �@
                            �?�э���?W            `b@                           �?:p�����?E            �]@������������������������       �EQEQ�?             E@������������������������       ������)�?,             S@                           �?
�b�m��?             =@������������������������       �      �?              @������������������������       �z'�L��?             5@                           �?�b_1��?�           8�@                           @����9�?6            @                           @�c��b�?�            �n@������������������������       ���|�'��?}            `i@������������������������       ���ճC��?             F@                          �9@��4ut��?�            `o@������������������������       ��:y��/�?}            �h@������������������������       �2+�QA�?             K@                           �?V��#�?           ��@                           @��Y3�M�?�            �x@������������������������       �rÄ��?�            �q@������������������������       ��P=���?C            �[@                          �>@	j*D��?�             j@������������������������       �v=m�ߧ�?�            @h@������������������������       �      �?             ,@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      =@      C@      ;@     �[@      �@      <@     H�@      (@      "@     �R@     �P@     @�@     �|@      *@     p@     �b@      5@      9@      7@     �V@     P~@      6@     ��@      "@      "@     @P@     �O@     @�@      v@      &@     �j@     �b@      4@      9@      7@     �U@     �|@      0@     ��@      @      "@      P@      N@     P@     �u@      &@      i@     @\@      0@      .@      6@      K@     pu@      ,@     (�@      @       @      D@      B@     �y@     `n@      @     �`@     �N@      @      @      1@      1@     �e@      "@     �t@                      (@      0@     �h@     �]@      @     �G@      J@      &@      $@      @     �B@     `e@      @     �o@      @       @      <@      4@     `j@     @_@      @     @U@      B@      @      $@      �?     �@@     �\@       @     @[@       @      @      8@      8@     @W@     �Y@      @     @Q@       @              @      �?      @      >@              (@              �?      @      "@      .@      6@       @      0@      <@      @      @              =@      U@       @     @X@       @      @      2@      .@     �S@      T@       @     �J@       @      �?                      @      <@      @     �O@      @              �?      @      3@      @              &@              �?                      @      :@      @     �F@      @              �?       @      3@      @              "@                                      @      @              8@                                      @      @              @              �?                              7@      @      5@      @              �?       @      ,@      �?              @       @                                       @       @      2@                              �?               @               @       @                                      �?              @                                               @                                                              �?       @      .@                              �?                               @     �G@       @      *@      @      5@     `g@      @     z@      @              $@      @      l@     �[@       @     �F@      =@      @      $@       @      0@     @T@      @      c@      @              "@       @     @W@     �O@              =@      (@       @       @       @       @      ?@       @     �R@       @              @             �H@      B@              0@      $@       @      @              @      :@       @     �P@       @              @             �E@      7@              *@       @              @       @      �?      @              @                       @              @      *@              @      1@      @       @               @      I@      �?     �S@      �?              @       @      F@      ;@              *@       @       @       @               @      G@      �?      J@      �?              @       @      C@      7@              $@      "@      �?                              @              ;@                                      @      @              @      2@      @      @       @      @     �Z@      @     �p@                      �?       @     ``@      H@       @      0@      *@      �?      @       @      @     �P@      @      f@                      �?       @     �R@      B@       @      *@      "@      �?      @       @      @     �@@      @     @`@                      �?       @      P@      :@              "@      @                                      A@              G@                                      $@      $@       @      @      @       @                       @     �C@              V@                                     �L@      (@              @      @       @                       @      C@              U@                                      H@      (@              @                                              �?              @                                      "@                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��uhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@2�;k܇�?�	           ��@       	                    �?��7U��?�           Z�@                            @eV�?1�?�           ̘@                            �?p��Ix�?�           ̑@������������������������       �u5H��?�            Pv@������������������������       �Ȱ����?�           p�@                           @�$I�$=�?            |@������������������������       ���lavW�?�            s@������������������������       ��1N�" �?Y            �a@
                            @/@�E��?�           �@                           @� �����?I           �@������������������������       ���#'�?w           ��@������������������������       �݊�6��?�           p�@                          �9@���9z�?Z           ��@������������������������       �5��}�?2           �~@������������������������       ��n���?(             R@                           �?�'���?           �y@                           @n�2&*�?q            `f@                           @�ue��?V            �`@������������������������       �H�N.���?>            @X@������������������������       �=J�L���?            �B@                          �=@\�D9�"�?            �F@������������������������       ��>4և��?             <@������������������������       �`3٫~�?
             1@                           @�R.���?�             m@                            @~��p��?�            �h@������������������������       ��X���?^            �`@������������������������       ��}j{3�?.            �P@                          �?@_��"�O�?             A@������������������������       �      �?             8@������������������������       �ףp=
��?             $@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@     �A@     �A@      6@      Z@     ��@      :@     �@      &@      "@     �Q@     �R@     ��@     �@      5@     q@     �f@      >@      A@      6@     �W@     ��@      9@     X�@      @       @     �O@     �Q@     `�@     �}@      2@      o@      X@      1@      9@      ,@     �J@     �s@      5@     pw@      @      @      =@      @@     @p@     �h@      "@     �`@     �R@      &@      ,@      ,@      E@      l@      0@     �o@      @      @      3@      >@     �d@      b@      "@     �[@      2@       @      @      @      &@      P@      @     �T@                      @       @     �P@     �N@       @      ;@     �L@      "@      &@      $@      ?@      d@      (@     @e@      @      @      ,@      6@      Y@     �T@      @     �T@      5@      @      &@              &@     @V@      @     �^@                      $@       @     �W@      K@              6@      .@       @      $@              "@     @Q@       @      Q@                       @             @Q@     �D@              (@      @      @      �?               @      4@      @     �K@                       @       @      9@      *@              $@      U@      *@      "@       @     �D@     �s@      @     ��@      �?      �?      A@     �C@     �x@     �q@      "@     @]@     @P@      $@       @      @     �B@     �k@      @     �v@      �?      �?      @@      ?@      p@     �j@      "@      X@     �E@      @      @      @      &@      X@             �d@                      $@      "@     �a@     @S@      @     �@@      6@      @      @       @      :@     @_@      @     �h@      �?      �?      6@      6@     @\@      a@      @     �O@      3@      @      �?       @      @     @X@      �?     �i@                       @       @      a@     �P@              5@      3@      @      �?       @       @     �V@      �?     �f@                       @       @      \@     �J@              2@                                       @      @              8@                                      8@      *@              @      0@      @      �?              $@     �Q@      �?     @c@      @      �?       @      @     @R@     �B@      @      8@      *@      @      �?              @      7@              M@                      @      �?      @@      6@      �?      ,@      (@      @      �?              @      2@             �C@                      @      �?      9@      &@      �?      (@      @      @      �?              @      0@              :@                      @      �?      2@      @      �?      &@      @                               @       @              *@                                      @      @              �?      �?                                      @              3@                                      @      &@               @                                              @              (@                                      @       @               @      �?                                                      @                                              "@                      @       @                      @      H@      �?      X@      @      �?      @      @     �D@      .@       @      $@      @       @                      @      A@      �?     �U@      �?      �?      @      @     �@@      .@       @      $@       @       @                      �?      1@      �?      K@      �?              @      @      8@      *@       @      "@      �?                               @      1@             �@@              �?                      "@       @              �?                                              ,@              "@      @                               @                                                                      "@              "@                                      @                                                                      @                      @                               @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJl �hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @B/Do�z�?�	           ��@       	                    @�_�����?           b�@                          �1@r��y���?;           ��@                           �?�;��KM�?�            �l@������������������������       �⃋��?T            �_@������������������������       �2�s�1�?D            @Y@                           �?ڼ�v���?�           �@������������������������       ������%�?7           @@������������������������       ��k��"e�?l           ��@
                          �<@������?�           �@                           �?b�r����?           ��@������������������������       ��	&q���?t             f@������������������������       �"����?           ��@                          �?@-��Y�"�?H            �Y@������������������������       ���>v��?-            �P@������������������������       �uk~X��?             B@                           �?*vW���?�           `�@                          �2@���Q��?�             t@                          �1@���-���?@            �W@������������������������       �333333�?             D@������������������������       ��#��M��?#            �K@                           �?��ӕ��?�             l@������������������������       ��������?             >@������������������������       �iOEA���?|            `h@                           �?bU&h���?�           ��@                           �?#��@���?!            �K@������������������������       �x9/���?	             ,@������������������������       �$E��~O�?            �D@                          �;@�<߮���?�           �@������������������������       ���<����?y           ��@������������������������       ��"��?@            �X@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@      ?@     �D@      :@     �X@     H�@      >@     `�@      2@       @      S@     �R@     `�@      @      5@     �m@     �c@      5@     �@@      4@      U@     �}@      :@     `�@      ,@      @     �Q@     �P@     ؀@     �w@      0@     �i@     �V@       @      9@      .@     �G@      m@      @     �t@      @      �?      ?@      <@     `p@     `a@      @      X@      7@      �?      @               @     �B@      @      F@                       @      *@     �G@      @@      �?      3@      &@      �?       @               @      0@      @      .@                      �?      @      >@      ;@      �?      ,@      (@               @                      5@              =@                      �?      "@      1@      @              @     �P@      @      5@      .@     �F@     �h@      �?     0r@      @      �?      =@      .@     �j@     �Z@      @     @S@      =@       @      1@      @      7@     �X@      �?     �_@      @      �?      4@      @     �T@     �F@      �?     �C@      C@      @      @       @      6@     �X@             �d@       @              "@      "@     �`@      O@       @      C@     �P@      *@       @      @     �B@     �n@      6@     �y@      "@      @      D@     �C@     Pq@     `n@      (@      [@     �P@      *@       @      @      B@     �l@      5@     �v@      @      @      C@     �C@     @p@      m@      (@     @Y@      $@                               @      3@      @     �K@      �?              @              C@      @@       @      @      L@      *@       @      @      <@     �j@      1@     ps@      @      @      A@     �C@     �k@      i@      $@     @X@                                      �?      .@      �?     �G@       @               @              1@      $@              @                                      �?      (@              ;@       @               @              ,@       @              @                                              @      �?      4@                                      @       @              �?      M@      $@       @      @      .@     @e@      @     �v@      @      @      @      @      n@      ]@      @      @@      *@      @      �?      @      @      J@       @     �W@                      @      @     �T@      F@              ,@      @              �?      @              2@              ?@                                      ?@      @              �?       @                                      "@              .@                                      &@      @                      �?              �?      @              "@              0@                                      4@      @              �?      $@      @                      @      A@       @     �O@                      @      @      J@     �B@              *@                                              @              @                                       @      ,@              �?      $@      @                      @      >@       @      N@                      @      @      F@      7@              (@     �F@      @      @      @      (@     �]@       @     �p@      @      @              @     �c@      R@      @      2@      @               @               @      @              ;@       @       @                      @      @                                       @               @                      @       @                                      �?                      @                                      @              4@               @                      @       @                     �D@      @      @      @      $@     �[@       @     `n@       @      �?              @      c@     @Q@      @      2@      =@      @      @      @      @     @X@       @     �h@      �?      �?              @      a@     @P@       @      0@      (@                              @      ,@              F@      �?                              .@      @      @       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJq�nkhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@M�T�{�?�	           ��@       	                     @=:����?�           �@                            �?�	J[)�?1           h�@                           @�m���?�           �@������������������������       ��/f�`�?y           ؕ@������������������������       ��y:m���?'           �|@                          �3@hw�H��?�           ��@������������������������       ��ӷ��?�            �o@������������������������       �f/�N�?�            pw@
                           �?����#�?a            �@                          �0@,V��a�?           �y@������������������������       �������?
             .@������������������������       �L?	�1�?           �x@                           @n���?S           H�@������������������������       ���m'��?           Pz@������������������������       �m0��2��?M            �`@                            @��@�F�?           }@                            �?�7<KQ�?�            �s@                          �?@i$��W�?I             ^@������������������������       ���c����?5            @V@������������������������       ��h70�?             ?@                          �=@�q�%�?t             h@������������������������       �     P�?;             X@������������������������       ��8��8~�?9             X@                           �?�Nh��
�?[             c@                           �?*L�9��?             6@������������������������       ��q�q�?             (@������������������������       ��Q����?             $@                           �?[!$��[�?L            ``@������������������������       �6��ѓ�?!            �M@������������������������       ����[���?+             R@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        l@      =@      H@      6@     @Y@     ��@      ?@     ��@      1@      @     �R@     �N@      �@     p@      .@     r@     `g@      ;@     �G@      6@     �V@     �@      =@     h�@      *@      @     �N@     �L@     ȃ@     �|@      ,@     �o@     �b@      1@     �D@      2@     @R@     z@      6@     ��@      $@      @     �G@      H@     `{@     �u@      (@     �j@     �Y@      *@      9@      0@     �G@     �u@      0@      �@      @              :@      <@     pu@      l@      @     �a@     �T@      @      4@      &@     �D@     0q@       @      y@      @              4@      6@     �o@      c@      @     �X@      5@       @      @      @      @     �Q@       @     �\@      �?              @      @     �V@      R@       @     �E@     �F@      @      0@       @      :@     �Q@      @     �[@      @      @      5@      4@     �W@      _@      @     �R@      3@       @      "@      �?      $@      B@      @     �F@              �?      (@      @      5@      C@      @      F@      :@       @      @      �?      0@     �A@      @     �P@      @       @      "@      *@     �R@     �U@      �?      >@     �C@      $@      @      @      2@     �c@      @     �u@      @              ,@      "@     `h@     �\@       @      D@      7@       @      @              .@     �R@      @     �]@      �?               @      @     @S@     �J@              5@      �?                                               @      �?                      �?      �?      @                      @      6@       @      @              .@     �R@       @     @]@      �?              @       @      R@     �J@              1@      0@       @      �?      @      @     @T@      @     �l@       @              @      @     �]@      O@       @      3@      $@       @      �?      @      @      Q@      @     �c@       @              @      @     �V@      I@       @      3@      @                                      *@             �Q@                      �?       @      <@      (@                      C@       @      �?              $@     �O@       @      f@      @      �?      *@      @     �R@      D@      �?      A@      :@       @      �?              @      E@       @     �X@       @              *@      @     �L@     �@@      �?      :@      �?                              @      3@              I@      �?              @      �?      6@      (@              @      �?                              @      1@             �B@      �?              @              1@       @              @                                               @              *@                              �?      @      $@                      9@       @      �?              @      7@       @      H@      �?              "@       @     �A@      5@      �?      3@      0@       @      �?                      .@              3@                      @       @      0@      *@              @      "@                              @       @       @      =@      �?              @              3@       @      �?      (@      (@                              @      5@             �S@       @      �?              �?      2@      @               @                                               @              "@                              �?       @      @              @                                                              @                              �?       @      �?              @                                               @              @                                               @                      (@                              @      3@             �Q@       @      �?                      0@      @              @      $@                               @      @              =@      �?                              @      @              @       @                               @      *@             �D@      �?      �?                      &@      �?                �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJp�hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @c��9c��?�	           ��@       	                    �?���?�           :�@                            �?F��H��?           �@                           @x�\���?           �|@������������������������       ����P�?�            �x@������������������������       �&�^YE��?&            �N@                            �?3x���?           ȉ@������������������������       �    0��?C            �@������������������������       ���&;��?�            �s@
                          �@@���;�}�?�           h�@                          �2@ìo��y�?�           (�@������������������������       �'P����?�            0w@������������������������       ����H&�?�           \�@������������������������       �      �?             0@                           �?����?�           ��@                          �;@]�����?�           x�@                          �9@���'�?[           `@������������������������       ���]����?8            |@������������������������       �$��m��?#             J@                          �@@��j�@u�?=            @V@������������������������       ��y���?5            �R@������������������������       �����S�?             ,@                           �?��u���?            �}@                           �?L�]B���?V            �a@������������������������       ����'F��?4            @T@������������������������       �N贁N�?"             N@                           �?��fG-B�?�             u@������������������������       ������?`             e@������������������������       ��ۓT"��?j            �d@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      ?@      D@      :@     @[@     ��@     �E@     ��@      8@      @     �Q@      R@      �@     �@      9@     �p@     �d@      4@      >@      9@     �U@     �}@     �B@     ��@      4@      @      O@      O@     �}@     �x@      7@     �l@      S@      ,@      7@      0@      M@     �k@      3@      q@      @       @      9@      ?@     `i@     �f@      (@     @^@      =@      �?      @      @      .@     �T@      $@     �^@                      *@      1@     �R@     �I@      @      ?@      8@      �?      @      @      (@     �P@      $@      X@                      *@      1@     �Q@      G@      @      >@      @                       @      @      .@              :@                                      @      @              �?     �G@      *@      4@      $@     �E@     `a@      "@      c@      @       @      (@      ,@      `@     @`@      "@     �V@     �@@      @      *@      @      >@     @W@      @     �Y@      @      �?      @      @      U@      Q@       @      K@      ,@      @      @      @      *@      G@      @      I@      @      �?      @       @      F@      O@      @      B@     �V@      @      @      "@      =@     `o@      2@     �|@      *@      @     �B@      ?@     0q@     �j@      &@     @[@     �V@      @      @      "@      =@     �n@      2@     �|@      *@      @     �B@      =@     �p@     �j@      &@     @[@     �D@      �?       @      �?      @      R@      @      V@                      (@      ,@     �K@      G@      @      =@     �H@      @      @       @      9@     �e@      .@     Pw@      *@      @      9@      .@     �j@     �d@       @      T@                                              @                                               @       @                              L@      &@      $@      �?      6@     �c@      @     �x@      @       @       @      $@     �l@     @]@       @      D@      C@      @       @      �?      $@     �P@      @     �m@      @       @       @      $@      [@     @Q@       @      8@      >@      @       @      �?       @     �M@      @     `g@       @      �?       @      "@     �X@     @P@      �?      6@      >@      @      @      �?      @      J@      @     �e@       @      �?       @      "@      T@     �L@      �?      4@               @       @              �?      @              (@                                      2@       @               @       @                               @       @             �I@      �?      �?              �?      $@      @      �?       @      @                               @       @             �C@      �?      �?              �?      "@      @      �?       @      �?                                                      (@                                      �?                              2@      @       @              (@     @V@       @     `c@      �?              @             �^@      H@              0@      *@      @                      @      3@             �@@                      @              E@      2@              @      $@      @                      �?      .@              &@                      @              6@      $@              @      @                               @      @              6@                                      4@       @              �?      @       @       @              "@     �Q@       @     �^@      �?              @              T@      >@              $@      �?      �?       @              @     �A@       @     �N@                       @              A@      0@               @      @      �?                       @     �A@             �N@      �?              �?              G@      ,@               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�"phG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@3Nb��x�?�	           ��@       	                     @�%{�]��?�           2�@                          �0@������?*           ��@                           @�
yW�?a             c@������������������������       ��ޔEǡ�?K            �]@������������������������       ��7�
t��?             A@                           �?����?�           x�@������������������������       �͔�?���?�           ��@������������������������       �d "�,�?4           l�@
                           @�Pi�aY�?m            �@                          �2@u��:���?           |@������������������������       �0_p��?V            `a@������������������������       �5�ԃ�E�?�            `s@                           �?����Sv�?U           �@������������������������       ��m��
�?�            �k@������������������������       �q�����?�            @r@                           �?7���B��?
            {@                          �=@�([bc�?�             o@                          �<@�*n��H�?E            @\@������������������������       ��Ĝ��?$             M@������������������������       �$�h���?!            �K@                           @G���U�?R             a@������������������������       ��q-�T�?<             Z@������������������������       �     ��?             @@                           @ڥ@G��?s            �f@                           �?SCp�j��?c            �c@������������������������       �0�����?/             R@������������������������       ��5;j��?4             U@                            �?�#*�6�?             ;@������������������������       ���S�ۿ?	             .@������������������������       ��q�q�?             (@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �i@      =@     �I@      1@      `@     ��@      =@     ��@      *@      @      V@     �P@     �@      ~@      1@     `m@     �g@      ;@     �E@      1@     @]@     ��@      =@     ��@       @      @     �R@      O@     (�@     `|@      .@      k@     �b@      .@     �A@      *@     �W@     �{@      5@     ��@       @      @     �P@      I@     0|@     �u@      ,@     �e@      &@       @      @       @      @      A@       @      3@                      @      @      8@      @@              @      "@       @      @       @      @      >@       @      .@                      @      @      2@      0@              @       @                              �?      @              @                                      @      0@              �?     @a@      *@      @@      &@      V@     �y@      3@     �@       @      @      O@     �E@     �z@     �s@      ,@      e@     @Q@       @      7@      @     �G@     �g@      &@     �j@      @      �?      9@      ;@     @f@      b@       @      Y@     @Q@      @      "@      @     �D@     �k@       @     �x@      �?       @     �B@      0@      o@      e@      @     @Q@      D@      (@       @      @      6@     �b@       @     t@                       @      (@     @l@     @[@      �?      E@      ,@      @      @       @      @      K@      @     �b@                      @      �?     �_@      I@              ;@      @              �?              �?      1@              D@                      �?             �J@      0@              @      "@      @      @       @      @     �B@      @      [@                      @      �?     @R@      A@              6@      :@       @       @       @      0@     @X@      @     �e@                      �?      &@      Y@     �M@      �?      .@      *@      @       @              $@     �K@      @      P@                      �?      @     �@@      :@              @      *@      @               @      @      E@      �?     @[@                              @     �P@     �@@      �?       @      0@       @       @              &@      N@             �e@      @      @      ,@      @      V@      :@       @      2@      .@       @       @              $@      D@              Y@              @      &@      @      ?@      *@       @      "@      @       @       @               @      7@              B@                      &@       @      (@      "@              @      @      �?                       @      (@              6@                      @               @      @               @              �?       @                      &@              ,@                      @       @      @      @              @      (@                               @      1@              P@              @              @      3@      @       @      @      $@                               @      $@             �J@              @               @      *@               @      @       @                                      @              &@                              �?      @      @              �?      �?                              �?      4@             �R@      @              @             �L@      *@              "@      �?                              �?      3@              J@      @              @             �J@      *@              "@      �?                              �?      @              ;@                                      8@      "@              @                                              0@              9@      @              @              =@      @               @                                              �?              6@                                      @                                                                                      ,@                                      �?                                                                      �?               @                                      @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�G�\hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �;@I�9���?�	           ��@       	                    @���\��?�           L�@                            @:}~}��?f           l�@                           !@�<m%��?Y           ��@������������������������       �e90z�?S           ��@������������������������       ���"e���?             "@                           �?�5��]�?           `�@������������������������       �M[��C�?�            �u@������������������������       ����z�r�?0           �~@
                           �?a����?:           ��@                          �7@ q�-Jl�?(           p|@������������������������       ��8��8K�?�             x@������������������������       �ۛ�3Q�?/            �Q@                          �4@HƵ�(�?           �z@������������������������       ��y>��?�            �n@������������������������       ���bi���?p            `f@                           �?l	�	O��?
           0z@                           �?ެ�Q�?.            �Q@                            �?     `�?             @@������������������������       ��P�n#�?	             1@������������������������       ��h$���?	             .@                           �?�(�	��?            �C@������������������������       ������H�?             "@������������������������       ���Wϊ�?             >@                            �?Mz�c��?�            �u@                            �?���u�?s            �f@������������������������       ������*�??             X@������������������������       ��s����?4             U@                           @LnR�-�?i             e@������������������������       �~ӝ�'#�?[            �b@������������������������       ��Q����?             4@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      ;@     �B@      4@     �W@     �@      C@     X�@      A@      @      X@      Q@     x�@     �@      4@     �n@     �h@      8@     �B@      3@      V@     �@     �B@     p�@      <@      @     @V@      O@     �@     �}@      *@     �l@      c@      2@      <@      .@      H@     �{@      >@     p�@      3@      @      O@      F@     ��@     �v@      @     �c@     �]@      (@      0@      *@      A@     �s@      9@     �y@      .@      �?     �I@      A@     @u@     �n@      @     ``@     �\@      (@      0@      *@      A@     �s@      6@     �y@      .@      �?     �I@      A@     @u@     �n@      @     ``@      @                                      �?      @                                                       @                      A@      @      (@       @      ,@      `@      @     `q@      @      @      &@      $@     @h@     �]@              9@      4@      @       @              $@      N@      @     @V@       @      @      @      �?     �T@      L@              "@      ,@       @      @       @      @      Q@       @     �g@       @              @      "@      \@      O@              0@      G@      @      "@      @      D@     ``@      @      p@      "@      �?      ;@      2@     `a@      [@      @      R@      6@       @      @      @      6@     �R@      @     �\@       @      �?      .@      (@      Q@     �L@      @     �C@      .@       @      @      @      5@     �P@      @     �Y@      @      �?      .@      (@     �I@     �G@      @      =@      @                              �?      @       @      *@      @                              1@      $@              $@      8@      @      @              2@     �L@             �a@      �?              (@      @     �Q@     �I@      @     �@@      5@              @              "@      A@             �U@      �?              "@      @      <@     �@@      @      0@      @      @                      "@      7@             �K@                      @      @     �E@      2@      �?      1@      6@      @              �?      @     @P@      �?      e@      @              @      @     �S@      ?@      @      2@      @      �?                              .@              4@                      @      @      &@       @              �?      @                                      $@              @                      @              @      �?                       @                                      @              �?                      @              @                              @                                      @              @                                      �?      �?                      �?      �?                              @              .@                              @      @      @              �?              �?                              �?              �?                              @       @      �?                      �?                                      @              ,@                                      @      @              �?      .@       @              �?      @      I@      �?     �b@      @               @      @     �P@      7@      @      1@      @       @              �?      @      :@              Q@      �?                      �?      F@      .@              "@                                      @      $@              F@      �?                      �?      ;@      @               @      @       @              �?      �?      0@              8@                                      1@      "@              @       @                                      8@      �?      T@      @               @       @      7@       @      @       @       @                                      5@      �?     @P@      @               @       @      5@       @      @       @                                              @              .@                                       @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��chG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @��mj��?�	           ��@       	                   �<@�i4�N#�?�           ��@                           �?N.���8�?h           �@                            �?�6D���?�             v@������������������������       �K0���o�?�             s@������������������������       �r�q�?              H@                           @2Q���9�?�           D�@������������������������       ��%�-��?|           Ȏ@������������������������       ��c�i?�?           $�@
                            �?JO�ݥ�?�            �j@                          �@@���_nw�?8            @W@������������������������       ����>4��?0             U@������������������������       ��2�tk~�?             "@                           �?�Ţ�B��?O            �]@������������������������       ����d;�?            �D@������������������������       �Z��Y���?2            �S@                          �2@Ƙ`F�?�           đ@                           @�?�Vc�?�            �q@                           �?&S���?�             i@������������������������       �r�q7�?=             X@������������������������       ��.y0���?I             Z@                           �?i�/���?3            @U@������������������������       �      �?              @������������������������       �K'"�/��?,            @S@                           �?��A`E��?           ��@                           @G����?�            �y@������������������������       ��&ih�?�             w@������������������������       �颋.���?             F@                          �4@���sT��?           `{@������������������������       �x9/���?:             U@������������������������       �Z�s���?�             v@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      C@      @@      3@     @Z@     �@      <@     Ȑ@      2@       @      X@     �L@     �@     ��@      9@     `q@     `e@      =@      6@      1@     �U@     0|@      7@     ��@      *@      @      S@     �F@     0@     �y@      9@     �l@     `c@      :@      5@      1@      U@     �z@      5@     H�@      *@      @      Q@     �E@     �|@      y@      7@      k@      6@       @      @      @      .@     �A@      @      W@      �?              *@             @S@     �H@      @      ?@      1@              @       @      ,@      =@      @     �U@                      $@             @Q@     �G@      @      5@      @       @      �?      �?      �?      @              @      �?              @               @       @       @      $@     �`@      8@      1@      ,@     @Q@     `x@      1@     �~@      (@      @     �K@     �E@     �w@     �u@      1@     @g@      R@      &@      .@      (@      A@     `h@      @     @l@      @              2@      .@      f@     �_@      @     �Q@     �N@      *@       @       @     �A@     `h@      (@     �p@      "@      @     �B@      <@     �i@      l@      *@     �\@      0@      @      �?              @      :@       @     �T@                       @       @     �C@      .@       @      (@                                       @      @      �?      H@                               @      4@      @              @                                       @      @      �?     �G@                                      4@      @              @                                               @              �?                               @              @              �?      0@      @      �?              �?      4@      �?     �A@                       @              3@       @       @      @       @       @      �?              �?       @              *@                      @               @      @               @       @      �?                              2@      �?      6@                       @              1@      @       @      @      J@      "@      $@       @      2@      h@      @     `y@      @       @      4@      (@     �m@      ]@             �H@      (@      �?      @      �?      @      H@      �?     �R@                      @       @     �U@      >@              (@      @              @      �?      @     �B@              I@                      @      �?     �Q@      *@              (@      �?              @              @      4@              :@                      @      �?      <@      @              @      @                      �?              1@              8@                                     �E@      $@              @      @      �?                       @      &@      �?      9@                      @      �?      0@      1@                                                       @      �?              @                                                                      @      �?                              $@      �?      4@                      @      �?      0@      1@                      D@       @      @      �?      *@      b@      @     �t@      @       @      *@      $@      c@     �U@             �B@      @@      @      @              (@      S@      @     `a@      �?              "@      @     �Q@      B@              7@      @@      @      @              @     @P@      @     ``@      �?              @      @     �P@      @@              1@              �?                      @      &@               @                      @              @      @              @       @      @       @      �?      �?      Q@      �?      h@      @       @      @      @     @T@      I@              ,@      @      �?      �?      �?              &@              <@       @               @       @      $@      1@              @      @      @      �?              �?     �L@      �?     �d@       @       @       @      @     �Q@     �@@              "@�t�bub�"     hhubh)��}�(hhhhhKhKhKhG        hh.hNhJP��rhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?� (cׄ�?�	           ��@       	                   �:@�e�>�?=           ��@                            @�|{\[�?�           $�@                            �?����?�           D�@������������������������       ��q,:�?�            0v@������������������������       ��玜��?�           p�@                           @�t�V� �?	           �w@������������������������       ��
t�Fp�?�             q@������������������������       �R�}e�.�?I             Z@
                           �?.Bm����?�            �l@                           �?�3�kf�?H            @[@������������������������       �"pc�
�?             F@������������������������       �mI����?-            @P@                          �>@�!�`��?I            �^@������������������������       �(vb'vb�?<             Z@������������������������       ��Kh/���?             2@                          �<@���� ��?z           2�@                            @ॼ�(��?�           4�@                            �?c�%O{�?�           ��@������������������������       ��՘b��?�           T�@������������������������       �W 
I��?�            �t@                          �9@����t��?X           P�@������������������������       �o[�(���?.           �~@������������������������       ������?*            �P@                            �?�����?�            �i@                           @ŏ1w-�?E             Y@������������������������       ��X����?<             V@������������������������       ��������?	             (@                           �?�q-�??             Z@������������������������       �r-�T��?!             J@������������������������       ��}e�.y�?             J@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@      ?@     �D@     �@@     �Z@     H�@      @@     \�@      2@      &@     �V@     �I@     ��@     @      .@     `p@     �Y@      2@      =@      *@      N@     `s@      1@     @y@      (@      @      F@      >@     Pr@     @l@      @     �a@     @U@      .@      <@      &@     �J@     �q@      1@     �s@      $@      @      B@      =@     p@      i@      @     �_@     �Q@      (@      8@      &@     �E@     @j@      ,@     �j@      "@      @      >@      <@     @f@     �b@      @     �Y@      4@       @      @      �?      .@     �N@       @     �U@                      @      ,@     @P@     �H@       @      <@     �I@      $@      3@      $@      <@     �b@      (@     �_@      "@      @      9@      ,@     @\@      Y@      @     �R@      ,@      @      @              $@     �R@      @     �Z@      �?              @      �?     �S@     �I@              8@      *@       @      @               @      M@       @     �P@      �?              @      �?     �J@      C@              6@      �?      �?                       @      0@      �?     �C@                      @              :@      *@               @      2@      @      �?       @      @      :@             @U@       @               @      �?      B@      :@              0@      *@      @      �?       @      @      ,@             �E@                       @      �?      "@      @              @                               @       @      @              5@                      @      �?      @                       @      *@      @      �?               @       @              6@                       @              @      @              @      @                              @      (@              E@       @                              ;@      5@              $@      @                              @      (@             �@@       @                              9@      0@              $@       @                                                      "@                                       @      @                     @X@      *@      (@      4@     �G@     0u@      .@     �@      @      @     �G@      5@     p}@     �p@      $@     �]@     @V@      *@      (@      4@     �F@     �r@      ,@     p�@       @      @     �D@      5@      {@     pp@       @      [@     �R@       @      "@      0@     �D@      l@      $@     �x@      �?      @      C@      .@      s@      j@      @     �V@     �K@      @      @      *@      7@     �f@      "@     �t@      �?              5@      (@     �n@     �b@      @     �M@      3@       @      @      @      2@      E@      �?      P@              @      1@      @      O@      N@      @      ?@      .@      @      @      @      @     @S@      @     �l@      �?              @      @      `@      K@       @      2@      .@      @      @      @      @     @P@      @     @j@      �?              @      @     �Y@     �G@       @      0@                                              (@              4@                                      9@      @               @       @                               @     �B@      �?     @U@      @      @      @             �B@       @       @      &@      @                                      5@      �?      @@                      �?              6@       @              "@      @                                      4@      �?      6@                      �?              5@       @              "@                                              �?              $@                                      �?                               @                               @      0@             �J@      @      @      @              .@               @       @                                               @              @@              @                      @               @      �?       @                               @       @              5@      @              @              "@                      �?�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�I�OhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @���z�?�	           ��@       	                   �<@%��[���?            �@                            �?0�?u           R�@                           @�v�x¸�?�           8�@������������������������       �i�7b1��?2           Ћ@������������������������       ���2�	��?�           P�@                           �?�H���?�           ؄@������������������������       �-�Q���?J            �_@������������������������       ��h�P,f�?^           �@
                          �@@8֊Hp��?�            �k@                           �?���qE�?{            �g@������������������������       ��[��?            �B@������������������������       �0���%��?b            @c@                           @F#߼��?             >@������������������������       ������?
             7@������������������������       �������?             @                           @�[����?�           �@                          �7@�P���s�?�           (�@                           �?�I��?<           @~@������������������������       �m��1��?�             j@������������������������       �y��`���?�            @q@                           �?v��^�?�            r@������������������������       �rz׾��?G            �]@������������������������       �?��hq�?k            `e@                           �?vT+��n�?�            �s@                          �<@�T����?f            �d@������������������������       �#2��0��?^            `b@������������������������       ���Kh/�?             2@                           @'D(~�)�?_             c@������������������������       �3��b���?6            �V@������������������������       �a��V{q�?)             O@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �f@      6@      B@      =@     �[@     ��@     �A@     ��@      6@      @      R@     �O@     ��@     ��@      :@     �p@     �a@      2@      9@      4@     @U@     0}@      <@     І@      5@      @      P@      L@     p@     �y@      6@      l@     �`@      2@      8@      4@     �T@     �z@      :@      �@      0@      @      M@      I@      }@      y@      5@     �j@     �Y@      @      ,@      2@      N@     �u@      5@     �@      &@      �?     �A@      8@     �u@     �q@      .@     �a@      J@      @      $@      &@     �@@     �e@      @     �o@       @              1@       @     �c@     �Y@      @     �K@      I@      @      @      @      ;@      f@      0@      p@      @      �?      2@      0@     �g@     �f@      $@     @U@      ?@      &@      $@       @      6@      S@      @     �`@      @       @      7@      :@     �^@     �]@      @     �R@      @      @      @              @      (@              2@      @              @      @      =@      *@      @      5@      <@      @      @       @      .@      P@      @      ]@      �?       @      4@      7@     @W@     @Z@      @     �J@      "@              �?              @     �E@       @     �U@      @              @      @     �B@      (@      �?      $@      "@              �?              @      A@       @     @T@      @              @      @      <@       @      �?       @      �?                                      $@              2@                       @       @       @      �?              �?       @              �?              @      8@       @     �O@      @              @      @      :@      @      �?      @                                              "@              @                              �?      "@      @               @                                               @              @                                      "@                       @                                              �?              �?                              �?              @                     �D@      @      &@      "@      9@     @h@      @     �x@      �?       @       @      @     �k@      ]@      @     �F@     �@@       @      $@      @      1@     @b@      @     @p@               @       @      @      b@     @X@      @      B@      5@       @      $@      @      "@     @W@      @     @b@               @       @      @      U@     @Q@       @      <@      "@      �?      @              "@      E@              G@               @      �?      @      ;@      F@              1@      (@      �?      @      @             �I@      @      Y@                      �?       @     �L@      9@       @      &@      (@                               @     �J@       @     �\@                              �?     �N@      <@       @       @      "@                              @      8@       @      A@                                      9@      1@       @      �?      @                              @      =@              T@                              �?      B@      &@              @       @       @      �?       @       @      H@      �?     �`@      �?              @      �?     @S@      3@              "@      @       @      �?       @      @      ;@      �?      L@                      @             �E@      &@              @      @       @      �?       @      @      ;@      �?      G@                      @              B@      $@              @                                                              $@                                      @      �?                      @                               @      5@             �S@      �?              �?      �?      A@       @              @      @                               @      @              J@                              �?      :@      @              �?                                              2@              ;@      �?              �?               @      @               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ
Ȳ%hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @~����?�	           ��@       	                   �0@_͌��?�           ��@                            �?ŕ`�|�?p            �g@                           @ԛ����?*            �R@������������������������       �c�=yX�?             I@������������������������       �j�t��?             9@                           �?C�/`?F�?F            �\@������������������������       �p��G��?            �E@������������������������       ��Kh/��?.             R@
                           !@l`�k*��?Y           4�@                           �?�lϕ���?R           �@������������������������       ��aCg?f�?�           0�@������������������������       ��T"f�?�           �@������������������������       �����W�?             *@                           �?��SO� �?�           đ@                          �=@�r��-�?B           �@                           @��DRJ��?+           �~@������������������������       �0	x]�?�            Pt@������������������������       ���7��?e             e@                           �?�>d?�?�?            �G@������������������������       �r�q��?             (@������������������������       �^�{�X�?            �A@                           �?FR�����?�           ��@                          �2@�(\��u�?9             T@������������������������       ������?             3@������������������������       �)���G��?+            �N@                           @n?��{��?L            �@������������������������       �0i��?�?�            �l@������������������������       ���l��(�?�            �q@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       @l@      C@     �A@      7@      X@     ��@      C@     �@      4@       @     �P@     �N@     ��@     @      8@     �o@      e@      6@      <@      4@      S@     @}@      >@     Ȅ@      .@      @     �M@      H@     x�@     �w@      5@     �j@       @              @       @      @      C@       @      0@      �?       @      @       @     �E@     �B@              6@      �?                      �?      @      ,@              &@                                      0@      3@              "@                              �?      @      @               @                                      0@      0@              @      �?                                      $@              "@                                              @               @      @              @      �?      @      8@       @      @      �?       @      @       @      ;@      2@              *@                      @               @      @              @      �?              @      �?      &@      $@               @      @                      �?      �?      3@       @       @               @       @      �?      0@       @              &@      d@      6@      9@      2@     @Q@     �z@      <@     H�@      ,@      @      J@      G@      �@     Pu@      5@      h@     �c@      6@      9@      2@     @Q@     �z@      6@     0�@      ,@      @      J@      G@     �@     Pu@      5@      h@     �S@      "@      5@      @     �E@     �i@      (@      n@      @       @      4@      ;@     �g@     �a@      "@     �V@      T@      *@      @      (@      :@     �k@      $@     `y@      "@      �?      @@      3@     pt@     �h@      (@     �Y@      �?                                       @      @      @                                      �?                              M@      0@      @      @      4@      h@       @      z@      @      @       @      *@     @l@     �]@      @      C@      C@      @      @      �?      *@     �X@      @      e@      @       @      @      "@     @X@     @P@       @      6@      9@      @      @      �?      &@     �V@      @      d@      @       @      @      @      V@     @P@              4@      6@      @      @      �?      @     �Q@      @     �T@                      @             �Q@      F@              .@      @      @      �?              @      4@      @     @S@      @       @              @      2@      5@              @      *@                               @      @              "@      �?                       @      "@               @       @                                      �?       @                      �?                       @      @                              *@                              �?      @              "@                                      @               @       @      4@      "@       @       @      @     �W@       @      o@      �?      �?      @      @      `@      K@      �?      0@      @               @              @      &@              A@                                      "@      @              @                                      @                      $@                                      �?      �?              @      @               @              �?      &@              8@                                       @      @              @      ,@      "@               @       @     �T@       @     �j@      �?      �?      @      @      ^@     �G@      �?      $@      @                      �?      �?      6@              Y@              �?      @      �?     �R@      1@              @      "@      "@              �?      �?     �N@       @     �\@      �?               @      @      G@      >@      �?      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJDH]\hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @�/��j�?�	           ��@       	                    @���(��?�           �@                          �4@d֑����?U           �@                            �?�|���+�?�           ��@������������������������       �mR�u���?0           ��@������������������������       ��H����?�            �t@                            �?^�!����?W           (�@������������������������       �������?V           ��@������������������������       ��X�R~��?           ��@
                            �?W�%�(V�?�            Pp@                          �;@������?C            �X@������������������������       ����Q8�?6             T@������������������������       ��GcT!)�?             3@                            �?��*���?d            @d@������������������������       ��sٞ��?A            �Z@������������������������       ����>4��?#             L@                           �?�#ve��?�           L�@                           @�0�_���?v             h@                           �?��eTs��?[            �b@������������������������       ���I!��?)            �R@������������������������       �D�.�?2            @S@                          �:@�e�J��?             E@������������������������       �     ��?             @@������������������������       �p=
ףp�?             $@                           �?�P5�R��?E           ��@                           �?}�L|�t�?�            �w@������������������������       �����4��?_             `@������������������������       �<㽀4��?�            �o@                          �2@�Dٴ��?L           ��@������������������������       ���� m�?P            �`@������������������������       �Վ�%��?�            �x@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �e@     �C@     �C@      5@     �X@     ��@      E@     ��@      2@      &@     �T@      J@     x�@      �@      1@     Pp@     �a@      <@      @@      1@     @T@      ~@     �C@      �@      .@      $@     @R@      D@     �@     Pw@      0@     �j@     �`@      :@      :@      .@     @S@     �{@     �@@     ؃@      ,@      $@     �P@     �A@     �}@     `u@      0@     �h@     �R@      *@      .@      @      C@      m@      .@     �p@      @      @      ?@      3@     `g@      h@      $@      U@     �K@       @      *@      @      8@      f@      &@     �k@      @       @      1@      "@     @a@     �`@      @      E@      4@      @       @              ,@     �K@      @      G@               @      ,@      $@     �H@      N@      @      E@     �M@      *@      &@      &@     �C@     `j@      2@     �v@      &@      @     �A@      0@     r@     �b@      @     @\@      <@      @      �?       @       @      X@      *@      e@      @              @      @      [@     �J@      @      =@      ?@      "@      $@      @      ?@     �\@      @     �h@       @      @      <@      $@     �f@      X@      @      U@      "@       @      @       @      @     �C@      @     @Y@      �?              @      @      ?@      ?@              1@      @       @      @       @       @      *@      @      <@      �?                      @      2@      ,@              @      @       @      @       @       @      (@      @      4@      �?                              (@      ,@              @                                              �?               @                              @      @                      �?      @              @               @      :@      @     @R@                      @       @      *@      1@              &@      �?                               @      ,@      @     �K@                      �?       @      (@      $@              @      @              @                      (@              2@                      @              �?      @              @      >@      &@      @      @      1@     �f@      @     �x@      @      �?      $@      (@     �n@     `a@      �?     �G@      @              �?              @     �A@             �L@                              �?     �C@      B@              *@      @              �?              @      =@             �D@                              �?     �@@      7@              *@      �?              �?              @      2@              1@                                      (@      ,@               @      @                              @      &@              8@                              �?      5@      "@              @      �?                                      @              0@                                      @      *@                      �?                                      @              "@                                      @      &@                                                              �?              @                                               @                      9@      &@      @      @      &@     `b@      @     0u@      @      �?      $@      &@     �i@     �Y@      �?      A@      3@      @      @       @      "@      M@      @     �Z@       @              @      @     �S@      K@      �?      8@      $@       @       @              �?      :@       @      5@                      @             �A@      0@               @      "@      @      @       @       @      @@      �?     �U@       @              �?      @      F@      C@      �?      0@      @      @               @       @     @V@              m@      �?      �?      @       @     �_@     �H@              $@       @                       @              5@              G@                      �?       @      G@      ,@              �?      @      @                       @      Q@             @g@      �?      �?       @      @      T@     �A@              "@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJK	 hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             @w{�k�?�	           ��@       	                    �?&��(M`�?M           �@                           @��i���?U           �@                           @��gs�?�           ��@������������������������       ��r��?�           ��@������������������������       �������?           �z@                           @�Q�w^��?}            �h@������������������������       �H6$ ��?;            @U@������������������������       �Y��fC��?B            �[@
                           �?�����?�            �@                          �;@Ӣv�-�?�           �@������������������������       �uԂ�a�?�           �@������������������������       ���8��X�?@             X@                          �2@cu��F�?,           0�@������������������������       �� ��r��?�            s@������������������������       �2�{ ���?j           ��@                            �?��'D�h�?f           ��@                           �?�!J[���?�            �n@                           @xX�L�?=            �W@������������������������       �窷uJ��?(            �L@������������������������       ���!CA[�?            �B@                           �?~�+r��?`             c@������������������������       ��KM�]�?             3@������������������������       �`@����?R            �`@                          �:@~'�£��?�           @�@                            @>(o����?o           �@������������������������       ���u�b�?�            �w@������������������������       ��W��٭�?w            `h@                           @�z���?Z            `a@������������������������       �8��P��?H            �\@������������������������       �9��8���?             8@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        i@      5@      D@      ;@      [@     h�@      >@     ԑ@      6@      @     �R@      L@      �@     �@      3@     �p@     @c@      *@      >@      8@     �W@     �@      0@     h�@      1@       @      L@      E@     X�@     `u@      *@      k@      S@       @      5@      2@     �O@      n@       @      u@      (@      �?      B@      ,@     �m@     �c@      @     �[@     �N@      @      5@      .@     �L@     @k@      @     `q@      &@      �?      8@      ,@     @j@     �`@      @     @V@     �B@       @      0@      $@      A@     �b@       @     `e@      @              2@      @      \@     �W@      @     �M@      8@      @      @      @      7@     @Q@      @     �Z@      @      �?      @      @     �X@     �C@      @      >@      .@      @              @      @      6@       @      N@      �?              (@              ;@      7@              6@      "@      �?              @      @      *@       @      ,@                      @              (@      &@              *@      @       @                      @      "@              G@      �?               @              .@      (@              "@     �S@      @      "@      @      ?@     �p@       @     ؀@      @      �?      4@      <@     �s@      g@      @     @Z@      E@      @      �?      @      3@     @^@      @     �l@              �?      "@      3@      a@     �T@      @     �O@     �D@      @      �?      @      2@     @Y@       @     @g@                      "@      1@     @_@     �T@             �J@      �?      �?                      �?      4@       @     �E@              �?               @      &@      �?      @      $@      B@               @      @      (@     �a@      @     `s@      @              &@      "@     �f@     �Y@      @      E@      5@              �?      �?      �?     �K@      �?     �W@                      @      @     �Q@      ?@       @      (@      .@              @       @      &@      V@      @     �j@      @              @       @     �[@     �Q@      �?      >@      G@       @      $@      @      ,@     �b@      ,@     �p@      @      @      2@      ,@     �f@     �e@      @      I@      &@      @      @      @      @      7@      �?     @R@                      @              N@     �F@              (@      @       @      @              @      $@              ;@                                      3@      .@              &@      @       @      �?                      @              4@                                      @      ,@              @                      @              @      @              @                                      .@      �?              @       @       @              @      �?      *@      �?      G@                      @             �D@      >@              �?                              �?      �?      �?      �?       @                      @               @      �?                       @       @               @              (@              C@                       @             �C@      =@              �?     �A@      @      @              $@     �_@      *@     �g@      @      @      (@      ,@     @^@      `@      @      C@      >@      @      @              $@     @Y@      (@      `@      @       @      (@      ,@     �W@     @\@      @      A@      7@      �?      @              @     �P@      &@     �Q@      @      �?      "@      "@     �K@     �S@      @      @@      @      @       @              @      A@      �?     �M@              �?      @      @      D@      A@               @      @                                      9@      �?      O@              �?                      :@      .@              @      @                                      4@              L@              �?                      3@      ,@                                                              @      �?      @                                      @      �?              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJM�B^hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @he"����?�	           ��@       	                   �0@��d���?           @�@                           �?�1xP�1�?x            �f@                           �?�(�!N�?7            �U@������������������������       �l	��g��?              I@������������������������       ��[��?            �B@                           @�-�)8D�?A            �W@������������������������       ��]�l�?             A@������������������������       ����h��?*            �N@
                           �?�zw�?�           Ԥ@                           @�	3Z"��?�           �@������������������������       ���b���?�           ��@������������������������       �
^N��)�?	             ,@                           �?-[jI(~�?�           ��@������������������������       ��t�@��?           �y@������������������������       �h���)c�?�           T�@                           @�qQR��?�           ��@                           �?G�n-�q�?0           p}@                           �?$I�$I�?�             l@������������������������       �ms�z�?            �G@������������������������       �T��k�V�?y             f@                          �0@���d�?�            �n@������������������������       �      �?              @������������������������       ���&�ѣ�?�            �m@                          �:@̖����?}           ��@                           @)�=9��?4           �~@������������������������       �x�@���?t             f@������������������������       �YV7E��?�            ps@                           @��2tm�?I            �Z@������������������������       �g\�5�?             :@������������������������       ��������?7             T@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �h@      @@     �G@     �@@      Z@     h�@      D@     h�@      3@      @     �U@     �T@     ��@     8�@      3@     �m@      c@      5@     �B@      ;@     �U@     �|@      ?@     ��@      (@      @      S@      Q@     ��@     pz@      2@     �h@      @      �?      �?      @      ,@      D@      @      8@      �?              @      @      >@      C@              *@      �?      �?      �?      �?      $@      9@       @      "@      �?              �?      @      &@      4@              �?              �?      �?      �?      $@      @       @      @      �?              �?               @      *@                      �?                                      3@              @                              @      @      @              �?      @                       @      @      .@      �?      .@                      @      �?      3@      2@              (@                                              @              �?                                      *@      (@              @      @                       @      @      &@      �?      ,@                      @      �?      @      @               @     @b@      4@      B@      8@      R@     `z@      <@     8�@      &@      @      R@      P@      @     x@      2@     @g@     @Q@      &@      6@      &@      E@     �g@      ,@     @o@      $@      @     �C@      =@     �h@      d@      @     �V@     @Q@      &@      6@      &@     �D@     �g@      $@      o@      $@      @     �C@      =@     �h@     `c@      @     �V@                                      �?       @      @      �?                                      �?      @                     @S@      "@      ,@      *@      >@     �l@      ,@     �z@      �?             �@@     �A@     �r@      l@      (@      X@      A@              @       @       @     �K@             �X@                      @      ,@     @Y@     �N@       @      :@     �E@      "@      &@      &@      6@      f@      ,@     �t@      �?              <@      5@     �h@     �d@      $@     �Q@     �G@      &@      $@      @      2@     �g@      "@     �u@      @      �?      $@      ,@      l@      `@      �?      D@      6@      �?      @      @      $@     @R@      @     `c@       @      �?      @       @      \@     �G@              9@      1@      �?      @      @       @      C@      @     �K@       @              @      �?     �F@      7@              0@       @                               @      $@              1@                      �?              @      @              @      .@      �?      @      @      @      <@      @      C@       @              @      �?     �C@      2@              (@      @              �?       @       @     �A@              Y@              �?              �?     �P@      8@              "@                                                              @                                      �?                              @              �?       @       @     �A@             @W@              �?              �?     �P@      8@              "@      9@      $@      @      �?       @     �]@      @      h@      @              @      (@     @\@     @T@      �?      .@      6@       @      @      �?       @      V@      @     �b@                      @      (@      X@     �S@              (@      "@      @              �?      @     �E@              H@                              @      B@      6@              @      *@      @      @               @     �F@      @     �Y@                      @       @      N@      L@              @      @       @                              >@              E@      @                              1@      @      �?      @      �?                                      &@              $@                                      �?       @              �?       @       @                              3@              @@      @                              0@      �?      �?       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ5u�9hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                              @���E��?�	           ��@       	                   �1@�2��?�           ��@                           �?
_؋x��?           0{@                          �0@�p� �?�            �m@������������������������       �^�;#1r�?A            @X@������������������������       �^�G���?U            `a@                           �?��DS_F�?�            �h@������������������������       ��o�����?             ;@������������������������       ��������?v            �e@
                            �?�)�����?�           ��@                           �?ݒ�;d�?T           ��@������������������������       ��^��8��?�           Ȉ@������������������������       ��2� ��?q           ��@                          �;@}�پt��?u           �@������������������������       ���D����?T           (�@������������������������       �����S�?!             L@                           �?X'I:|7�?�           <�@                          �>@A߲�L�?D           `@                          �=@��|�`�?8           ~@������������������������       ��먥�R�?2           �}@������������������������       �      �?              @������������������������       �e�J��?             5@                          �2@`��e�?�           Ȃ@                           @�`0AC�?`            @b@������������������������       �,����?3            @R@������������������������       ��r�j`�?-            @R@                          �<@7�Dg���?+           p|@������������������������       �v��
���?	           @y@������������������������       �t�e��?"            �I@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        j@      >@     �D@      ;@     @\@     ��@      A@     ��@      1@      @     �U@      R@     ��@     ~@      6@      n@      d@      :@      ?@      3@     �U@      @      >@      �@      ,@      @     �S@     @P@     @�@     �u@      5@     �h@      @@      @      @       @      *@     �T@      @      U@      �?       @       @      2@     �M@     @S@      @     �C@      .@       @      @      �?      *@      D@      @      =@      �?       @       @      ,@      A@      E@       @      =@      @       @              �?       @      0@      @      &@      �?                      @      5@      3@              @      &@              @              @      8@       @      2@               @       @      $@      *@      7@       @      6@      1@      �?      �?      �?              E@      �?     �K@                      @      @      9@     �A@      �?      $@      "@                                      @               @                                      @       @      �?      �?       @      �?      �?      �?             �A@      �?     �J@                      @      @      4@     �@@              "@      `@      7@      9@      1@     @R@      z@      8@     ��@      *@      @     �Q@     �G@     �|@     �p@      2@      d@     @V@      5@      0@      0@      F@      u@      2@     P@      "@             �F@      :@     �v@     �d@      ,@     @Z@      H@      "@      $@      $@      9@      e@       @     `i@       @              9@      *@     �a@     �P@      @      N@     �D@      (@      @      @      3@     �d@      $@     �r@      @              4@      *@     �k@      Y@      $@     �F@     �C@       @      "@      �?      =@      T@      @     �^@      @      @      :@      5@     @X@     @Z@      @     �K@      @@       @      "@      �?      =@     �R@      @     @Y@      @      @      6@      2@     �V@     �Y@      @     �I@      @                                      @      �?      6@                      @      @      @       @      �?      @     �H@      @      $@       @      ;@     @h@      @     �w@      @      �?       @      @     `m@     �`@      �?      E@      ;@      @      $@      @      4@     @Y@      @     �a@       @      �?      @      @      X@      M@              9@      8@      @      $@      @      4@      Y@      @     @`@       @      �?      @       @     @W@      M@              8@      7@      @      $@      @      1@      Y@      @      `@       @      �?      @       @     �V@      M@              8@      �?                              @                      �?                                      @                              @                                      �?              (@                              �?      @                      �?      6@                      @      @     @W@      �?     `m@      �?               @      @     `a@     �R@      �?      1@      @                      @      @      3@              F@                      �?             �I@      *@              @       @                      �?              @              5@                                      A@      "@               @      @                      @      @      .@              7@                      �?              1@      @              @      0@                              @     �R@      �?     �g@      �?              �?      @      V@      O@      �?      (@      0@                              @      L@      �?     `e@      �?              �?      @     �S@     �N@      �?      $@                                      �?      2@              4@                                      "@      �?               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��2jhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �=@�<h
t�?�	           ��@       	                    @ܤ��5��?	           ��@                            @4�E�4t�?�           إ@                          �:@:U���?�           ��@������������������������       ��1��
��?h           �@������������������������       ��������?k            @e@                           �?������?�           ��@������������������������       ��9
�`�?�            @t@������������������������       ���۴��?4           �@
                           �?������?4           ��@                           @��u�?�            �u@������������������������       ��L��m�?m            `d@������������������������       ��ˤ2k��?y            �g@                          �;@^bf�8�?N           ��@������������������������       ��&��d�?:           @@������������������������       ��;c�W�?             =@                           @��X���?�            �m@                           @6�X�{�?�            �i@                           �?�@�m��?/             Q@������������������������       ��鿈���?             �G@������������������������       �G���H�?             5@                           �?8�
t�F�?Q             a@������������������������       ���8��8�?             8@������������������������       �����>t�?A             \@                          �>@W3g	�?            �@@������������������������       ���!pc�?             &@������������������������       ��J����?             6@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      ?@      E@      2@      Z@     ��@     �@@     �@      9@      @     @U@     �I@     ��@     �@      3@      n@      g@      >@      E@      2@     �X@     ��@      >@     �@      3@      @      U@      G@     ��@      @      .@     �l@     �c@      .@     �A@      .@     �S@     0�@      1@     �@      ,@      @      P@      A@     p�@     u@      @     �e@     �]@      "@      <@      *@     �O@     �v@      (@     �~@      (@      @     �L@      @@     �v@     �o@      @      a@     @Y@      @      7@      *@      N@     �u@      (@     �|@      $@      @     �I@      @@     �s@     @m@      @     @^@      2@       @      @              @      3@              ?@       @              @             �G@      4@      �?      0@      D@      @      @       @      .@     @c@      @     Pq@       @              @       @      h@     �T@              B@      (@      @              �?      @      H@      @     @X@                      @      �?     @V@      A@              ;@      <@      @      @      �?      &@     �Z@       @     �f@       @               @      �?     �Y@     �H@              "@      9@      .@      @      @      5@     �b@      *@     `k@      @              4@      (@     `d@      d@      "@     �L@      .@      @      @              "@      P@      @      P@      @              @      @      R@     @P@      @      ;@      (@      @      @              @     �@@      @      <@       @                      @      8@      =@              1@      @       @      �?              @      ?@      @      B@      �?              @      @      H@      B@      @      $@      $@       @      @      @      (@     �U@      @     `c@       @              1@      @     �V@      X@      @      >@      $@       @      @      @      (@      S@      @     `a@       @              0@      @     �V@     �W@      @      >@                                              $@              0@                      �?              �?      �?                      @      �?                      @      @@      @     @Z@      @              �?      @     �F@      (@      @      &@      @      �?                      @      4@      @      X@      �?              �?      @     �D@      $@      @      &@      @      �?                      @       @      @      8@                              @      ,@      �?              @      @      �?                      @      @      @      3@                              �?      @                      @                                      �?      �?              @                              @      @      �?              @      @                                      (@              R@      �?              �?      �?      ;@      "@      @      @      �?                                       @              $@                                      @      @              �?      @                                      $@              O@      �?              �?      �?      7@      @      @      @                                      �?      (@              "@      @                              @       @                                                      �?                      @                                       @       @                                                              (@              @      @                               @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ��6hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?O�+�w�?�	           ��@       	                   �:@��y�?(           ܚ@                           @茨Tn8�?�           ,�@                          �5@�ŪF�?�           X�@������������������������       �ɂ�?��?�            �x@������������������������       ����v�{�?�             p@                           @u���]�?�            �@������������������������       � �6��f�?i            �f@������������������������       ��ک�� �?�           X�@
                            �?�x��?�            �m@                           @_B{	�%�?"             K@������������������������       �����=��?            �F@������������������������       ������H�?             "@                            �?&��M��?t            �f@������������������������       �zZcK~�?-            @S@������������������������       �
��o0:�?G            @Z@                            @P�=�x��?]           $�@                           @�n��?�           �@                          �0@�J܃K�?�           p�@������������������������       ����=A�?             C@������������������������       ��P�w#�?�           @�@                          �<@daE�(��?#           ��@������������������������       �,W�$��?�           �@������������������������       ���Bu��?5             U@                           @̡ր_<�?�           h�@                           �?�D@f�L�?�            �q@������������������������       ��;m[��?k            `e@������������������������       �/�����?C             \@                           @��}y��?�             w@������������������������       �|�f�p�?z            �i@������������������������       ���@��,�?l            `d@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �g@      8@     �F@      9@     �]@     ��@      D@     ؑ@      1@      &@     �S@      P@     `�@     �@      ,@     `o@     �V@      *@      @@      ,@     �R@     �t@      7@     pz@      "@      @      C@      ?@     �o@     @o@      @     �_@     �S@      $@      =@      ,@     @Q@     �s@      7@     �t@      @      @      =@      ?@     �j@     �k@      @     �Z@      J@      @      0@      @      7@     �a@      @     �^@      @              $@      "@     @X@     �[@             �I@      @@      @      &@              3@      S@      @     �T@                      @       @     �F@     �N@              E@      4@      �?      @      @      @      P@              D@      @              @      �?      J@      I@              "@      ;@      @      *@      $@      G@      f@      1@     �i@      @      @      3@      6@     �]@     @[@      @     �K@       @      �?      @      �?      ,@      J@       @     �D@                      �?       @      9@      3@      @       @      9@       @      "@      "@      @@      _@      "@     �d@      @      @      2@      4@     @W@     �V@             �G@      &@      @      @              @      3@             �W@      @              "@             �B@      >@              5@                                      @       @              ?@                      �?              @       @              @                                      @      @              7@                      �?              @       @              @                                              �?               @                                                                      &@      @      @              @      &@             �O@      @               @             �@@      <@              0@       @      �?       @              �?      @              $@       @               @              0@      0@              @      @       @      �?               @      @             �J@      �?                              1@      (@              "@      Y@      &@      *@      &@      F@     �v@      1@     x�@       @      @      D@     �@@      {@     pp@      &@      _@     �U@      $@      &@       @      B@     �p@      1@     �z@      @      @      C@      9@     @r@     �h@      &@     �Y@      K@      @      @      @      *@      \@      @     �h@      @              &@      (@     @^@     �N@      @      H@      @                                      (@              @                      �?       @      @       @              @     �I@      @      @      @      *@      Y@      @     `h@      @              $@      $@     @]@     �J@      @      F@      @@      @      @      @      7@     �c@      ,@     �l@       @      @      ;@      *@     `e@      a@      @      K@      @@      @      @      @      7@     �a@      (@     �h@       @      @      :@      *@     @c@      `@      @     �H@                                              0@       @     �A@                      �?              1@       @              @      ,@      �?       @      @       @      W@             r@      @      @       @       @     �a@     �P@              6@      @               @      �?      @      =@             �]@              @      �?      @     @S@      8@              ,@      @                      �?      �?      *@             @S@              @      �?      �?      C@      3@              ,@       @               @              @      0@              E@                               @     �C@      @                      "@      �?               @      @     �O@             @e@      @              �?      @     �O@      E@               @      @      �?               @       @      @@             @[@       @                              :@      6@              @      @                              �?      ?@             �N@      �?              �?      @     �B@      4@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                             �?�/��?�	           ��@       	                    @���-<G�?4           \�@                            @`�t�?=�?�           x�@                            �?�h�ű��?�           `�@������������������������       ��;_�`�?�            @v@������������������������       �@~��]��?�           ��@                          �1@�Q\.��?�            `x@������������������������       �\")�i��?             G@������������������������       �k�F	��?�            �u@
                          �<@���Q!�?�             o@                          �7@Tg�I �?�            �l@������������������������       �j b	�?w            @g@������������������������       ��GN��?!             F@                            �?x�"w���?             3@������������������������       �      �?              @������������������������       �}��7�?             &@                           �?iϢ;���?Y           d�@                            @L�+�n �?t           ��@                          �2@̣���m�?           0|@������������������������       �;��¤�?Q             a@������������������������       �K�rg`�?�            �s@                           �?n�����?b             b@������������������������       �ı��{i�?=            @U@������������������������       ��%ʍ8�?%            �M@                          �;@��B��?�           |�@                          �8@�7��8�?[           �@������������������������       ��;ͼ�?�           ��@������������������������       ��Q����?�            @l@                            @�>\^��?�            �k@������������������������       ���7OP �?V             a@������������������������       �,U,?��?4            �T@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �j@      >@      C@      :@     �V@     ؄@      E@     4�@      6@      .@     �T@     �P@     h�@     `|@      =@     �q@     @X@      2@      :@      ,@      K@     �s@      6@     �w@      1@      $@      C@      5@     �r@     @j@      "@      c@      T@      0@      7@      "@     �C@     `p@      4@     �u@      1@       @     �@@      4@     @n@     �f@      "@     �`@     �K@      $@      6@      "@     �@@     �g@      *@      l@      0@      @      <@      4@     `d@     @`@      @     �^@      .@       @      �?      @      (@     �O@      @     �Z@                      "@       @     �P@      ?@      �?      ?@      D@       @      5@      @      5@     �_@      "@     @]@      0@      @      3@      (@     @X@     �X@      @     �V@      9@      @      �?              @     @R@      @      ^@      �?      �?      @             �S@     �I@       @      *@              @                      @      @              4@                      �?                       @              @      9@      @      �?              �?      Q@      @      Y@      �?      �?      @             �S@     �E@       @      "@      1@       @      @      @      .@     �L@       @     �C@               @      @      �?      K@      =@              2@      .@       @      @      @      ,@     �L@       @     �@@               @      @      �?      H@      9@              2@      *@               @      @      ,@     �H@              :@               @      @      �?      B@      4@              *@       @       @      �?                       @       @      @                                      (@      @              @       @                              �?                      @                                      @      @                      �?                                                      @                                      �?      @                      �?                              �?                      @                                      @      �?                     @]@      (@      (@      (@      B@     �u@      4@     p�@      @      @     �F@      G@     P|@     �n@      4@     �`@      H@       @       @      @      $@     �U@      �?      e@                      "@      @     @b@      R@      �?     �C@      F@       @       @      @       @      S@      �?     �[@                      @      @     �Z@     �J@      �?      ?@      6@              �?      �?              B@              :@                      �?      �?     �@@      $@              @      6@       @      �?       @       @      D@      �?     @U@                      @      @     �R@     �E@      �?      :@      @                      �?       @      &@             �L@                       @      �?     �C@      3@               @                              �?              @              B@                       @              2@      .@               @      @                               @      @              5@                              �?      5@      @                     @Q@      $@      $@       @      :@     Pp@      3@     0�@      @      @      B@      D@     0s@     �e@      3@     �W@     �P@      $@      $@      @      7@     �k@      0@     `|@      @      @      >@     �C@     �p@      d@      3@     @S@      K@      $@      $@      @      2@     �g@      ,@     `x@      @      @      >@      A@     `j@      `@      3@     �O@      *@                              @      A@       @      P@                              @     �L@      @@              ,@       @                      �?      @     �C@      @      X@      �?      �?      @      �?     �C@      &@              1@       @                      �?      �?      3@      @     �I@      �?              @      �?      <@      "@              .@                                       @      4@             �F@              �?                      &@       @               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJ���qhG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                              @��I���?�	           ��@       	                    �?�F���?�            �@                            �?�8p�W�?*           ��@                           @x�����?           �{@������������������������       �w��$�?�            �o@������������������������       �ߗ���?z            @g@                          �=@4
j�$��?           ��@������������������������       �Rw�S��?           �@������������������������       �����W�?             :@
                            �?уI���?�           ��@                           @͆U��?�           ܒ@������������������������       �8bA���?>           (�@������������������������       �6ɱ�k�?�             s@                          �4@�JY���?�            �v@������������������������       �2�����?c            `d@������������������������       �����e�?�            �h@                           @D(^��?�           �@                           �?���[#�?.           }@                           �?iJ�`�?�            `r@������������������������       ��5[|/��?W            �`@������������������������       �0���?c            @d@                          �;@��"�P��?t            `e@������������������������       �F�B��?k            `c@������������������������       �     ��?	             0@                           �?��*k��?~           @�@                           @�i4��?�            @o@������������������������       ��~��[�?�            �l@������������������������       ��zv�X�?             6@                          @@@S�l�`�?�            �v@������������������������       ��@�n\�?�            @v@������������������������       �p=
ףp�?             $@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        k@     �C@      F@      7@      Z@     ��@      C@     x�@      <@      @     �T@     �K@     ��@     @      2@     �o@     �d@      <@     �@@      4@      V@     ~@      ?@     ��@      1@      @     �P@     �H@     8�@     �w@      1@     �j@     �Q@      0@      ?@      *@     �J@      n@      0@     pr@       @       @      ;@      :@     �i@      d@      @     @W@      8@      @      @      @      2@     �U@      @     �^@      �?              $@      @     @Q@      N@              8@      ,@      @      @      �?       @     �A@      @      U@                      @      @     �C@     �C@              $@      $@                      @      $@     �I@              C@      �?              @      @      >@      5@              ,@      G@      (@      9@       @     �A@     @c@      &@     �e@      @       @      1@      4@      a@      Y@      @     @Q@     �E@      (@      9@       @     �A@     �b@      &@      d@      @       @      1@      4@     �`@     �X@      @     �P@      @                                      @              *@                                      @       @               @     �W@      (@       @      @     �A@      n@      .@     �z@      "@       @     �C@      7@     �s@      k@      $@     �^@     @P@      &@      �?      @      3@     `g@      *@     �v@       @              6@      &@     p@     @c@      @     �T@      L@      @      �?      @      ,@      c@      $@      o@      @              ,@       @     @j@      ^@       @     �I@      "@      @              @      @     �A@      @      ]@      @               @      @     �G@      A@      @      ?@      =@      �?      �?              0@      K@       @     �O@      �?       @      1@      (@      L@     �O@      @      D@      1@              �?              @      ;@      �?      <@                      &@      @      &@      >@      @      7@      (@      �?                      $@      ;@      �?     �A@      �?       @      @      @     �F@     �@@       @      1@      J@      &@      &@      @      0@      f@      @     �x@      &@       @      0@      @     �j@      ^@      �?     �C@      .@      �?       @      �?      @     �O@      @      h@      @               @      @     �W@     �F@              5@      $@              @      �?      @      ?@      �?      a@      @              @       @     �G@      ?@              *@      @              @              @      4@      �?     �G@      @              @      �?      4@      1@              @      @              �?      �?       @      &@             �V@                      @      �?      ;@      ,@              "@      @      �?       @                      @@       @      L@                       @      �?      H@      ,@               @      @      �?      �?                      @@       @      F@                       @      �?     �G@      ,@              @                      �?                                      (@                                      �?                       @     �B@      $@      @       @      &@     @\@      @     @i@      @       @       @      @      ^@     �R@      �?      2@      5@      @       @              @     �E@      @     �P@      @       @       @       @     �C@     �A@      �?      ,@      4@      @       @              @     �C@      @     �N@      @       @       @       @      =@     �A@      �?      (@      �?                                      @              @                                      $@                       @      0@      @      �?       @      @     �Q@      �?      a@      @                      �?     @T@      D@              @      .@      @      �?       @      @     �Q@      �?     �`@      @                      �?     �R@      D@              @      �?                                                       @                                      @                        �t�bub��+      hhubh)��}�(hhhhhKhKhKhG        hh.hNhJ�5hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�B�                            �<@r��D��?�	           ��@                          �7@�^'a��?�           $�@                           !@�P�x��?�           ��@                            @�$(��?�           `�@������������������������       ��U��/�?�           @�@������������������������       ��I�O{�?�            �@������������������������       �����p9�?	             3@                          �8@������?           x�@	       
                    @ '�hG��?�            �m@������������������������       �Ą�A`��?�            �i@������������������������       ��.�?��?             >@                           @[H&�V��?�           �@������������������������       ��%M*��?U           Ȁ@������������������������       ���ě��?1            �R@                           @�[¶��?�            ps@                           @v�N�?�?�            �p@                           �?[V:��A�?I            �Z@������������������������       �j�V���?             6@������������������������       �,)&# �?=            @U@                          �?@R���Q�?l             d@������������������������       �>-\Tu�?D            �X@������������������������       �6��Hn�?(            �N@                           �?]t�E]�?             F@������������������������       �9��8���?             8@                            �?�(\����?             4@������������������������       ����Q��?             $@������������������������       �ףp=
��?             $@�t�bh�h4h7K ��h9��R�(KKKK��h��B�        f@     �B@      D@     �D@     �[@     ��@     �C@     ��@      7@      (@     �V@     �Q@     X�@      ~@      .@     `p@     �c@      B@     �C@     �D@     �Y@     ��@     �A@     P�@      4@      &@     @S@     �P@     ��@     �|@      &@     �n@     @`@      5@      B@      <@     �T@      {@      >@      �@      ,@      $@      O@      N@     Ȁ@     �u@      $@     �j@      _@      5@      B@      <@     �T@     �z@      ;@     �@      ,@      $@      O@      N@     Ȁ@     �u@      $@     �j@     �X@      0@      @@      6@      N@     t@      3@     �~@      *@      "@     �H@      K@     @w@      q@      $@     �d@      :@      @      @      @      6@      Z@       @     @o@      �?      �?      *@      @     �d@     �S@             �G@      @                                      @      @       @                                                              �?      ;@      .@      @      *@      4@     �e@      @     `p@      @      �?      .@      @     �c@     �[@      �?     �@@      @      @       @      @      @     �H@       @     @V@                       @      @     �B@      ,@              &@      @      @              @      @     �F@       @     @Q@                       @      @     �A@      ,@              "@                       @                      @              4@                                       @                       @      7@      "@      �?      $@      ,@     �^@      @     �e@      @      �?      @       @     �]@     @X@      �?      6@      5@      "@      �?       @      (@     �\@      @     �a@      @      �?      @       @     �Z@     @U@      �?      4@       @                       @       @       @              @@                       @              (@      (@               @      3@      �?      �?              "@      @@      @     ``@      @      �?      *@      @      K@      3@      @      0@      0@      �?      �?              @      8@      @     �]@      @      �?      *@      @     �C@      .@      @      0@      @      �?      �?              @      $@      �?      @@       @      �?      "@      @      0@      @      @      $@      �?                               @      @              �?                      @      �?       @      @              @      @      �?      �?              @      @      �?      ?@       @      �?      @       @      ,@      @      @      @      &@                              �?      ,@      @     �U@      �?              @      �?      7@       @      �?      @      "@                              �?      $@             �L@      �?              @              @      @      �?      @       @                                      @      @      >@                              �?      1@      @              �?      @                               @       @              (@                                      .@      @                      @                               @      �?              @                                      @      @                                                              @              @                                       @                                                                      @                                                      @                                                                      @              @                                       @                        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh.hNhJY��&hG        hNhG        h/Kh0Kh1h4h7K ��h9��R�(KK��hR�C�              �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@�t�bhFhWhZC       ���R�h_Kh`hcKh4h7K ��h9��R�(KK��hZ�C       �t�bK��R�}�(hKhmKhnh4h7K ��h9��R�(KK��hu�BX                             @sw��ͪ�?�	           ��@       	                    �?��:d���?�           $�@                           @�JĞ ��?V           ��@                          �:@��ÿ�?           �z@������������������������       ��.)kh��?�            �v@������������������������       �     ��?+             P@                            �?0mY0ɍ�?F            �[@������������������������       �	�����?(             N@������������������������       ����p��?            �I@
                           �?�Կ Y��?u           ��@                           �?P�R*�?B           `�@������������������������       �������?�            �t@������������������������       �$}����?x           �@                           @0~s}���?3           ��@������������������������       �|�"c��?D           H�@������������������������       �jpjC��?�           �@                          �:@��Tze|�?�            ps@                           @�Kg�
�?�            �n@                            �?��7Z�4�?]            �b@������������������������       ��D����?9            @W@������������������������       �>4և���?$             L@                          �3@�o�G`�?A            �X@������������������������       ���8��x�?             H@������������������������       ��{�Pk�?"             I@                            �?     L�?*             P@������������������������       �"P7��?             3@                           @��ӭ�a�?            �F@������������������������       ��vG�
�?            �@@������������������������       �      �?             (@�t�bh�h4h7K ��h9��R�(KKKK��h��B�       �k@      9@     �E@      ;@     @Z@     ��@      H@     ��@      6@      "@      S@      S@     ��@     8�@      5@      o@      k@      8@      D@      :@     �X@     �@      D@     x�@      4@      "@     �Q@     �Q@     X�@     ~@      5@     �k@     �@@      @      @       @      (@     �Q@       @     �`@      @              &@      @     �[@     @Y@      �?     �C@      7@      @      @       @      $@      N@      �?     �X@       @              &@      @      Y@     @P@      �?     �B@      2@      @      @       @      $@     �D@      �?      V@       @              @      @     @U@      O@      �?      >@      @              �?                      3@              $@                      @              .@      @              @      $@                               @      $@      �?     �A@      @                              &@      B@               @      @                                      @      �?      9@       @                              @      ,@              �?      @                               @      @              $@       @                              @      6@              �?      g@      5@      A@      8@     �U@     ��@      C@     P�@      ,@      "@     �M@     @P@     ��@     �w@      4@     �f@     �K@      @      (@      "@      2@     @e@      &@     @r@       @      @       @      &@     @e@      [@      @      H@      =@      @      (@      @      &@      O@      @     �V@       @       @      @      �?      F@      D@      �?      4@      :@      @              @      @      [@      @     @i@      @      @      @      $@     �_@      Q@      @      <@      `@      ,@      6@      .@     @Q@     �v@      ;@     0�@      @      @     �I@      K@      y@      q@      *@     �`@      B@      @      @      @      @     �W@      "@      \@       @              "@      (@     @_@     �Q@      @      >@     @W@      &@      3@      $@      O@     �p@      2@     `{@      @      @      E@      E@     Pq@      i@      $@      Z@      @      �?      @      �?      @      ?@       @     @Z@       @              @      @     @R@      C@              ;@      @      �?      @      �?      @      9@       @     �Q@       @              @      @     �N@      B@              7@       @      �?      @      �?       @      1@      @     �A@      �?              �?              J@      3@               @       @                      �?      �?      (@      @      7@      �?              �?              >@       @              @              �?      @              �?      @              (@                                      6@      &@              �?      @                              @       @      �?      B@      �?               @      @      "@      1@              .@      �?                              @      @      �?      8@                      �?              @       @              @       @                                      @              (@      �?              �?      @      @      "@              (@                                      �?      @              A@                      @       @      (@       @              @                                      �?      �?              @                      @       @      @      �?              �?                                              @              =@                                      @      �?              @                                              @              4@                                      @      �?                                                                              "@                                                              @�t�bubhhubehhub.