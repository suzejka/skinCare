���J      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K
�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�Ch                                                                	       
                     �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K
�
node_count�Kq�nodes�hhK ��h��R�(KKq��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B�         H                   �5@��=	c��?�             c@       E                    @��I���?g            �Y@       0                     @�.����?c            �X@                           �?.�r?��?E            @Q@       
                    �?����X�?             ,@                           �?      �?             @������������������������       �                     �?       	                    3@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?                           �?z�G�z�?
             $@������������������������       ��q�q�?             @������������������������       �                     @                           @Ȅ���?7            �K@                           @r֛w���?             ?@                          �2@�q�q�?             5@                           �?      �?              @������������������������       �      �?             @������������������������       �      �?             @                           �?�n_Y�K�?             *@                           �?�q�q�?	             "@                            �?      �?             @������������������������       ��q�q�?             @������������������������       �                     �?                           @z�G�z�?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �      �?             @                           �?ףp=
�?
             $@������������������������       �                     @������������������������       �r�q��?             @        !                     �?r�q��?             8@������������������������       �                     �?"       '                   �1@`������?             7@#       &                    @�8��8��?             @$       %                    �?���Q��?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     �?(       -                    �?�"�O�|�?             1@)       *                     �?      �?             @������������������������       �                     @+       ,                     @      �?              @������������������������       �                     �?������������������������       �                     �?.       /                    @�C��2(�?             &@������������������������       �                     @������������������������       �      �?             @1       :                    �?z5�h$�?             >@2       3                    �?��.k���?             1@������������������������       �                      @4       9                    3@��S���?             .@5       6                    �?      �?             ,@������������������������       �և���X�?             @7       8                   �1@և���X�?             @������������������������       �      �?              @������������������������       ����Q��?             @������������������������       �                     �?;       <                    @޾�z�<�?             *@������������������������       �                     @=       @                    @�8��8��?             @>       ?                    3@      �?              @������������������������       �                     �?������������������������       �                     �?A       D                    �?      �?             @B       C                   �3@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     �?F       G                    !@      �?             @������������������������       �                      @������������������������       �      �?              @I       ^                     �?���9#J�?2             I@J       [                    @��,d!�?             7@K       Z                    A@ԍx��?             3@L       O                    �?k��\��?             1@M       N                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @P       Q                   �6@t�E]t�?             &@������������������������       �                     @R       S                   �7@      �?              @������������������������       �                     �?T       Y                    @�$I�$I�?             @U       X                   �8@{�G�z�?             @V       W                    �?      �?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @\       ]                    9@      �?             @������������������������       �                      @������������������������       �                      @_       h                     @���v^��?             ;@`       g                   �8@     ��?             0@a       d                    @��Q��?
             $@b       c                    �?z�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @e       f                     @���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @i       n                    �?��!pc�?             &@j       m                    @      �?             @k       l                    �?�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                     �?o       p                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @�t�b�values�hhK ��h��R�(KKqKK��hV�B�-        3@      S@      *@      �?      @      �?      5@      @      @      �?       @      �?      �?      .@      Q@       @      �?      @              &@                      �?                      �?      .@      Q@       @              @              "@                                              �?      @      I@      �?              @              "@                                              �?      @      $@                                                                                               @       @                                                                                                      �?                                                                                               @      �?                                                                                              �?      �?                                                                                              �?                                                                                                       @       @                                                                                               @      @                                                                                                      @                                                                                                      D@      �?              @              "@                                              �?              7@                                       @                                                              ,@                                      @                                                              @                                       @                                                              @                                      �?                                                              @                                      �?                                                               @                                      @                                                              @                                      @                                                               @                                       @                                                               @                                      �?                                                                                                      �?                                                              @                                      �?                                                              �?                                                                                                      @                                      �?                                                               @                                       @                                                              "@                                      �?                                                              @                                                                                                      @                                      �?                                                              1@      �?              @              �?                                              �?                                                                                                      �?              1@      �?              @              �?                                                              @                       @              �?                                                              @                       @                                                                                                      �?                                                                              @                      �?                                                                                                                      �?                                                              ,@      �?               @                                                                              @      �?              �?                                                                              @                                                                                                              �?              �?                                                                                                      �?                                                                                      �?                                                                                              $@                      �?                                                                              @                                                                                                      @                      �?                                                                      &@      2@      �?                                                                                      "@       @                                                                                               @                                                                                                      @       @                                                                                              @      @                                                                                              @      @                                                                                              @      @                                                                                              �?      �?                                                                                               @      @                                                                                                      �?                                                                                               @      $@      �?                                                                                              @                                                                                               @      @      �?                                                                                      �?              �?                                                                                                      �?                                                                                      �?                                                                                                      �?      @                                                                                              �?       @                                                                                              �?      �?                                                                                                      �?                                                                                                      �?                                                                                                                      �?                       @                      �?                                                                               @                                                                              �?                                              �?                              @       @      &@              @      �?      $@      @      @               @      �?               @       @       @                      �?      "@              @               @      �?                       @       @                      �?      "@              @                      �?                       @                              �?      "@              @                      �?                                                               @              @                                                                                       @                                                                                                                      @                                               @                              �?      @                                      �?                                                              @                                                               @                              �?      @                                      �?                                                      �?                                                                       @                                      @                                      �?                       @                                       @                                      �?                       @                                       @                                                              �?                                                                                                      �?                                       @                                                                                                                                              �?                                                               @                                                                       @                                                                                       @                                                                               @                       @                                                                                                                                                                                       @                       @      @      "@              @              �?      @                                                      @      "@              @                                                                              @      @              @                                                                              @                      �?                                                                               @                      �?                                                                               @                                                                                                              @               @                                                                                                       @                                                                                      @                                                                                                      @                                                                                       @       @                                      �?      @                                              �?       @                                      �?                                                               @                                      �?                                                              �?                                                                                                      �?                                      �?                                                      �?                                                                                                      �?                                                      @                                              �?                                                                                                                                                              @                                        �t�bub�_sklearn_version��1.1.0�ub.