���]      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C�                                           	       
                                                                      �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K�
node_count�Kw�nodes�hhK ��h��R�(KKw��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B         >                   �4@J��%7)�?�             e@       +                    @���k�?T             U@       $                    @::P��P�?7            �K@                           �?�� =[�?"             A@                           �?�b-�I�?             3@       	                    �?�q�q�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?
                            �?      �?             @������������������������       �                     �?                            @�q�q�?             @������������������������       �                     �?������������������������       �      �?              @                           @g\�5�?             *@                          �3@{�G�z�?
             $@                           2@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �:/����?             @                            �?�q�q�?             @������������������������       �                     �?������������������������       �                      @       #                      @�'}�'}�?             .@                           @*x9/��?             ,@                            �?{�G�z�?             @������������������������       �                      @                           �?�q�q�?             @������������������������       �      �?              @������������������������       �                     �?       "                     �?�<ݚ�?	             "@        !                    �?����X�?             @������������������������       �      �?              @������������������������       �z�G�z�?             @������������������������       �                      @������������������������       �                     �?%       (                    �?��s����?             5@&       '                    �?      �?             (@������������������������       �r�q��?             @������������������������       ��q�q�?             @)       *                    �?�����H�?	             "@������������������������       �z�G�z�?             @������������������������       �                     @,       1                    @΃�\�?             =@-       0                    �?@4և���?             ,@.       /                     @      �?              @������������������������       �r�q��?             @������������������������       �                      @������������������������       �                     @2       9                    @�X�%��?             .@3       6                     �?ffffff�?
             $@4       5                    @�Q����?             @������������������������       �      �?             @������������������������       �                     �?7       8                    �?z�G�z�?             @������������������������       �                      @������������������������       ��q�q�?             @:       ;                    @z�G�z�?             @������������������������       �                      @<       =                    �?�q�q�?             @������������������������       �                     �?������������������������       �      �?              @?       F                     �?
�Sy'�?T             U@@       A                   �5@�8��8��?             8@������������������������       �                     @B       C                    �?>F?�!��?             5@������������������������       �                     @D       E                   �@@�����H�?             2@������������������������       �                     0@������������������������       �                      @G       Z                    7@8�&���?<             N@H       S                     @����p9�?             3@I       R                    @T�r
^N�?             ,@J       O                     �?r�q��?             (@K       L                    �?�����H�?	             "@������������������������       �                     @M       N                    @z�G�z�?             @������������������������       �                      @������������������������       ��q�q�?             @P       Q                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @T       Y                   �5@
ףp=
�?             @U       X                     @      �?             @V       W                    �?�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                     �?������������������������       �                     �?[       b                     �?��!�Ɔ�?)            �D@\       _                    �?��Q��?
             $@]       ^                    �?      �?             @������������������������       �                      @������������������������       �                      @`       a                    ?@r�q��?             @������������������������       �                     @������������������������       �                     �?c       d                    �?�߸�ǒ�?             ?@������������������������       �      �?             @e       t                   �<@T�����?             ;@f       i                    �?I�O���?             7@g       h                    @      �?              @������������������������       �                     �?������������������������       �                     �?j       s                    @Cu��?             5@k       n                     @P�|�@�?             1@l       m                    �?�q�q�?             @������������������������       �      �?              @������������������������       �                     �?o       p                     @��X��?             ,@������������������������       ��q�q�?             @q       r                    @      �?              @������������������������       �{�G�z�?             @������������������������       �VUUUUU�?             @������������������������       �                     @u       v                    @      �?             @������������������������       �                     �?������������������������       �                     @�t�b�values�hhK ��h��R�(KKwKK��hV�B8?        .@      @      @      *@      5@      (@      7@      @       @       @      @       @      @      ,@      (@      6@      @      .@                      $@      1@      @      7@                                      @      @      @              �?               @                      $@      *@      @      7@                                      �?      @                                       @                      $@      "@      @      @                                      �?      @                                       @                      �?      @      �?      @                                              @                                       @                               @      �?                                                      �?                                                                              �?                                                      �?                                                                              �?                                                                                                                                                                                              �?                                       @                               @                                                                                                                                      �?                                                                                                       @                              �?                                                                                                      �?                                                                                                                                      �?                              �?                                                                                                                              �?      @              @                                               @                                                                      @              @                                               @                                                                       @              �?                                                                                                                      �?              �?                                                                                                                      �?                                                                                                                                       @              @                                               @                                                              �?                       @                                                                                                              �?                                                                                                                                                               @                                                                                                              "@      @       @                                              �?                                                                      "@      @       @                                                                                                                       @      �?       @                                                                                                                                       @                                                                                                                       @      �?                                                                                                                              �?      �?                                                                                                                              �?                                                                                                                                      @       @                                                                                                                              @       @                                                                                                                              �?      �?                                                                                                                              @      �?                                                                                                                               @                                                                                                                                                                                                      �?                                                                              @              1@                                                                                                                      @              "@                                                                                                                      �?              @                                                                                                                       @              @                                                                                                                      �?               @                                                                                                                      �?              @                                                                                                                                      @                                                                                      *@                              @      @                                              @              @              �?              *@                              �?                                                                                                      @                              �?                                                                                                      @                              �?                                                                                                       @                                                                                                                                      @                                                                                                                                                                      @      @                                              @              @              �?                                               @      @                                                              @              �?                                              �?      @                                                                              �?                                              �?      @                                                                                                                                                                                                                      �?                                              �?                                                                      @                                                                                                                                       @                                                              �?                                                                       @                                                              �?                                                      @                                                                                                                                       @                                                                              �?                                                       @                                                                                                                                      �?                                                                              �?                                                      �?                                                      @      @      @      @      @              @       @       @      @      @      �?      $@      (@      5@      @               @              @              @                                                                              0@                                      @                                                                                                                       @                              @                                                                              0@                                                      @                                                                                                       @                                                                                                              0@                                                                                                                                      0@                       @                                                                                                                                      �?      @              @      @              @       @       @      @      @      �?      $@      (@      @      @                      �?               @       @                                               @      �?      "@               @                                              �?                                                       @              "@               @                                              �?                                                       @              "@                                                              �?                                                                       @                                                                                                                                      @                                                              �?                                                                      @                                                                                                                                       @                                                              �?                                                                       @                                                                                                                       @              �?                                                                                                                       @                                                                                                                                                      �?                                                                                                                                                       @                              �?              �?       @                                                      �?                                                      �?              �?       @                                                                                                                              �?       @                                                                                                                                      �?                                                                                                                              �?      �?                                                                                                              �?                                                                                                                                                                                                                      �?                                              �?      @               @      �?              @       @       @      @      �?              �?      (@      @      @              �?       @                                      @               @                                                                               @                                                       @                                                                               @                                                                                                                                                                                               @                                                                      �?                                              @                                                                                                                                      @                                                                                      �?                                                                                                                                               @               @      �?                       @              @      �?              �?      (@      @      @                       @                                               @                                                                                                       @      �?                                      @      �?              �?      (@      @      @                                       @      �?                                      @      �?              �?      &@              @                                              �?                                                              �?                                                                      �?                                                                                                                                                                                                      �?                                                               @                                              @      �?                      &@              @                                       @                                              @      �?                      @              @                                       @                                                      �?                                                                              �?                                                      �?                                                                              �?                                                                                                                                                                                      @                              @              @                                                                                       @                              @                                                                                                       @                              @              @                                                                                      �?                               @               @                                                                                      �?                              �?              �?                                                                                                                      @                                                                                                                                      �?      @                                                                                                                              �?                                                                                                                                              @        �t�bub�_sklearn_version��1.1.0�ub.