���      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C                              �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K�
node_count�K7�nodes�hhK ��h��R�(KK7��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B         "                     @�aZ�y�?s            �\@                           �?���`��?Q            @T@                            �?b���i��?,             F@       	                    �?Hx�5?�?$             B@                           3@���Q��?             @������������������������       �                     �?                            �?      �?             @������������������������       �      �?              @������������������������       �      �?              @
                           @w���<�?             ?@                           @hE#߼�?             >@������������������������       �>4և���?             <@������������������������       �      �?              @������������������������       �                     �?                           @      �?              @                           @      �?             @������������������������       �      �?              @������������������������       �      �?              @                           2@      �?             @������������������������       �                     �?                           5@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?                            �?�i����?%            �B@������������������������       �                     ,@                           @K����?             7@                           �?���Q��?
             $@������������������������       ��q�q�?             @������������������������       �      �?             @       !                   �2@.y0��k�?             *@                            @�Q����?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                      @#       ,                    �?Lj�����?"             A@$       '                    �?     ��?             0@%       &                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @(       +                   �2@ףp=
�?
             $@)       *                    �?�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                     @-       0                    @�[��"e�?             2@.       /                    �?      �?             @������������������������       �      �?              @������������������������       �                      @1       6                   �5@և���X�?             ,@2       5                   �2@�n_Y�K�?             *@3       4                    �?�eP*L��?             &@������������������������       ����Q��?             @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �                     �?�t�b�values�hhK ��h��R�(KK7KK��hV�B�        4@     @R@      .@      @      @     �L@      ,@      @      @      :@      "@      @      @      8@      @       @      @       @                      �?                               @       @                      �?      �?                      �?      �?                              6@      @       @              6@      @       @              5@      @      �?              �?              �?                      �?                       @       @      @               @               @              �?              �?              �?              �?                       @       @                      �?                              �?       @                      �?      �?                              �?              ?@      @      �?              ,@                              1@      @      �?              @      @                      @       @                       @       @                      &@      �?      �?              @      �?      �?                      �?                      @              �?               @                      1@      0@      �?              &@      @                       @      @                       @                                      @                      "@      �?                       @      �?                      �?                              �?      �?                      @                              @      &@      �?                      @      �?                      �?      �?                       @                      @       @                      @       @                      @      @                      @       @                       @      @                               @                      �?                        �t�bub�_sklearn_version��1.1.0�ub.