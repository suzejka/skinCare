���+      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��entropy��splitter��best��	max_depth�K�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�Ch                                                                	       
                     �t�b�
n_classes_�h�scalar���h%C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C       �t�bK��R�}�(h	K�
node_count�K?�nodes�hhK ��h��R�(KK?��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B�         8                   �8@c���J�@�             e@                           @AD$�@�            �a@                          �5@<f4P�@G            �Q@                           �?[q��g@+            �E@                           �?�:1]@             9@                           3@�ڰ`+��?
             $@������������������������       �                      @������������������������       �c�YB�d�?              @	       
                    �?������@             .@������������������������       ����� ��?             @������������������������       �//�jsx @	             "@                           �?�o�9M�?             2@                            �?M�)9��?	             "@������������������������       �                     @������������������������       ��Z���?             @                          �4@��!zȓ@	             "@������������������������       ���b}�?              @������������������������       �                     �?                           �?�� Rf��?             <@                            �?z&F�Y�?             @������������������������       �|%��b�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                           �?o�$��V�?             7@                           @*����?             6@������������������������       ��{���?             .@������������������������       �                     @������������������������       �                     �?       )                     �?��=R	@E            @Q@       $                    @�~~�x @             6@        !                     �?��!zȓ@	             "@������������������������       �                     �?"       #                    �?��b}�?              @������������������������       ��,�4�?             @������������������������       �                     �?%       (                    !@� �P��?             *@&       '                    �?�v��T��?             (@������������������������       ���'4���?              @������������������������       �                     @������������������������       �                     �?*       1                    �?v� N@/            �G@+       .                    @e%P�d�?             9@,       -                    �?z&F�Y�?             .@������������������������       ���&��?             @������������������������       �p-�"�?
             $@/       0                    6@�ڰ`+��?
             $@������������������������       �N�y�ΐ�?	             "@������������������������       �                     �?2       5                     @Dv�@� @             6@3       4                    @�J�'~x�?             0@������������������������       ��1H����?              @������������������������       ���b}�?              @6       7                    �?_�z|�X�?             @������������������������       �|%��b�?             @������������������������       �|%��b�?             @9       <                     �?��t�wK�?             <@:       ;                   �@@�!]]t�?	             "@������������������������       �                     @������������������������       �                      @=       >                     @��$�	�?             3@������������������������       �                     2@������������������������       �                     �?�t�b�values�hhK ��h��R�(KK?KK��hV�B�        �?      @      ;@      @      7@      9@      @      &@      �?      �?       @      0@     �I@      �?      @      ;@      @      7@      @      @      &@      �?      �?       @      0@      F@              @      @      @      &@      �?      @      @              �?       @      $@      ?@              @       @              "@      �?      �?      @                       @      $@      (@              @       @              @                      �?                       @      $@       @                                      �?                                               @      @                                                                                               @                                                      �?                                                      @                      @       @              @                      �?                              @       @              @      �?                                                                      �?      �?                      �?              @                      �?                               @      �?                                      @      �?      �?       @                                      $@                                      �?                                                               @                                                                                                      @                                      �?                                                              @                                      @      �?      �?       @                                       @                                      @      �?               @                                       @                                                      �?                                                                      �?      @       @               @                      �?                      3@                      �?               @                                                               @                                      �?                                                               @                      �?              �?                                                                                                      �?                                                                                      �?                                                                                                              @                       @                      �?                      1@                              @                       @                                              1@                              @                       @                                              $@                                                                                                      @                                                                              �?                              �?              8@              (@      @               @      �?                      @      *@      �?               @              @                              �?                      @      &@      �?              �?               @                                                      @       @      �?                                                                                                                      �?               @                                                      @       @                      �?               @                                                       @       @                                                                                              �?                              �?               @                              �?                              "@                      �?               @                                                              "@                      �?               @                                                              @                                                                                                      @                                                                      �?                                                      6@               @      @               @                              @       @                      *@              @                       @                              �?                              @              @                      @                                                               @                                      @                                                              @              @                      @                                                              @                                       @                              �?                              @                                      �?                              �?                                                                      �?                                                              "@              @      @                                               @       @                      "@               @      @                                                      �?                      @              �?                                                              �?                      @              �?      @                                                                                              @                                                       @      �?                                      �?                                                       @                                               @                                                              �?                              �?              4@                                                      @                                               @                                                      @                                                                                                      @                                               @                                                                                      �?              2@                                                                                                      2@                                                                                      �?                                                                        �t�bub�_sklearn_version��1.1.0�ub.